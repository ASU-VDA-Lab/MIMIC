module real_jpeg_16131_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_258;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_0),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_1),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_2),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g23 ( 
.A(n_4),
.B(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_4),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_4),
.B(n_63),
.Y(n_62)
);

AND2x4_ASAP7_75t_SL g66 ( 
.A(n_4),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_4),
.B(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_4),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_4),
.B(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_4),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_5),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_5),
.B(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_5),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_6),
.Y(n_92)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_7),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_7),
.Y(n_162)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_7),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_8),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_8),
.B(n_50),
.Y(n_49)
);

AND2x4_ASAP7_75t_SL g58 ( 
.A(n_8),
.B(n_59),
.Y(n_58)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_8),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_8),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_8),
.B(n_31),
.Y(n_107)
);

NAND2x1p5_ASAP7_75t_L g127 ( 
.A(n_8),
.B(n_128),
.Y(n_127)
);

NAND2x1_ASAP7_75t_L g170 ( 
.A(n_8),
.B(n_171),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_9),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_10),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_10),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_10),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_10),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_10),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_10),
.B(n_253),
.Y(n_252)
);

BUFx8_ASAP7_75t_L g171 ( 
.A(n_11),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_11),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_11),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_222),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_220),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_183),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_147),
.B(n_182),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_116),
.B(n_146),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_88),
.B(n_115),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_53),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_21),
.B(n_53),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.C(n_46),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_22),
.B(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_26),
.B1(n_36),
.B2(n_37),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_23),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_23),
.A2(n_36),
.B1(n_135),
.B2(n_139),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_23),
.A2(n_98),
.B(n_107),
.C(n_136),
.Y(n_154)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_27),
.A2(n_28),
.B1(n_122),
.B2(n_131),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_27),
.B(n_131),
.C(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_28),
.B(n_32),
.C(n_36),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_44),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_29),
.B(n_177),
.Y(n_176)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_32),
.A2(n_33),
.B1(n_159),
.B2(n_163),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_33),
.B(n_195),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g257 ( 
.A1(n_33),
.A2(n_258),
.B(n_259),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_35),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_38),
.A2(n_46),
.B1(n_47),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_38),
.A2(n_39),
.B(n_42),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_48),
.B1(n_49),
.B2(n_52),
.Y(n_47)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_42),
.A2(n_43),
.B1(n_57),
.B2(n_58),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_42),
.A2(n_43),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_43),
.B(n_207),
.C(n_211),
.Y(n_233)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_48),
.A2(n_49),
.B1(n_94),
.B2(n_96),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_58),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_49),
.B(n_94),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_50),
.Y(n_175)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_72),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_54),
.B(n_73),
.C(n_87),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_65),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_56),
.A2(n_104),
.B(n_108),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_56),
.A2(n_66),
.B(n_71),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_66),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_66),
.A2(n_91),
.B(n_93),
.C(n_98),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_91),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_66),
.A2(n_70),
.B1(n_91),
.B2(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_69),
.B(n_122),
.C(n_127),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_86),
.B2(n_87),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_85),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_75),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_75),
.B(n_79),
.C(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_79),
.A2(n_235),
.B1(n_236),
.B2(n_240),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_79),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_81),
.Y(n_179)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_82),
.A2(n_143),
.B1(n_158),
.B2(n_164),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_85),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_102),
.B(n_114),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_99),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_91),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_91),
.B(n_106),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g190 ( 
.A(n_91),
.B(n_107),
.C(n_170),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_91),
.A2(n_112),
.B1(n_194),
.B2(n_200),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_91),
.B(n_196),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_94),
.A2(n_96),
.B1(n_159),
.B2(n_163),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_94),
.B(n_143),
.C(n_159),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_110),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_109),
.B(n_113),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_106),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_106),
.A2(n_107),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_112),
.B(n_195),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_118),
.Y(n_146)
);

XOR2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_133),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_132),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_132),
.C(n_133),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_126),
.B1(n_127),
.B2(n_131),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_122),
.Y(n_131)
);

OR2x6_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_140),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_141),
.C(n_145),
.Y(n_151)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_149),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_165),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_152),
.C(n_165),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_157),
.C(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_181),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_173),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_173),
.C(n_181),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_172),
.Y(n_167)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_176),
.B(n_180),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_176),
.Y(n_180)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_180),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_185),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_203),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_186),
.B(n_204),
.C(n_219),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_201),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_192),
.C(n_201),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_194),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_219),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_215),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_217),
.C(n_218),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_261),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_260),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_225),
.B(n_260),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_244),
.B2(n_245),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_231)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_236),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_241),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2x1_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_256),
.B2(n_257),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);


endmodule