module fake_aes_4821_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
NOR2xp33_ASAP7_75t_L g4 ( .A(n_0), .B(n_2), .Y(n_4) );
HB1xp67_ASAP7_75t_L g5 ( .A(n_3), .Y(n_5) );
AOI22xp33_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
AOI322xp5_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_7), .A3(n_6), .B1(n_4), .B2(n_1), .C1(n_0), .C2(n_2), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
AO21x2_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_0), .B(n_1), .Y(n_11) );
endmodule