module real_aes_8036_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_379;
wire n_374;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_449;
wire n_363;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_0), .A2(n_180), .B1(n_181), .B2(n_182), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_0), .Y(n_180) );
INVx1_ASAP7_75t_L g227 ( .A(n_1), .Y(n_227) );
AOI21xp33_ASAP7_75t_L g271 ( .A1(n_2), .A2(n_243), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g200 ( .A(n_3), .Y(n_200) );
AND2x6_ASAP7_75t_L g221 ( .A(n_3), .B(n_198), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_3), .B(n_530), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_4), .A2(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g277 ( .A(n_5), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_6), .B(n_306), .Y(n_305) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_6), .Y(n_525) );
AO22x2_ASAP7_75t_L g85 ( .A1(n_7), .A2(n_26), .B1(n_86), .B2(n_87), .Y(n_85) );
INVx1_ASAP7_75t_L g213 ( .A(n_8), .Y(n_213) );
INVx1_ASAP7_75t_L g331 ( .A(n_9), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_10), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_11), .A2(n_80), .B1(n_177), .B2(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_11), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_12), .B(n_248), .Y(n_319) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_13), .A2(n_27), .B1(n_86), .B2(n_90), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_14), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_15), .B(n_243), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_16), .B(n_255), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g328 ( .A1(n_17), .A2(n_329), .B(n_330), .C(n_332), .Y(n_328) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_18), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_19), .B(n_231), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_20), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_21), .A2(n_51), .B1(n_151), .B2(n_155), .Y(n_150) );
INVx1_ASAP7_75t_L g266 ( .A(n_22), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_23), .Y(n_97) );
AOI211xp5_ASAP7_75t_L g81 ( .A1(n_24), .A2(n_82), .B(n_96), .C(n_123), .Y(n_81) );
INVx2_ASAP7_75t_L g219 ( .A(n_25), .Y(n_219) );
OAI221xp5_ASAP7_75t_L g191 ( .A1(n_27), .A2(n_40), .B1(n_50), .B2(n_192), .C(n_193), .Y(n_191) );
INVxp67_ASAP7_75t_L g194 ( .A(n_27), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g289 ( .A1(n_28), .A2(n_221), .B(n_223), .C(n_290), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g140 ( .A1(n_29), .A2(n_55), .B1(n_141), .B2(n_146), .Y(n_140) );
INVx1_ASAP7_75t_L g264 ( .A(n_30), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_31), .B(n_231), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g111 ( .A1(n_32), .A2(n_56), .B1(n_112), .B2(n_117), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_33), .B(n_106), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g267 ( .A(n_34), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_35), .B(n_243), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_36), .Y(n_124) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_37), .A2(n_223), .B1(n_233), .B2(n_262), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g298 ( .A(n_38), .Y(n_298) );
CKINVDCx16_ASAP7_75t_R g215 ( .A(n_39), .Y(n_215) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_40), .A2(n_61), .B1(n_86), .B2(n_90), .Y(n_93) );
INVxp67_ASAP7_75t_L g195 ( .A(n_40), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_41), .A2(n_80), .B1(n_176), .B2(n_177), .Y(n_79) );
CKINVDCx14_ASAP7_75t_R g176 ( .A(n_41), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_42), .A2(n_251), .B(n_275), .C(n_276), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_43), .Y(n_322) );
INVx1_ASAP7_75t_L g273 ( .A(n_44), .Y(n_273) );
INVx1_ASAP7_75t_L g198 ( .A(n_45), .Y(n_198) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_46), .Y(n_183) );
OAI22xp5_ASAP7_75t_SL g182 ( .A1(n_47), .A2(n_183), .B1(n_184), .B2(n_185), .Y(n_182) );
INVx1_ASAP7_75t_L g185 ( .A(n_47), .Y(n_185) );
INVx1_ASAP7_75t_L g212 ( .A(n_48), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_49), .Y(n_192) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_50), .A2(n_66), .B1(n_86), .B2(n_87), .Y(n_95) );
INVx1_ASAP7_75t_L g172 ( .A(n_52), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_SL g247 ( .A1(n_53), .A2(n_248), .B(n_249), .C(n_251), .Y(n_247) );
INVxp67_ASAP7_75t_L g250 ( .A(n_54), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_57), .Y(n_269) );
INVx1_ASAP7_75t_L g315 ( .A(n_58), .Y(n_315) );
A2O1A1Ixp33_ASAP7_75t_L g316 ( .A1(n_59), .A2(n_221), .B(n_223), .C(n_317), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_60), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_62), .B(n_228), .Y(n_291) );
INVx2_ASAP7_75t_L g210 ( .A(n_63), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_64), .A2(n_179), .B1(n_186), .B2(n_187), .Y(n_178) );
INVx1_ASAP7_75t_L g186 ( .A(n_64), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_64), .B(n_248), .Y(n_292) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_65), .A2(n_221), .B(n_223), .C(n_226), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_67), .B(n_238), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_68), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_69), .A2(n_221), .B(n_223), .C(n_303), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_70), .Y(n_310) );
INVx1_ASAP7_75t_L g246 ( .A(n_71), .Y(n_246) );
CKINVDCx16_ASAP7_75t_R g327 ( .A(n_72), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_73), .B(n_228), .Y(n_304) );
INVx1_ASAP7_75t_L g537 ( .A(n_73), .Y(n_537) );
INVx1_ASAP7_75t_L g86 ( .A(n_74), .Y(n_86) );
INVx1_ASAP7_75t_L g88 ( .A(n_74), .Y(n_88) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_75), .B(n_241), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_76), .A2(n_243), .B(n_244), .Y(n_242) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_188), .B1(n_201), .B2(n_517), .C(n_523), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_178), .Y(n_78) );
INVx1_ASAP7_75t_L g177 ( .A(n_80), .Y(n_177) );
AOI22xp5_ASAP7_75t_SL g524 ( .A1(n_80), .A2(n_177), .B1(n_525), .B2(n_526), .Y(n_524) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_138), .Y(n_80) );
BUFx3_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
AND2x6_ASAP7_75t_L g83 ( .A(n_84), .B(n_91), .Y(n_83) );
AND2x4_ASAP7_75t_L g120 ( .A(n_84), .B(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g84 ( .A(n_85), .B(n_89), .Y(n_84) );
INVx2_ASAP7_75t_L g103 ( .A(n_85), .Y(n_103) );
AND2x2_ASAP7_75t_L g116 ( .A(n_85), .B(n_93), .Y(n_116) );
INVx1_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx1_ASAP7_75t_L g90 ( .A(n_88), .Y(n_90) );
AND2x2_ASAP7_75t_L g102 ( .A(n_89), .B(n_103), .Y(n_102) );
OR2x2_ASAP7_75t_L g110 ( .A(n_89), .B(n_103), .Y(n_110) );
INVx1_ASAP7_75t_L g115 ( .A(n_89), .Y(n_115) );
INVx2_ASAP7_75t_L g130 ( .A(n_89), .Y(n_130) );
AND2x6_ASAP7_75t_L g162 ( .A(n_91), .B(n_109), .Y(n_162) );
AND2x4_ASAP7_75t_L g165 ( .A(n_91), .B(n_102), .Y(n_165) );
AND2x2_ASAP7_75t_L g171 ( .A(n_91), .B(n_145), .Y(n_171) );
AND2x2_ASAP7_75t_L g91 ( .A(n_92), .B(n_94), .Y(n_91) );
AND2x2_ASAP7_75t_L g104 ( .A(n_92), .B(n_95), .Y(n_104) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_93), .B(n_95), .Y(n_149) );
AND2x2_ASAP7_75t_L g154 ( .A(n_93), .B(n_122), .Y(n_154) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g122 ( .A(n_95), .Y(n_122) );
INVx1_ASAP7_75t_L g129 ( .A(n_95), .Y(n_129) );
OAI211xp5_ASAP7_75t_L g96 ( .A1(n_97), .A2(n_98), .B(n_105), .C(n_111), .Y(n_96) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
BUFx3_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
NAND2x1p5_ASAP7_75t_L g101 ( .A(n_102), .B(n_104), .Y(n_101) );
AND2x2_ASAP7_75t_L g153 ( .A(n_102), .B(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g145 ( .A(n_103), .B(n_130), .Y(n_145) );
AND2x4_ASAP7_75t_L g108 ( .A(n_104), .B(n_109), .Y(n_108) );
AND2x4_ASAP7_75t_L g144 ( .A(n_104), .B(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx4_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_116), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x6_ASAP7_75t_L g156 ( .A(n_115), .B(n_149), .Y(n_156) );
AND2x4_ASAP7_75t_L g127 ( .A(n_116), .B(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g136 ( .A(n_116), .B(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B1(n_131), .B2(n_132), .Y(n_123) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
INVx1_ASAP7_75t_L g137 ( .A(n_129), .Y(n_137) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx12f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NOR3xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_157), .C(n_166), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_150), .Y(n_139) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx4_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_L g147 ( .A(n_145), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_145), .B(n_154), .Y(n_175) );
BUFx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx8_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B1(n_163), .B2(n_164), .Y(n_157) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx11_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx6_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B1(n_172), .B2(n_173), .Y(n_166) );
INVx1_ASAP7_75t_SL g168 ( .A(n_169), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_179), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_183), .Y(n_184) );
CKINVDCx16_ASAP7_75t_R g188 ( .A(n_189), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_190), .Y(n_189) );
AND3x1_ASAP7_75t_SL g190 ( .A(n_191), .B(n_196), .C(n_199), .Y(n_190) );
INVxp67_ASAP7_75t_L g530 ( .A(n_191), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
INVx1_ASAP7_75t_SL g531 ( .A(n_196), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_196), .A2(n_534), .B(n_536), .Y(n_533) );
INVx1_ASAP7_75t_L g543 ( .A(n_196), .Y(n_543) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_197), .B(n_200), .Y(n_536) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OR2x2_ASAP7_75t_SL g542 ( .A(n_199), .B(n_543), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_200), .Y(n_199) );
OR4x1_ASAP7_75t_L g201 ( .A(n_202), .B(n_406), .C(n_466), .D(n_493), .Y(n_201) );
NAND4xp25_ASAP7_75t_SL g202 ( .A(n_203), .B(n_354), .C(n_385), .D(n_402), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_279), .B(n_281), .C(n_334), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_257), .Y(n_204) );
INVx1_ASAP7_75t_L g396 ( .A(n_205), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_205), .A2(n_437), .B1(n_485), .B2(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_239), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_206), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g347 ( .A(n_206), .B(n_259), .Y(n_347) );
AND2x2_ASAP7_75t_L g389 ( .A(n_206), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_206), .B(n_280), .Y(n_401) );
INVx1_ASAP7_75t_L g441 ( .A(n_206), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_206), .B(n_495), .Y(n_494) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g369 ( .A(n_207), .B(n_259), .Y(n_369) );
INVx3_ASAP7_75t_L g373 ( .A(n_207), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_207), .B(n_431), .Y(n_430) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_214), .B(n_235), .Y(n_207) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_208), .A2(n_260), .B(n_268), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_208), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g296 ( .A(n_208), .Y(n_296) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_209), .Y(n_241) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
AND2x2_ASAP7_75t_SL g238 ( .A(n_210), .B(n_211), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_222), .Y(n_214) );
OAI22xp33_ASAP7_75t_L g260 ( .A1(n_216), .A2(n_253), .B1(n_261), .B2(n_267), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_216), .A2(n_315), .B(n_316), .Y(n_314) );
NAND2x1p5_ASAP7_75t_L g216 ( .A(n_217), .B(n_221), .Y(n_216) );
AND2x4_ASAP7_75t_L g243 ( .A(n_217), .B(n_221), .Y(n_243) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_220), .Y(n_217) );
INVx1_ASAP7_75t_L g522 ( .A(n_218), .Y(n_522) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g224 ( .A(n_219), .Y(n_224) );
INVx1_ASAP7_75t_L g234 ( .A(n_219), .Y(n_234) );
INVx1_ASAP7_75t_L g225 ( .A(n_220), .Y(n_225) );
INVx3_ASAP7_75t_L g229 ( .A(n_220), .Y(n_229) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_220), .Y(n_231) );
INVx1_ASAP7_75t_L g248 ( .A(n_220), .Y(n_248) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_220), .Y(n_263) );
INVx4_ASAP7_75t_SL g253 ( .A(n_221), .Y(n_253) );
INVx5_ASAP7_75t_L g245 ( .A(n_223), .Y(n_245) );
AND2x6_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_224), .Y(n_252) );
BUFx3_ASAP7_75t_L g295 ( .A(n_224), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_230), .C(n_232), .Y(n_226) );
INVx5_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_229), .B(n_250), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_229), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g275 ( .A(n_231), .Y(n_275) );
INVx4_ASAP7_75t_L g306 ( .A(n_231), .Y(n_306) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_237), .B(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_237), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g300 ( .A(n_238), .Y(n_300) );
OA21x2_ASAP7_75t_L g323 ( .A1(n_238), .A2(n_324), .B(n_333), .Y(n_323) );
AND2x2_ASAP7_75t_L g460 ( .A(n_239), .B(n_270), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_239), .B(n_373), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_239), .B(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g280 ( .A(n_240), .B(n_259), .Y(n_280) );
INVx1_ASAP7_75t_L g342 ( .A(n_240), .Y(n_342) );
BUFx2_ASAP7_75t_L g346 ( .A(n_240), .Y(n_346) );
AND2x2_ASAP7_75t_L g390 ( .A(n_240), .B(n_258), .Y(n_390) );
OR2x2_ASAP7_75t_L g429 ( .A(n_240), .B(n_258), .Y(n_429) );
AND2x2_ASAP7_75t_L g454 ( .A(n_240), .B(n_270), .Y(n_454) );
AND2x2_ASAP7_75t_L g513 ( .A(n_240), .B(n_343), .Y(n_513) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_254), .Y(n_240) );
INVx4_ASAP7_75t_L g256 ( .A(n_241), .Y(n_256) );
BUFx2_ASAP7_75t_L g325 ( .A(n_243), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_247), .C(n_253), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g272 ( .A1(n_245), .A2(n_253), .B(n_273), .C(n_274), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g326 ( .A1(n_245), .A2(n_253), .B(n_327), .C(n_328), .Y(n_326) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_252), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_253), .B(n_521), .Y(n_520) );
OA21x2_ASAP7_75t_L g270 ( .A1(n_255), .A2(n_271), .B(n_278), .Y(n_270) );
INVx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_SL g297 ( .A(n_256), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g488 ( .A(n_257), .Y(n_488) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_270), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_258), .B(n_270), .Y(n_374) );
AND2x2_ASAP7_75t_L g384 ( .A(n_258), .B(n_373), .Y(n_384) );
BUFx2_ASAP7_75t_L g395 ( .A(n_258), .Y(n_395) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g417 ( .A(n_259), .B(n_270), .Y(n_417) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_259), .Y(n_472) );
OAI22xp5_ASAP7_75t_SL g262 ( .A1(n_263), .A2(n_264), .B1(n_265), .B2(n_266), .Y(n_262) );
INVx2_ASAP7_75t_L g265 ( .A(n_263), .Y(n_265) );
INVx4_ASAP7_75t_L g329 ( .A(n_263), .Y(n_329) );
INVx2_ASAP7_75t_L g519 ( .A(n_265), .Y(n_519) );
AND2x2_ASAP7_75t_SL g279 ( .A(n_270), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_SL g343 ( .A(n_270), .Y(n_343) );
BUFx2_ASAP7_75t_L g368 ( .A(n_270), .Y(n_368) );
INVx2_ASAP7_75t_L g387 ( .A(n_270), .Y(n_387) );
AND2x2_ASAP7_75t_L g449 ( .A(n_270), .B(n_373), .Y(n_449) );
AOI321xp33_ASAP7_75t_L g468 ( .A1(n_279), .A2(n_469), .A3(n_470), .B1(n_471), .B2(n_473), .C(n_474), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_280), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_280), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g462 ( .A(n_280), .B(n_441), .Y(n_462) );
AND2x2_ASAP7_75t_L g495 ( .A(n_280), .B(n_387), .Y(n_495) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_311), .Y(n_282) );
OR2x2_ASAP7_75t_L g397 ( .A(n_283), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_299), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx3_ASAP7_75t_L g349 ( .A(n_286), .Y(n_349) );
AND2x2_ASAP7_75t_L g359 ( .A(n_286), .B(n_313), .Y(n_359) );
AND2x2_ASAP7_75t_L g364 ( .A(n_286), .B(n_339), .Y(n_364) );
INVx1_ASAP7_75t_L g381 ( .A(n_286), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_286), .B(n_362), .Y(n_400) );
AND2x2_ASAP7_75t_L g405 ( .A(n_286), .B(n_338), .Y(n_405) );
OR2x2_ASAP7_75t_L g437 ( .A(n_286), .B(n_426), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_286), .B(n_350), .Y(n_476) );
AND2x2_ASAP7_75t_L g510 ( .A(n_286), .B(n_336), .Y(n_510) );
OR2x6_ASAP7_75t_L g286 ( .A(n_287), .B(n_297), .Y(n_286) );
AOI21xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_289), .B(n_296), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_292), .B(n_293), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_293), .A2(n_318), .B(n_319), .Y(n_317) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g332 ( .A(n_295), .Y(n_332) );
INVx1_ASAP7_75t_L g320 ( .A(n_296), .Y(n_320) );
INVx1_ASAP7_75t_L g337 ( .A(n_299), .Y(n_337) );
INVx2_ASAP7_75t_L g352 ( .A(n_299), .Y(n_352) );
AND2x2_ASAP7_75t_L g392 ( .A(n_299), .B(n_363), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_299), .B(n_339), .Y(n_414) );
AO21x2_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B(n_309), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_308), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B(n_307), .Y(n_303) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g498 ( .A(n_312), .B(n_349), .Y(n_498) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_323), .Y(n_312) );
INVx2_ASAP7_75t_L g339 ( .A(n_313), .Y(n_339) );
AND2x2_ASAP7_75t_L g492 ( .A(n_313), .B(n_352), .Y(n_492) );
AO21x2_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_320), .B(n_321), .Y(n_313) );
AND2x2_ASAP7_75t_L g338 ( .A(n_323), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g353 ( .A(n_323), .Y(n_353) );
INVx1_ASAP7_75t_L g363 ( .A(n_323), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_329), .B(n_331), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_340), .B1(n_344), .B2(n_348), .Y(n_334) );
OAI22xp33_ASAP7_75t_L g489 ( .A1(n_335), .A2(n_453), .B1(n_490), .B2(n_491), .Y(n_489) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g404 ( .A(n_337), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_338), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g399 ( .A(n_339), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_339), .B(n_352), .Y(n_426) );
INVx1_ASAP7_75t_L g442 ( .A(n_339), .Y(n_442) );
AND2x2_ASAP7_75t_L g383 ( .A(n_341), .B(n_384), .Y(n_383) );
INVx3_ASAP7_75t_SL g422 ( .A(n_341), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_341), .B(n_347), .Y(n_499) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g508 ( .A(n_344), .Y(n_508) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_345), .B(n_441), .Y(n_483) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx3_ASAP7_75t_SL g388 ( .A(n_347), .Y(n_388) );
NAND2x1_ASAP7_75t_SL g348 ( .A(n_349), .B(n_350), .Y(n_348) );
AND2x2_ASAP7_75t_L g409 ( .A(n_349), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g416 ( .A(n_349), .B(n_353), .Y(n_416) );
AND2x2_ASAP7_75t_L g421 ( .A(n_349), .B(n_362), .Y(n_421) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_349), .Y(n_470) );
OAI311xp33_ASAP7_75t_L g493 ( .A1(n_350), .A2(n_494), .A3(n_496), .B1(n_497), .C1(n_507), .Y(n_493) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g506 ( .A(n_351), .B(n_379), .Y(n_506) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
AND2x2_ASAP7_75t_L g362 ( .A(n_352), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g410 ( .A(n_352), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g465 ( .A(n_352), .Y(n_465) );
INVx1_ASAP7_75t_L g358 ( .A(n_353), .Y(n_358) );
INVx1_ASAP7_75t_L g378 ( .A(n_353), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_353), .B(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g411 ( .A(n_353), .Y(n_411) );
AOI221xp5_ASAP7_75t_SL g354 ( .A1(n_355), .A2(n_357), .B1(n_365), .B2(n_370), .C(n_375), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_360), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx4_ASAP7_75t_L g379 ( .A(n_359), .Y(n_379) );
AND2x2_ASAP7_75t_L g473 ( .A(n_359), .B(n_392), .Y(n_473) );
AND2x2_ASAP7_75t_L g480 ( .A(n_359), .B(n_362), .Y(n_480) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_362), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g391 ( .A(n_364), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_367), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g516 ( .A(n_369), .B(n_460), .Y(n_516) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g501 ( .A(n_373), .B(n_429), .Y(n_501) );
OAI211xp5_ASAP7_75t_L g466 ( .A1(n_374), .A2(n_467), .B(n_468), .C(n_481), .Y(n_466) );
AOI21xp33_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_380), .B(n_382), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NOR2xp67_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g445 ( .A(n_379), .Y(n_445) );
OAI221xp5_ASAP7_75t_L g474 ( .A1(n_380), .A2(n_475), .B1(n_476), .B2(n_477), .C(n_478), .Y(n_474) );
AND2x2_ASAP7_75t_L g451 ( .A(n_381), .B(n_392), .Y(n_451) );
AND2x2_ASAP7_75t_L g504 ( .A(n_381), .B(n_399), .Y(n_504) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_384), .B(n_422), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_389), .B(n_391), .C(n_393), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
AND2x2_ASAP7_75t_L g432 ( .A(n_387), .B(n_390), .Y(n_432) );
OR2x2_ASAP7_75t_L g475 ( .A(n_387), .B(n_429), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_388), .B(n_454), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_388), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_SL g419 ( .A(n_389), .Y(n_419) );
INVx1_ASAP7_75t_L g485 ( .A(n_392), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_397), .B1(n_400), .B2(n_401), .Y(n_393) );
INVx1_ASAP7_75t_L g408 ( .A(n_394), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_395), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g471 ( .A(n_396), .B(n_472), .Y(n_471) );
INVxp67_ASAP7_75t_L g457 ( .A(n_398), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_399), .B(n_485), .Y(n_484) );
OAI22xp33_ASAP7_75t_L g458 ( .A1(n_400), .A2(n_459), .B1(n_461), .B2(n_463), .Y(n_458) );
INVx1_ASAP7_75t_L g467 ( .A(n_403), .Y(n_467) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
AND2x2_ASAP7_75t_L g509 ( .A(n_404), .B(n_504), .Y(n_509) );
AOI222xp33_ASAP7_75t_L g438 ( .A1(n_405), .A2(n_439), .B1(n_442), .B2(n_443), .C1(n_446), .C2(n_447), .Y(n_438) );
NAND4xp25_ASAP7_75t_SL g406 ( .A(n_407), .B(n_427), .C(n_438), .D(n_450), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_412), .B2(n_417), .C(n_418), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_410), .B(n_445), .Y(n_444) );
INVxp67_ASAP7_75t_L g436 ( .A(n_411), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_412), .A2(n_482), .B1(n_484), .B2(n_486), .C(n_489), .Y(n_481) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g424 ( .A(n_416), .B(n_425), .Y(n_424) );
OAI21xp33_ASAP7_75t_L g478 ( .A1(n_417), .A2(n_479), .B(n_480), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B1(n_422), .B2(n_423), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI21xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B(n_433), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g469 ( .A(n_440), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_441), .B(n_460), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_441), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_445), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g477 ( .A(n_449), .Y(n_477) );
AOI221xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B1(n_455), .B2(n_457), .C(n_458), .Y(n_450) );
INVxp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI222xp33_ASAP7_75t_L g497 ( .A1(n_460), .A2(n_498), .B1(n_499), .B2(n_500), .C1(n_502), .C2(n_505), .Y(n_497) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_464), .B(n_504), .Y(n_503) );
INVxp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g496 ( .A(n_470), .Y(n_496) );
INVxp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVxp33_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AOI221xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B1(n_510), .B2(n_511), .C(n_514), .Y(n_507) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVxp67_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
INVx1_ASAP7_75t_L g535 ( .A(n_518), .Y(n_535) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_521), .B(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OAI322xp33_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_527), .A3(n_531), .B1(n_532), .B2(n_537), .C1(n_538), .C2(n_540), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_525), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
endmodule