module fake_aes_3649_n_33 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
BUFx3_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_3), .B(n_4), .Y(n_13) );
AND2x2_ASAP7_75t_R g14 ( .A(n_3), .B(n_7), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_1), .Y(n_15) );
BUFx6f_ASAP7_75t_L g16 ( .A(n_12), .Y(n_16) );
AND2x4_ASAP7_75t_L g17 ( .A(n_11), .B(n_0), .Y(n_17) );
INVx2_ASAP7_75t_SL g18 ( .A(n_12), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
AOI22xp33_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_11), .B1(n_13), .B2(n_15), .Y(n_20) );
AOI22xp33_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_17), .B1(n_18), .B2(n_16), .Y(n_21) );
NOR5xp2_ASAP7_75t_SL g22 ( .A(n_19), .B(n_14), .C(n_1), .D(n_2), .E(n_4), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_21), .B(n_17), .Y(n_23) );
AND4x1_ASAP7_75t_L g24 ( .A(n_22), .B(n_0), .C(n_17), .D(n_18), .Y(n_24) );
NOR2xp33_ASAP7_75t_R g25 ( .A(n_23), .B(n_5), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
CKINVDCx20_ASAP7_75t_R g28 ( .A(n_25), .Y(n_28) );
NOR4xp75_ASAP7_75t_L g29 ( .A(n_28), .B(n_22), .C(n_8), .D(n_9), .Y(n_29) );
NOR3xp33_ASAP7_75t_SL g30 ( .A(n_27), .B(n_16), .C(n_6), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
OR2x6_ASAP7_75t_L g32 ( .A(n_30), .B(n_16), .Y(n_32) );
OAI22xp5_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_16), .B1(n_28), .B2(n_32), .Y(n_33) );
endmodule