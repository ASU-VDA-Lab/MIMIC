module real_aes_1186_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_453;
wire n_374;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_564;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_552;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
AO22x2_ASAP7_75t_L g102 ( .A1(n_0), .A2(n_55), .B1(n_90), .B2(n_103), .Y(n_102) );
AOI22xp33_ASAP7_75t_L g120 ( .A1(n_1), .A2(n_20), .B1(n_121), .B2(n_124), .Y(n_120) );
INVx1_ASAP7_75t_L g185 ( .A(n_2), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_3), .B(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g267 ( .A(n_4), .Y(n_267) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_5), .A2(n_16), .B1(n_90), .B2(n_100), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_6), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g108 ( .A1(n_7), .A2(n_48), .B1(n_109), .B2(n_114), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_8), .B(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g200 ( .A(n_9), .Y(n_200) );
INVx1_ASAP7_75t_L g246 ( .A(n_10), .Y(n_246) );
INVx1_ASAP7_75t_L g243 ( .A(n_11), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_11), .A2(n_80), .B1(n_163), .B2(n_243), .Y(n_551) );
INVx1_ASAP7_75t_SL g218 ( .A(n_12), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_13), .B(n_221), .Y(n_327) );
AOI33xp33_ASAP7_75t_L g295 ( .A1(n_14), .A2(n_39), .A3(n_206), .B1(n_214), .B2(n_296), .B3(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g276 ( .A(n_15), .Y(n_276) );
OAI221xp5_ASAP7_75t_L g177 ( .A1(n_16), .A2(n_55), .B1(n_57), .B2(n_178), .C(n_180), .Y(n_177) );
OR2x2_ASAP7_75t_L g201 ( .A(n_17), .B(n_70), .Y(n_201) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_17), .A2(n_70), .B(n_200), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_18), .B(n_204), .Y(n_203) );
INVx3_ASAP7_75t_L g90 ( .A(n_19), .Y(n_90) );
AOI22xp33_ASAP7_75t_L g155 ( .A1(n_21), .A2(n_35), .B1(n_156), .B2(n_158), .Y(n_155) );
INVx1_ASAP7_75t_SL g95 ( .A(n_22), .Y(n_95) );
INVx1_ASAP7_75t_L g187 ( .A(n_23), .Y(n_187) );
AND2x2_ASAP7_75t_L g209 ( .A(n_23), .B(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g227 ( .A(n_23), .B(n_185), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g278 ( .A(n_24), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_25), .A2(n_64), .B1(n_169), .B2(n_170), .Y(n_168) );
INVx1_ASAP7_75t_L g170 ( .A(n_25), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_26), .B(n_204), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_27), .A2(n_230), .B1(n_236), .B2(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_28), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_29), .B(n_221), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_30), .A2(n_45), .B1(n_149), .B2(n_151), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g84 ( .A1(n_31), .A2(n_68), .B1(n_85), .B2(n_104), .Y(n_84) );
OAI22xp5_ASAP7_75t_L g79 ( .A1(n_32), .A2(n_80), .B1(n_162), .B2(n_163), .Y(n_79) );
INVx1_ASAP7_75t_L g162 ( .A(n_32), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_33), .B(n_264), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g126 ( .A1(n_34), .A2(n_66), .B1(n_127), .B2(n_130), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_36), .B(n_221), .Y(n_268) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_37), .A2(n_57), .B1(n_90), .B2(n_91), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_38), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_40), .B(n_221), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_41), .Y(n_135) );
INVx1_ASAP7_75t_L g207 ( .A(n_42), .Y(n_207) );
INVx1_ASAP7_75t_L g223 ( .A(n_42), .Y(n_223) );
AND2x2_ASAP7_75t_L g308 ( .A(n_43), .B(n_198), .Y(n_308) );
INVx1_ASAP7_75t_L g167 ( .A(n_44), .Y(n_167) );
AOI221xp5_ASAP7_75t_L g265 ( .A1(n_44), .A2(n_59), .B1(n_204), .B2(n_212), .C(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g96 ( .A(n_46), .Y(n_96) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_47), .B(n_204), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_49), .B(n_230), .Y(n_285) );
AOI21xp5_ASAP7_75t_SL g255 ( .A1(n_50), .A2(n_212), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g239 ( .A(n_51), .Y(n_239) );
INVx1_ASAP7_75t_L g306 ( .A(n_52), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_53), .A2(n_80), .B1(n_163), .B2(n_558), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_53), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_54), .A2(n_212), .B(n_305), .Y(n_304) );
INVxp33_ASAP7_75t_L g182 ( .A(n_55), .Y(n_182) );
INVx1_ASAP7_75t_L g210 ( .A(n_56), .Y(n_210) );
INVx1_ASAP7_75t_L g225 ( .A(n_56), .Y(n_225) );
INVxp67_ASAP7_75t_L g181 ( .A(n_57), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_58), .B(n_204), .Y(n_298) );
AND2x2_ASAP7_75t_L g228 ( .A(n_60), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g240 ( .A(n_61), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_62), .A2(n_212), .B(n_217), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g325 ( .A1(n_63), .A2(n_212), .B(n_290), .C(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g169 ( .A(n_64), .Y(n_169) );
AND2x2_ASAP7_75t_SL g253 ( .A(n_65), .B(n_229), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_67), .A2(n_212), .B1(n_293), .B2(n_294), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_69), .B(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g257 ( .A(n_71), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_72), .A2(n_165), .B1(n_172), .B2(n_173), .Y(n_164) );
INVx1_ASAP7_75t_L g172 ( .A(n_72), .Y(n_172) );
AND2x2_ASAP7_75t_L g299 ( .A(n_73), .B(n_229), .Y(n_299) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_74), .A2(n_274), .B(n_275), .C(n_277), .Y(n_273) );
BUFx2_ASAP7_75t_SL g179 ( .A(n_75), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_76), .B(n_221), .Y(n_258) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_174), .B1(n_188), .B2(n_549), .C(n_550), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_164), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_80), .Y(n_163) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NAND2xp5_ASAP7_75t_L g81 ( .A(n_82), .B(n_133), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_119), .Y(n_82) );
NAND2xp5_ASAP7_75t_SL g83 ( .A(n_84), .B(n_108), .Y(n_83) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
INVx3_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_97), .Y(n_87) );
AND2x2_ASAP7_75t_L g111 ( .A(n_88), .B(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_L g157 ( .A(n_88), .B(n_105), .Y(n_157) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_92), .Y(n_88) );
INVx2_ASAP7_75t_L g107 ( .A(n_89), .Y(n_107) );
BUFx2_ASAP7_75t_L g117 ( .A(n_89), .Y(n_117) );
AND2x2_ASAP7_75t_L g138 ( .A(n_89), .B(n_93), .Y(n_138) );
INVx1_ASAP7_75t_L g91 ( .A(n_90), .Y(n_91) );
OAI22x1_ASAP7_75t_L g93 ( .A1(n_90), .A2(n_94), .B1(n_95), .B2(n_96), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_90), .Y(n_94) );
INVx2_ASAP7_75t_L g100 ( .A(n_90), .Y(n_100) );
INVx1_ASAP7_75t_L g103 ( .A(n_90), .Y(n_103) );
AND2x4_ASAP7_75t_L g106 ( .A(n_92), .B(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
AND2x2_ASAP7_75t_L g123 ( .A(n_93), .B(n_107), .Y(n_123) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_93), .Y(n_146) );
AND2x4_ASAP7_75t_L g122 ( .A(n_97), .B(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g129 ( .A(n_97), .B(n_106), .Y(n_129) );
AND2x4_ASAP7_75t_L g137 ( .A(n_97), .B(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g97 ( .A(n_98), .B(n_101), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x4_ASAP7_75t_L g105 ( .A(n_99), .B(n_101), .Y(n_105) );
INVx1_ASAP7_75t_L g113 ( .A(n_99), .Y(n_113) );
AND2x2_ASAP7_75t_L g118 ( .A(n_99), .B(n_102), .Y(n_118) );
INVxp67_ASAP7_75t_L g161 ( .A(n_101), .Y(n_161) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g112 ( .A(n_102), .B(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
AND2x2_ASAP7_75t_L g142 ( .A(n_105), .B(n_123), .Y(n_142) );
AND2x4_ASAP7_75t_L g125 ( .A(n_106), .B(n_118), .Y(n_125) );
AND2x4_ASAP7_75t_L g132 ( .A(n_106), .B(n_112), .Y(n_132) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g150 ( .A(n_112), .B(n_123), .Y(n_150) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_113), .Y(n_154) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx5_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
AND2x2_ASAP7_75t_L g145 ( .A(n_118), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_126), .Y(n_119) );
BUFx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx8_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_SL g130 ( .A(n_131), .Y(n_130) );
INVx8_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_147), .Y(n_133) );
OAI211xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B(n_139), .C(n_143), .Y(n_134) );
INVx2_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g152 ( .A(n_138), .B(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_L g160 ( .A(n_138), .B(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx12f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_155), .Y(n_147) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_SL g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx6_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_165), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B1(n_168), .B2(n_171), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_168), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_176), .Y(n_175) );
AND3x1_ASAP7_75t_SL g176 ( .A(n_177), .B(n_183), .C(n_186), .Y(n_176) );
INVxp67_ASAP7_75t_L g556 ( .A(n_177), .Y(n_556) );
CKINVDCx8_ASAP7_75t_R g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
CKINVDCx16_ASAP7_75t_R g554 ( .A(n_183), .Y(n_554) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_183), .A2(n_322), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g205 ( .A(n_184), .B(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_SL g561 ( .A(n_184), .B(n_186), .Y(n_561) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g216 ( .A(n_185), .B(n_207), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_186), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2x1p5_ASAP7_75t_L g213 ( .A(n_187), .B(n_214), .Y(n_213) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OR3x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_414), .C(n_485), .Y(n_190) );
NAND3x1_ASAP7_75t_SL g191 ( .A(n_192), .B(n_341), .C(n_363), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_331), .Y(n_192) );
AOI22xp33_ASAP7_75t_SL g193 ( .A1(n_194), .A2(n_260), .B1(n_309), .B2(n_313), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_194), .A2(n_517), .B1(n_518), .B2(n_520), .Y(n_516) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_232), .Y(n_194) );
AND2x2_ASAP7_75t_L g332 ( .A(n_195), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_195), .B(n_379), .Y(n_398) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g316 ( .A(n_196), .Y(n_316) );
AND2x2_ASAP7_75t_L g366 ( .A(n_196), .B(n_234), .Y(n_366) );
INVx1_ASAP7_75t_L g405 ( .A(n_196), .Y(n_405) );
OR2x2_ASAP7_75t_L g442 ( .A(n_196), .B(n_252), .Y(n_442) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_196), .Y(n_454) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_196), .Y(n_478) );
AND2x2_ASAP7_75t_L g535 ( .A(n_196), .B(n_362), .Y(n_535) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_202), .B(n_228), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_198), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_SL g199 ( .A(n_200), .B(n_201), .Y(n_199) );
AND2x4_ASAP7_75t_L g236 ( .A(n_200), .B(n_201), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_211), .Y(n_202) );
INVx1_ASAP7_75t_L g286 ( .A(n_204), .Y(n_286) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_208), .Y(n_204) );
INVx1_ASAP7_75t_L g322 ( .A(n_205), .Y(n_322) );
OR2x6_ASAP7_75t_L g219 ( .A(n_206), .B(n_215), .Y(n_219) );
INVxp33_ASAP7_75t_L g296 ( .A(n_206), .Y(n_296) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x4_ASAP7_75t_L g248 ( .A(n_207), .B(n_224), .Y(n_248) );
INVx1_ASAP7_75t_L g323 ( .A(n_208), .Y(n_323) );
BUFx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g215 ( .A(n_210), .Y(n_215) );
AND2x6_ASAP7_75t_L g245 ( .A(n_210), .B(n_222), .Y(n_245) );
INVxp67_ASAP7_75t_L g284 ( .A(n_212), .Y(n_284) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_212), .Y(n_549) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_216), .Y(n_212) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_213), .Y(n_564) );
INVx1_ASAP7_75t_L g297 ( .A(n_214), .Y(n_297) );
INVx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_SL g217 ( .A1(n_218), .A2(n_219), .B(n_220), .C(n_226), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_219), .A2(n_239), .B1(n_240), .B2(n_241), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_219), .A2(n_226), .B(n_257), .C(n_258), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_SL g266 ( .A1(n_219), .A2(n_226), .B(n_267), .C(n_268), .Y(n_266) );
INVxp67_ASAP7_75t_L g274 ( .A(n_219), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g305 ( .A1(n_219), .A2(n_226), .B(n_306), .C(n_307), .Y(n_305) );
INVx2_ASAP7_75t_L g329 ( .A(n_219), .Y(n_329) );
INVx1_ASAP7_75t_L g241 ( .A(n_221), .Y(n_241) );
AND2x4_ASAP7_75t_L g221 ( .A(n_222), .B(n_224), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_226), .B(n_236), .Y(n_249) );
INVx1_ASAP7_75t_L g293 ( .A(n_226), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_226), .A2(n_327), .B(n_328), .Y(n_326) );
INVx5_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_227), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_229), .A2(n_273), .B1(n_278), .B2(n_279), .Y(n_272) );
INVx3_ASAP7_75t_L g279 ( .A(n_229), .Y(n_279) );
INVx4_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_230), .B(n_282), .Y(n_281) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
BUFx4f_ASAP7_75t_L g264 ( .A(n_231), .Y(n_264) );
NOR2x1_ASAP7_75t_L g232 ( .A(n_233), .B(n_250), .Y(n_232) );
INVx1_ASAP7_75t_L g410 ( .A(n_233), .Y(n_410) );
AND2x2_ASAP7_75t_L g436 ( .A(n_233), .B(n_252), .Y(n_436) );
NAND2x1_ASAP7_75t_L g452 ( .A(n_233), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g333 ( .A(n_234), .B(n_319), .Y(n_333) );
INVx3_ASAP7_75t_L g362 ( .A(n_234), .Y(n_362) );
NOR2x1_ASAP7_75t_SL g481 ( .A(n_234), .B(n_252), .Y(n_481) );
AND2x4_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_236), .A2(n_255), .B(n_259), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_242), .B(n_249), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_241), .B(n_276), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B1(n_246), .B2(n_247), .Y(n_242) );
INVxp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OAI222xp33_ASAP7_75t_L g550 ( .A1(n_246), .A2(n_551), .B1(n_552), .B2(n_557), .C1(n_559), .C2(n_562), .Y(n_550) );
INVxp67_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_250), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g360 ( .A(n_251), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx4_ASAP7_75t_L g330 ( .A(n_252), .Y(n_330) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_252), .Y(n_375) );
AND2x2_ASAP7_75t_L g447 ( .A(n_252), .B(n_319), .Y(n_447) );
AND2x4_ASAP7_75t_L g464 ( .A(n_252), .B(n_408), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_252), .B(n_406), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_252), .B(n_315), .Y(n_540) );
OR2x6_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_260), .A2(n_357), .B1(n_428), .B2(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_287), .Y(n_260) );
INVx2_ASAP7_75t_L g430 ( .A(n_261), .Y(n_430) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_270), .Y(n_261) );
BUFx3_ASAP7_75t_L g420 ( .A(n_262), .Y(n_420) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_263), .B(n_289), .Y(n_312) );
INVx2_ASAP7_75t_L g336 ( .A(n_263), .Y(n_336) );
INVx1_ASAP7_75t_L g348 ( .A(n_263), .Y(n_348) );
AND2x4_ASAP7_75t_L g355 ( .A(n_263), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g372 ( .A(n_263), .B(n_271), .Y(n_372) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_263), .Y(n_386) );
INVxp67_ASAP7_75t_L g394 ( .A(n_263), .Y(n_394) );
OA21x2_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_265), .B(n_269), .Y(n_263) );
INVx2_ASAP7_75t_SL g290 ( .A(n_264), .Y(n_290) );
AND2x2_ASAP7_75t_L g423 ( .A(n_270), .B(n_339), .Y(n_423) );
AND2x2_ASAP7_75t_L g439 ( .A(n_270), .B(n_340), .Y(n_439) );
NOR2xp67_ASAP7_75t_L g526 ( .A(n_270), .B(n_339), .Y(n_526) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x4_ASAP7_75t_L g335 ( .A(n_271), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g346 ( .A(n_271), .Y(n_346) );
INVx1_ASAP7_75t_L g359 ( .A(n_271), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_271), .B(n_301), .Y(n_396) );
OR2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_280), .Y(n_271) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_279), .A2(n_302), .B(n_308), .Y(n_301) );
AO21x2_ASAP7_75t_L g339 ( .A1(n_279), .A2(n_302), .B(n_308), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_284), .B1(n_285), .B2(n_286), .Y(n_280) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g519 ( .A(n_287), .Y(n_519) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_300), .Y(n_287) );
AND2x2_ASAP7_75t_L g393 ( .A(n_288), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g422 ( .A(n_288), .Y(n_422) );
AND2x2_ASAP7_75t_L g524 ( .A(n_288), .B(n_339), .Y(n_524) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_289), .B(n_301), .Y(n_384) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B(n_299), .Y(n_289) );
AO21x2_ASAP7_75t_L g340 ( .A1(n_290), .A2(n_291), .B(n_299), .Y(n_340) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_292), .B(n_298), .Y(n_291) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx3_ASAP7_75t_L g310 ( .A(n_300), .Y(n_310) );
NAND2x1p5_ASAP7_75t_L g499 ( .A(n_300), .B(n_420), .Y(n_499) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_301), .Y(n_413) );
AND2x2_ASAP7_75t_L g440 ( .A(n_301), .B(n_386), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AND2x2_ASAP7_75t_L g354 ( .A(n_310), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g370 ( .A(n_310), .Y(n_370) );
AND2x2_ASAP7_75t_L g458 ( .A(n_310), .B(n_335), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_310), .B(n_478), .Y(n_483) );
AND2x2_ASAP7_75t_L g493 ( .A(n_310), .B(n_372), .Y(n_493) );
OR2x2_ASAP7_75t_L g530 ( .A(n_310), .B(n_430), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_311), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g490 ( .A(n_311), .B(n_346), .Y(n_490) );
AND2x2_ASAP7_75t_L g506 ( .A(n_311), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g500 ( .A(n_312), .B(n_396), .Y(n_500) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_317), .Y(n_313) );
INVx1_ASAP7_75t_L g382 ( .A(n_314), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_314), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g480 ( .A(n_314), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_314), .B(n_361), .Y(n_505) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_315), .Y(n_352) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_316), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_317), .A2(n_350), .B1(n_368), .B2(n_371), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_317), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_SL g484 ( .A(n_317), .Y(n_484) );
AND2x4_ASAP7_75t_SL g317 ( .A(n_318), .B(n_330), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g361 ( .A(n_319), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g381 ( .A(n_319), .Y(n_381) );
INVx1_ASAP7_75t_L g408 ( .A(n_319), .Y(n_408) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_325), .Y(n_319) );
NOR3xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .C(n_324), .Y(n_321) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_330), .Y(n_350) );
AND2x4_ASAP7_75t_L g407 ( .A(n_330), .B(n_408), .Y(n_407) );
NOR2x1_ASAP7_75t_L g468 ( .A(n_330), .B(n_437), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
AND2x2_ASAP7_75t_L g432 ( .A(n_332), .B(n_375), .Y(n_432) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_332), .A2(n_513), .B(n_514), .Y(n_512) );
INVx2_ASAP7_75t_L g390 ( .A(n_333), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_334), .A2(n_444), .B1(n_448), .B2(n_451), .Y(n_443) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_335), .Y(n_401) );
AND2x2_ASAP7_75t_L g411 ( .A(n_335), .B(n_412), .Y(n_411) );
INVx3_ASAP7_75t_L g450 ( .A(n_335), .Y(n_450) );
NAND2x1_ASAP7_75t_SL g475 ( .A(n_335), .B(n_344), .Y(n_475) );
AND2x2_ASAP7_75t_L g371 ( .A(n_337), .B(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NOR2x1_ASAP7_75t_L g347 ( .A(n_339), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g344 ( .A(n_340), .Y(n_344) );
INVx2_ASAP7_75t_L g356 ( .A(n_340), .Y(n_356) );
AOI21xp5_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_349), .B(n_353), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_344), .B(n_538), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_345), .A2(n_434), .B1(n_438), .B2(n_441), .Y(n_433) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
BUFx2_ASAP7_75t_L g538 ( .A(n_346), .Y(n_538) );
INVx1_ASAP7_75t_SL g545 ( .A(n_346), .Y(n_545) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_347), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OA21x2_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_357), .B(n_360), .Y(n_353) );
AND2x2_ASAP7_75t_L g357 ( .A(n_355), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g399 ( .A(n_355), .B(n_395), .Y(n_399) );
AND2x2_ASAP7_75t_L g514 ( .A(n_355), .B(n_412), .Y(n_514) );
AND2x2_ASAP7_75t_L g517 ( .A(n_355), .B(n_423), .Y(n_517) );
AND2x4_ASAP7_75t_L g525 ( .A(n_355), .B(n_526), .Y(n_525) );
OAI21xp33_ASAP7_75t_L g479 ( .A1(n_357), .A2(n_480), .B(n_482), .Y(n_479) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g507 ( .A(n_359), .Y(n_507) );
AND2x2_ASAP7_75t_L g523 ( .A(n_359), .B(n_524), .Y(n_523) );
INVx4_ASAP7_75t_L g437 ( .A(n_361), .Y(n_437) );
INVx1_ASAP7_75t_L g406 ( .A(n_362), .Y(n_406) );
AND2x2_ASAP7_75t_L g428 ( .A(n_362), .B(n_381), .Y(n_428) );
NOR2x1_ASAP7_75t_L g363 ( .A(n_364), .B(n_387), .Y(n_363) );
OAI21xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_367), .B(n_373), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g374 ( .A(n_366), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_SL g527 ( .A(n_366), .B(n_379), .Y(n_527) );
AND2x2_ASAP7_75t_L g548 ( .A(n_366), .B(n_464), .Y(n_548) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g474 ( .A(n_371), .Y(n_474) );
OAI21xp5_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_376), .B(n_383), .Y(n_373) );
OR2x6_ASAP7_75t_L g426 ( .A(n_375), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_382), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
OR2x2_ASAP7_75t_L g449 ( .A(n_384), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g546 ( .A(n_384), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_385), .B(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_400), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B1(n_397), .B2(n_399), .Y(n_388) );
OR2x2_ASAP7_75t_L g460 ( .A(n_390), .B(n_461), .Y(n_460) );
INVx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_392), .Y(n_417) );
NAND2x1p5_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
INVx1_ASAP7_75t_L g466 ( .A(n_395), .Y(n_466) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_409), .B2(n_411), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_407), .Y(n_403) );
AND2x4_ASAP7_75t_SL g404 ( .A(n_405), .B(n_406), .Y(n_404) );
AND2x2_ASAP7_75t_L g409 ( .A(n_407), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g470 ( .A(n_410), .B(n_464), .Y(n_470) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_415), .B(n_455), .Y(n_414) );
NOR2xp67_ASAP7_75t_L g415 ( .A(n_416), .B(n_429), .Y(n_415) );
AOI21xp33_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_418), .B(n_424), .Y(n_416) );
OR2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND2x1p5_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI22xp33_ASAP7_75t_SL g494 ( .A1(n_426), .A2(n_495), .B1(n_497), .B2(n_500), .Y(n_494) );
NOR2x1_ASAP7_75t_L g441 ( .A(n_427), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g477 ( .A(n_428), .B(n_478), .Y(n_477) );
OAI211xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_431), .B(n_433), .C(n_443), .Y(n_429) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2xp33_ASAP7_75t_SL g434 ( .A(n_435), .B(n_437), .Y(n_434) );
INVxp33_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g446 ( .A(n_437), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g457 ( .A1(n_438), .A2(n_458), .B1(n_459), .B2(n_462), .C(n_465), .Y(n_457) );
AND2x4_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g498 ( .A(n_439), .Y(n_498) );
INVx2_ASAP7_75t_SL g496 ( .A(n_442), .Y(n_496) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
NAND2x1_ASAP7_75t_L g495 ( .A(n_446), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g492 ( .A(n_452), .Y(n_492) );
INVx1_ASAP7_75t_L g521 ( .A(n_453), .Y(n_521) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NOR2x1_ASAP7_75t_L g455 ( .A(n_456), .B(n_471), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_469), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g510 ( .A(n_461), .Y(n_510) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g531 ( .A(n_464), .B(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g536 ( .A(n_464), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVxp33_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g489 ( .A(n_468), .Y(n_489) );
OAI21xp5_ASAP7_75t_SL g471 ( .A1(n_472), .A2(n_476), .B(n_479), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_L g532 ( .A(n_478), .Y(n_532) );
AND2x2_ASAP7_75t_L g520 ( .A(n_481), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_R g482 ( .A(n_483), .B(n_484), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_501), .C(n_528), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_494), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_488), .B(n_491), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
OR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_515), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_503), .B(n_512), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g503 ( .A1(n_504), .A2(n_506), .B1(n_508), .B2(n_509), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NOR2x1_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
INVxp67_ASAP7_75t_SL g513 ( .A(n_511), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_516), .B(n_522), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_525), .B(n_527), .Y(n_522) );
INVx1_ASAP7_75t_L g541 ( .A(n_525), .Y(n_541) );
AOI211xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_531), .B(n_533), .C(n_542), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_537), .B1(n_539), .B2(n_541), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_547), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
INVxp67_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_563), .Y(n_562) );
endmodule