module fake_jpeg_9085_n_108 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx4f_ASAP7_75t_SL g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx4f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

AOI21xp33_ASAP7_75t_L g22 ( 
.A1(n_20),
.A2(n_0),
.B(n_1),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_26),
.B1(n_15),
.B2(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_11),
.B(n_0),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_14),
.C(n_18),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_32),
.Y(n_42)
);

BUFx2_ASAP7_75t_SL g41 ( 
.A(n_29),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_15),
.B1(n_18),
.B2(n_14),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_25),
.B1(n_13),
.B2(n_20),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_23),
.C(n_26),
.Y(n_32)
);

INVx2_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_27),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_44),
.B1(n_17),
.B2(n_2),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_13),
.B(n_19),
.C(n_16),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_33),
.B(n_32),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_17),
.B(n_12),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_23),
.B(n_21),
.C(n_10),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_19),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_25),
.B1(n_21),
.B2(n_23),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_10),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_57),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_1),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_70),
.B1(n_55),
.B2(n_51),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_42),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_69),
.C(n_53),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_39),
.B(n_50),
.C(n_46),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_74),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_40),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_54),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_79),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_76),
.B(n_53),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_56),
.C(n_43),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_45),
.B(n_68),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_61),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_85),
.C(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_60),
.Y(n_84)
);

BUFx24_ASAP7_75t_SL g87 ( 
.A(n_84),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_85),
.C(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_89),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_72),
.B(n_77),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_91),
.B(n_62),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_83),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_64),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_94),
.Y(n_97)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_96),
.A2(n_75),
.B1(n_63),
.B2(n_47),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_99),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_74),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_95),
.Y(n_101)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_96),
.A3(n_8),
.B1(n_6),
.B2(n_7),
.C1(n_5),
.C2(n_3),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_92),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_103),
.B(n_7),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_74),
.C(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_106),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_104),
.Y(n_108)
);


endmodule