module fake_jpeg_3577_n_683 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_683);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_683;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_19),
.B(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_14),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_59),
.Y(n_158)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_61),
.B(n_62),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_64),
.B(n_66),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_65),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_20),
.B(n_56),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_67),
.B(n_95),
.C(n_98),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_68),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_10),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_69),
.B(n_75),
.Y(n_190)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g138 ( 
.A(n_70),
.Y(n_138)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_71),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_47),
.B(n_10),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_73),
.B(n_76),
.Y(n_133)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_32),
.B(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_21),
.B(n_10),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_25),
.B(n_11),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_77),
.B(n_84),
.Y(n_171)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_78),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g172 ( 
.A(n_79),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_80),
.B(n_82),
.Y(n_191)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_26),
.B(n_11),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_26),
.B(n_11),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_86),
.B(n_87),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_30),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g88 ( 
.A(n_22),
.Y(n_88)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_89),
.Y(n_177)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_37),
.Y(n_90)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_91),
.Y(n_173)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_92),
.Y(n_176)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_93),
.Y(n_144)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_1),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_96),
.Y(n_184)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_97),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_1),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_99),
.Y(n_193)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_30),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_102),
.B(n_104),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_103),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_30),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_106),
.Y(n_231)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_108),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_109),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_48),
.B(n_12),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_110),
.B(n_112),
.Y(n_227)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_34),
.Y(n_111)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_111),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_50),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_2),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_113),
.B(n_130),
.C(n_3),
.Y(n_216)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_114),
.Y(n_217)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_115),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_46),
.B(n_2),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_116),
.B(n_118),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_46),
.B(n_2),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_23),
.Y(n_119)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_119),
.Y(n_223)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_23),
.Y(n_123)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_123),
.Y(n_230)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_126),
.Y(n_197)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_44),
.Y(n_127)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_127),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_128),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_51),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_129),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_51),
.B(n_2),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_29),
.Y(n_131)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_131),
.Y(n_209)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_36),
.Y(n_132)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_80),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_135),
.B(n_113),
.Y(n_234)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_137),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_52),
.B1(n_38),
.B2(n_35),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_139),
.A2(n_157),
.B1(n_138),
.B2(n_168),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_36),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_142),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_29),
.B1(n_49),
.B2(n_35),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_147),
.B(n_207),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_38),
.B1(n_49),
.B2(n_41),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_155),
.A2(n_178),
.B1(n_179),
.B2(n_188),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_67),
.A2(n_29),
.B1(n_49),
.B2(n_35),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_94),
.A2(n_42),
.B1(n_41),
.B2(n_38),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g294 ( 
.A1(n_168),
.A2(n_175),
.B1(n_185),
.B2(n_195),
.Y(n_294)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_63),
.Y(n_170)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_170),
.Y(n_245)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_81),
.Y(n_174)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_174),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_97),
.A2(n_42),
.B1(n_127),
.B2(n_106),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_67),
.A2(n_41),
.B1(n_53),
.B2(n_32),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_71),
.A2(n_99),
.B1(n_89),
.B2(n_128),
.Y(n_179)
);

INVx6_ASAP7_75t_SL g180 ( 
.A(n_60),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_180),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_114),
.A2(n_54),
.B1(n_27),
.B2(n_28),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_85),
.Y(n_186)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_186),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_65),
.A2(n_43),
.B1(n_54),
.B2(n_27),
.Y(n_188)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_194),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_70),
.A2(n_28),
.B1(n_39),
.B2(n_53),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_93),
.A2(n_28),
.B1(n_44),
.B2(n_43),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_196),
.A2(n_199),
.B1(n_203),
.B2(n_206),
.Y(n_302)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_198),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_72),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_120),
.Y(n_200)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_200),
.Y(n_295)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_201),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_59),
.A2(n_12),
.B1(n_17),
.B2(n_5),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_90),
.Y(n_204)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_204),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_78),
.A2(n_12),
.B1(n_17),
.B2(n_5),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_103),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_207),
.A2(n_215),
.B1(n_199),
.B2(n_195),
.Y(n_255)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_129),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_68),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_214),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_117),
.A2(n_125),
.B1(n_109),
.B2(n_88),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_216),
.B(n_208),
.Y(n_282)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_88),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_218),
.Y(n_292)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_79),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_219),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_95),
.B(n_13),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_220),
.B(n_98),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_100),
.A2(n_13),
.B1(n_16),
.B2(n_7),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_221),
.A2(n_126),
.B1(n_122),
.B2(n_121),
.Y(n_243)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_131),
.Y(n_226)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_105),
.Y(n_228)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_95),
.A2(n_9),
.B(n_16),
.C(n_7),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_113),
.B(n_98),
.C(n_8),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g324 ( 
.A1(n_232),
.A2(n_266),
.B(n_272),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_152),
.Y(n_233)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_233),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_234),
.B(n_282),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_235),
.B(n_248),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_146),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_237),
.B(n_251),
.Y(n_348)
);

INVx2_ASAP7_75t_R g238 ( 
.A(n_142),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_238),
.Y(n_320)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_141),
.Y(n_239)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_239),
.Y(n_373)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_158),
.Y(n_240)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_240),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_188),
.A2(n_184),
.B1(n_230),
.B2(n_223),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_242),
.A2(n_291),
.B1(n_224),
.B2(n_172),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_243),
.A2(n_265),
.B1(n_267),
.B2(n_271),
.Y(n_358)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_152),
.Y(n_246)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_246),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_111),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_220),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_249),
.B(n_253),
.Y(n_319)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_148),
.Y(n_250)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_250),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_187),
.B(n_8),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_189),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_255),
.A2(n_278),
.B1(n_172),
.B2(n_298),
.Y(n_332)
);

A2O1A1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_171),
.A2(n_229),
.B(n_133),
.C(n_227),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_L g351 ( 
.A1(n_256),
.A2(n_298),
.B(n_294),
.C(n_315),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_151),
.B(n_3),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_257),
.B(n_260),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_161),
.B(n_211),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_212),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_261),
.B(n_268),
.Y(n_357)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_181),
.Y(n_262)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_262),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_181),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_264),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_191),
.A2(n_8),
.B1(n_9),
.B2(n_14),
.Y(n_265)
);

OAI21xp33_ASAP7_75t_L g266 ( 
.A1(n_190),
.A2(n_9),
.B(n_14),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_217),
.A2(n_15),
.B1(n_18),
.B2(n_4),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_136),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_169),
.Y(n_269)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_269),
.Y(n_343)
);

INVx8_ASAP7_75t_L g270 ( 
.A(n_160),
.Y(n_270)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_270),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_217),
.A2(n_18),
.B1(n_205),
.B2(n_167),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_173),
.B(n_192),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_274),
.B(n_277),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_209),
.Y(n_275)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_275),
.Y(n_333)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_149),
.Y(n_276)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_276),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_176),
.B(n_143),
.Y(n_277)
);

INVx11_ASAP7_75t_L g279 ( 
.A(n_137),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_279),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_209),
.Y(n_280)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_280),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_160),
.Y(n_281)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_281),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_177),
.Y(n_283)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_283),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_177),
.Y(n_284)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_284),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_226),
.Y(n_285)
);

INVx13_ASAP7_75t_L g326 ( 
.A(n_285),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_231),
.A2(n_144),
.B1(n_138),
.B2(n_208),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_286),
.A2(n_300),
.B1(n_306),
.B2(n_312),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_140),
.B(n_145),
.C(n_162),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g341 ( 
.A(n_287),
.B(n_238),
.CI(n_260),
.CON(n_341),
.SN(n_341)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_150),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_288),
.B(n_293),
.Y(n_369)
);

INVx5_ASAP7_75t_SL g290 ( 
.A(n_148),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_290),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_159),
.A2(n_166),
.B1(n_164),
.B2(n_193),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_219),
.B(n_144),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_L g298 ( 
.A1(n_185),
.A2(n_196),
.B(n_221),
.C(n_206),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_159),
.B(n_134),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_299),
.B(n_313),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_156),
.A2(n_175),
.B1(n_222),
.B2(n_158),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_215),
.B(n_203),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_301),
.B(n_303),
.Y(n_345)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_165),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_222),
.B(n_156),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_304),
.B(n_310),
.Y(n_354)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_163),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_305),
.Y(n_330)
);

BUFx12f_ASAP7_75t_L g306 ( 
.A(n_172),
.Y(n_306)
);

INVx6_ASAP7_75t_L g308 ( 
.A(n_193),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_308),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_183),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_309),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_154),
.B(n_182),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_154),
.B(n_182),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_311),
.B(n_315),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_165),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_134),
.B(n_153),
.Y(n_313)
);

AND2x2_ASAP7_75t_SL g314 ( 
.A(n_197),
.B(n_225),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_314),
.B(n_296),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_197),
.B(n_153),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_224),
.B(n_225),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_317),
.B(n_239),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_272),
.A2(n_278),
.B1(n_282),
.B2(n_297),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_325),
.A2(n_332),
.B1(n_335),
.B2(n_363),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g424 ( 
.A(n_328),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_247),
.A2(n_302),
.B1(n_301),
.B2(n_274),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_331),
.A2(n_340),
.B1(n_350),
.B2(n_362),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_282),
.A2(n_253),
.B1(n_257),
.B2(n_300),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g338 ( 
.A1(n_294),
.A2(n_232),
.B(n_277),
.Y(n_338)
);

O2A1O1Ixp33_ASAP7_75t_L g429 ( 
.A1(n_338),
.A2(n_327),
.B(n_353),
.C(n_323),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_299),
.A2(n_313),
.B1(n_249),
.B2(n_256),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_341),
.B(n_250),
.C(n_306),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_241),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_346),
.B(n_371),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_294),
.A2(n_269),
.B1(n_288),
.B2(n_244),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_351),
.B(n_359),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_294),
.A2(n_315),
.B1(n_305),
.B2(n_303),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_352),
.A2(n_252),
.B(n_292),
.Y(n_388)
);

A2O1A1Ixp33_ASAP7_75t_L g359 ( 
.A1(n_287),
.A2(n_254),
.B(n_259),
.C(n_245),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_291),
.A2(n_314),
.B1(n_254),
.B2(n_259),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_314),
.A2(n_308),
.B1(n_246),
.B2(n_244),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_262),
.A2(n_273),
.B1(n_289),
.B2(n_295),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_364),
.A2(n_367),
.B1(n_368),
.B2(n_372),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_366),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_245),
.A2(n_307),
.B1(n_295),
.B2(n_289),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_273),
.A2(n_307),
.B1(n_276),
.B2(n_316),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_316),
.B(n_236),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_370),
.B(n_379),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_241),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_270),
.A2(n_233),
.B1(n_284),
.B2(n_283),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_292),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_377),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_236),
.B(n_263),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_281),
.A2(n_312),
.B1(n_240),
.B2(n_263),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_380),
.A2(n_327),
.B1(n_328),
.B2(n_323),
.Y(n_416)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_321),
.Y(n_381)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_381),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_336),
.Y(n_383)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_383),
.Y(n_454)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_321),
.Y(n_385)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_385),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_370),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_386),
.B(n_394),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_388),
.A2(n_395),
.B(n_419),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_319),
.B(n_252),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_389),
.B(n_411),
.C(n_417),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_361),
.B(n_280),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_392),
.B(n_396),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_357),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_325),
.A2(n_275),
.B1(n_285),
.B2(n_290),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_361),
.B(n_258),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_329),
.B(n_258),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_397),
.B(n_403),
.Y(n_443)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_379),
.Y(n_398)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_398),
.Y(n_445)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_344),
.Y(n_399)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_399),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_368),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_400),
.B(n_410),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_351),
.A2(n_345),
.B(n_335),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_401),
.A2(n_373),
.B(n_347),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_322),
.B(n_348),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_402),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_319),
.B(n_250),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_349),
.Y(n_404)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_404),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_405),
.B(n_389),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_329),
.B(n_306),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_406),
.B(n_408),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_332),
.A2(n_279),
.B1(n_306),
.B2(n_345),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_344),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_409),
.Y(n_449)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_318),
.B(n_340),
.C(n_337),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_349),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_412),
.B(n_415),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_337),
.B(n_338),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_413),
.B(n_414),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_352),
.A2(n_338),
.B1(n_318),
.B2(n_341),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_342),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g450 ( 
.A(n_416),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_322),
.B(n_354),
.Y(n_417)
);

NOR2x1p5_ASAP7_75t_L g419 ( 
.A(n_362),
.B(n_338),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_341),
.A2(n_374),
.B1(n_366),
.B2(n_354),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_SL g433 ( 
.A1(n_420),
.A2(n_421),
.B1(n_423),
.B2(n_414),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_374),
.A2(n_377),
.B1(n_358),
.B2(n_365),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_343),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_422),
.B(n_425),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_324),
.A2(n_369),
.B1(n_320),
.B2(n_339),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_339),
.B(n_369),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_375),
.B(n_342),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_426),
.B(n_394),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_363),
.A2(n_330),
.B1(n_380),
.B2(n_334),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_427),
.A2(n_430),
.B(n_367),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_359),
.B(n_346),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_428),
.B(n_376),
.Y(n_457)
);

AOI21xp33_ASAP7_75t_L g455 ( 
.A1(n_429),
.A2(n_333),
.B(n_353),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_371),
.A2(n_330),
.B(n_334),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_407),
.A2(n_424),
.B1(n_413),
.B2(n_428),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_432),
.A2(n_465),
.B1(n_416),
.B2(n_418),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_433),
.A2(n_435),
.B(n_440),
.Y(n_481)
);

XOR2x2_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_347),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_SL g489 ( 
.A(n_437),
.B(n_423),
.C(n_419),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_356),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_441),
.B(n_456),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_425),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_444),
.B(n_453),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_390),
.A2(n_355),
.B(n_373),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_446),
.A2(n_463),
.B(n_388),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_SL g448 ( 
.A1(n_421),
.A2(n_376),
.B1(n_333),
.B2(n_356),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_SL g484 ( 
.A1(n_448),
.A2(n_467),
.B1(n_391),
.B2(n_387),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_451),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_382),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_455),
.B(n_460),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_420),
.B(n_360),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_457),
.B(n_470),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_417),
.B(n_360),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_390),
.A2(n_355),
.B(n_326),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_407),
.A2(n_372),
.B1(n_378),
.B2(n_336),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_SL g467 ( 
.A1(n_408),
.A2(n_326),
.B1(n_378),
.B2(n_387),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_382),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_468),
.B(n_444),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_386),
.B(n_326),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_469),
.B(n_471),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_398),
.B(n_392),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_406),
.B(n_405),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_472),
.B(n_418),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_433),
.A2(n_395),
.B1(n_419),
.B2(n_400),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_473),
.A2(n_479),
.B1(n_488),
.B2(n_510),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_469),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_474),
.B(n_475),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_439),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_434),
.Y(n_476)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_476),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_439),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_478),
.B(n_483),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_453),
.A2(n_419),
.B1(n_396),
.B2(n_427),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_434),
.Y(n_480)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_480),
.Y(n_535)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_438),
.Y(n_482)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_482),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_484),
.Y(n_536)
);

CKINVDCx14_ASAP7_75t_R g487 ( 
.A(n_436),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_487),
.Y(n_522)
);

XNOR2x1_ASAP7_75t_L g529 ( 
.A(n_489),
.B(n_437),
.Y(n_529)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_438),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_492),
.B(n_494),
.Y(n_514)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_442),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_464),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_495),
.B(n_501),
.Y(n_516)
);

CKINVDCx14_ASAP7_75t_R g496 ( 
.A(n_436),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_496),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_432),
.A2(n_397),
.B1(n_429),
.B2(n_384),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_497),
.A2(n_445),
.B1(n_431),
.B2(n_467),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_450),
.A2(n_435),
.B1(n_468),
.B2(n_458),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_498),
.A2(n_503),
.B1(n_511),
.B2(n_431),
.Y(n_533)
);

CKINVDCx14_ASAP7_75t_R g499 ( 
.A(n_442),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_499),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_500),
.B(n_461),
.Y(n_523)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_464),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_454),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_502),
.B(n_505),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_450),
.A2(n_429),
.B1(n_403),
.B2(n_393),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_504),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_470),
.B(n_452),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_471),
.B(n_393),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_506),
.Y(n_546)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_449),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_507),
.B(n_509),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_447),
.A2(n_430),
.B(n_415),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_508),
.A2(n_457),
.B(n_440),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_443),
.B(n_445),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_459),
.A2(n_381),
.B1(n_385),
.B2(n_422),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_458),
.A2(n_391),
.B1(n_399),
.B2(n_409),
.Y(n_511)
);

XOR2x2_ASAP7_75t_L g512 ( 
.A(n_486),
.B(n_459),
.Y(n_512)
);

XNOR2x1_ASAP7_75t_L g552 ( 
.A(n_512),
.B(n_529),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_486),
.B(n_472),
.Y(n_513)
);

MAJx2_ASAP7_75t_L g553 ( 
.A(n_513),
.B(n_531),
.C(n_541),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_490),
.B(n_451),
.C(n_441),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_519),
.B(n_524),
.C(n_525),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_521),
.A2(n_483),
.B(n_481),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_SL g559 ( 
.A(n_523),
.B(n_524),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_477),
.B(n_472),
.C(n_461),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_477),
.B(n_460),
.C(n_456),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_527),
.A2(n_549),
.B1(n_479),
.B2(n_507),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_485),
.Y(n_530)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_530),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_500),
.B(n_456),
.Y(n_531)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_533),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_508),
.A2(n_455),
.B(n_437),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_534),
.A2(n_503),
.B(n_496),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_475),
.B(n_443),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g563 ( 
.A(n_537),
.B(n_485),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_488),
.A2(n_465),
.B1(n_446),
.B2(n_463),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_538),
.A2(n_544),
.B1(n_484),
.B2(n_498),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_477),
.B(n_447),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_506),
.B(n_462),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_542),
.B(n_545),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_473),
.A2(n_448),
.B1(n_462),
.B2(n_449),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_510),
.B(n_449),
.C(n_410),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_478),
.B(n_466),
.C(n_404),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_547),
.B(n_511),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_499),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_548),
.B(n_494),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_498),
.A2(n_466),
.B1(n_454),
.B2(n_383),
.Y(n_549)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_550),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_530),
.B(n_505),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_554),
.B(n_560),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_543),
.B(n_493),
.Y(n_555)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_555),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_556),
.A2(n_575),
.B(n_534),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_557),
.A2(n_564),
.B1(n_527),
.B2(n_521),
.Y(n_591)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_517),
.Y(n_558)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_558),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_SL g586 ( 
.A(n_559),
.B(n_565),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_523),
.B(n_509),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_517),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_SL g604 ( 
.A(n_561),
.B(n_566),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_563),
.A2(n_569),
.B1(n_576),
.B2(n_579),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_515),
.A2(n_497),
.B1(n_504),
.B2(n_493),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_SL g565 ( 
.A(n_541),
.B(n_481),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_526),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_516),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_567),
.Y(n_594)
);

BUFx24_ASAP7_75t_SL g568 ( 
.A(n_546),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_568),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_SL g570 ( 
.A(n_531),
.B(n_491),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_SL g602 ( 
.A(n_570),
.B(n_552),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_573),
.B(n_542),
.Y(n_601)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_514),
.Y(n_574)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_574),
.Y(n_606)
);

OAI21xp33_ASAP7_75t_L g576 ( 
.A1(n_528),
.A2(n_491),
.B(n_474),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_543),
.B(n_487),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_577),
.B(n_578),
.Y(n_590)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_518),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_519),
.B(n_482),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_520),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_580),
.B(n_581),
.Y(n_595)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_520),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_L g615 ( 
.A1(n_582),
.A2(n_592),
.B(n_532),
.Y(n_615)
);

BUFx12_ASAP7_75t_L g584 ( 
.A(n_572),
.Y(n_584)
);

CKINVDCx16_ASAP7_75t_R g619 ( 
.A(n_584),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_562),
.B(n_513),
.C(n_525),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_585),
.B(n_587),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_562),
.B(n_559),
.C(n_572),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_553),
.B(n_547),
.C(n_545),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_588),
.B(n_593),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_SL g620 ( 
.A1(n_591),
.A2(n_538),
.B1(n_522),
.B2(n_511),
.Y(n_620)
);

AOI321xp33_ASAP7_75t_L g592 ( 
.A1(n_558),
.A2(n_546),
.A3(n_548),
.B1(n_539),
.B2(n_522),
.C(n_532),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_553),
.B(n_528),
.C(n_512),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_565),
.B(n_529),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g625 ( 
.A(n_596),
.B(n_601),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_571),
.A2(n_515),
.B1(n_536),
.B2(n_539),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_598),
.A2(n_599),
.B1(n_544),
.B2(n_569),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_564),
.A2(n_557),
.B1(n_533),
.B2(n_551),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_602),
.B(n_512),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_595),
.B(n_555),
.Y(n_607)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_607),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_608),
.A2(n_620),
.B1(n_591),
.B2(n_599),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_601),
.B(n_573),
.C(n_551),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_609),
.B(n_613),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_595),
.B(n_577),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_610),
.B(n_614),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_582),
.A2(n_575),
.B(n_556),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_611),
.A2(n_612),
.B(n_615),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_SL g612 ( 
.A1(n_600),
.A2(n_550),
.B(n_489),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_588),
.B(n_570),
.C(n_552),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_590),
.Y(n_614)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_590),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_616),
.B(n_617),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_594),
.B(n_578),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_618),
.B(n_622),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_589),
.B(n_549),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_603),
.B(n_580),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_623),
.B(n_627),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_587),
.B(n_581),
.C(n_540),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_624),
.B(n_619),
.C(n_609),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_593),
.B(n_540),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_629),
.B(n_634),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_SL g654 ( 
.A1(n_630),
.A2(n_635),
.B1(n_640),
.B2(n_637),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_624),
.B(n_605),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_632),
.B(n_636),
.Y(n_649)
);

NOR2x1_ASAP7_75t_L g634 ( 
.A(n_614),
.B(n_600),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_615),
.A2(n_603),
.B1(n_597),
.B2(n_583),
.Y(n_635)
);

AO221x1_ASAP7_75t_L g636 ( 
.A1(n_627),
.A2(n_604),
.B1(n_606),
.B2(n_592),
.C(n_584),
.Y(n_636)
);

BUFx24_ASAP7_75t_SL g639 ( 
.A(n_621),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_639),
.B(n_625),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_622),
.A2(n_597),
.B1(n_606),
.B2(n_596),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_626),
.B(n_620),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_641),
.B(n_642),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_SL g642 ( 
.A1(n_611),
.A2(n_610),
.B1(n_607),
.B2(n_612),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_613),
.B(n_412),
.Y(n_643)
);

XNOR2xp5_ASAP7_75t_L g653 ( 
.A(n_643),
.B(n_535),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_629),
.B(n_585),
.C(n_625),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_647),
.B(n_650),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_SL g663 ( 
.A(n_648),
.B(n_657),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_630),
.B(n_586),
.C(n_618),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_SL g651 ( 
.A1(n_634),
.A2(n_623),
.B(n_602),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g667 ( 
.A1(n_651),
.A2(n_628),
.B(n_638),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_633),
.B(n_586),
.C(n_584),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_652),
.B(n_655),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_653),
.B(n_654),
.Y(n_666)
);

XOR2xp5_ASAP7_75t_L g655 ( 
.A(n_631),
.B(n_637),
.Y(n_655)
);

XNOR2xp5_ASAP7_75t_L g656 ( 
.A(n_631),
.B(n_535),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_656),
.B(n_659),
.Y(n_660)
);

INVx11_ASAP7_75t_L g657 ( 
.A(n_635),
.Y(n_657)
);

XNOR2xp5_ASAP7_75t_L g659 ( 
.A(n_640),
.B(n_502),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_646),
.B(n_658),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_661),
.B(n_662),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_649),
.B(n_645),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_655),
.B(n_642),
.Y(n_664)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_664),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_656),
.B(n_644),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_665),
.A2(n_650),
.B(n_659),
.Y(n_674)
);

NOR4xp25_ASAP7_75t_L g671 ( 
.A(n_667),
.B(n_628),
.C(n_657),
.D(n_651),
.Y(n_671)
);

MAJIxp5_ASAP7_75t_L g670 ( 
.A(n_668),
.B(n_647),
.C(n_652),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_670),
.A2(n_666),
.B(n_667),
.Y(n_677)
);

A2O1A1O1Ixp25_ASAP7_75t_L g678 ( 
.A1(n_671),
.A2(n_666),
.B(n_660),
.C(n_495),
.D(n_501),
.Y(n_678)
);

AOI21x1_ASAP7_75t_L g676 ( 
.A1(n_674),
.A2(n_675),
.B(n_669),
.Y(n_676)
);

NOR3xp33_ASAP7_75t_L g675 ( 
.A(n_663),
.B(n_476),
.C(n_480),
.Y(n_675)
);

XOR2xp5_ASAP7_75t_L g679 ( 
.A(n_676),
.B(n_678),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_677),
.Y(n_680)
);

MAJIxp5_ASAP7_75t_L g681 ( 
.A(n_680),
.B(n_672),
.C(n_673),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_681),
.B(n_679),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_682),
.A2(n_492),
.B(n_383),
.Y(n_683)
);


endmodule