module real_jpeg_24233_n_16 (n_5, n_4, n_8, n_0, n_12, n_353, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_353;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_2),
.A2(n_26),
.B1(n_39),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_2),
.A2(n_70),
.B1(n_79),
.B2(n_80),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_70),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_70),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

INVx8_ASAP7_75t_SL g33 ( 
.A(n_4),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_5),
.A2(n_55),
.B1(n_56),
.B2(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_5),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_5),
.A2(n_75),
.B(n_80),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_5),
.B(n_89),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_5),
.A2(n_121),
.B1(n_144),
.B2(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_5),
.A2(n_34),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_5),
.B(n_45),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_6),
.A2(n_55),
.B1(n_56),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_6),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_6),
.A2(n_79),
.B1(n_80),
.B2(n_109),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_109),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_6),
.A2(n_26),
.B1(n_39),
.B2(n_109),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_7),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_7),
.A2(n_25),
.B1(n_34),
.B2(n_35),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_7),
.A2(n_25),
.B1(n_79),
.B2(n_80),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_7),
.A2(n_25),
.B1(n_55),
.B2(n_56),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_10),
.A2(n_55),
.B1(n_56),
.B2(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_10),
.A2(n_79),
.B1(n_80),
.B2(n_118),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_118),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_10),
.A2(n_23),
.B1(n_118),
.B2(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_11),
.A2(n_79),
.B1(n_80),
.B2(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_11),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_126),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_126),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_11),
.A2(n_26),
.B1(n_126),
.B2(n_259),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_13),
.A2(n_27),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_13),
.A2(n_68),
.B1(n_79),
.B2(n_80),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_13),
.A2(n_55),
.B1(n_56),
.B2(n_68),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_68),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_43),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_14),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_14),
.A2(n_43),
.B1(n_79),
.B2(n_80),
.Y(n_128)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_15),
.Y(n_124)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_15),
.Y(n_130)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_15),
.Y(n_149)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_15),
.Y(n_278)
);

XNOR2x2_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_92),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_91),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_46),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_20),
.B(n_46),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_40),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_21),
.A2(n_30),
.B(n_66),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_22),
.B(n_45),
.Y(n_86)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_23),
.Y(n_243)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_26),
.Y(n_259)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_28),
.A2(n_45),
.B1(n_65),
.B2(n_69),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_28),
.A2(n_69),
.B(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_28),
.A2(n_45),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_28),
.A2(n_45),
.B1(n_230),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_29),
.A2(n_30),
.B1(n_242),
.B2(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_29),
.A2(n_40),
.B(n_258),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_29),
.A2(n_86),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_38),
.Y(n_29)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_30)
);

OAI32xp33_ASAP7_75t_L g210 ( 
.A1(n_31),
.A2(n_35),
.A3(n_67),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_32),
.B(n_34),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_34),
.A2(n_35),
.B1(n_54),
.B2(n_58),
.Y(n_62)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_34),
.A2(n_54),
.A3(n_56),
.B1(n_164),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_35),
.B(n_105),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_39),
.A2(n_105),
.B(n_211),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_41),
.Y(n_306)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_42),
.B(n_105),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_84),
.C(n_87),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_47),
.A2(n_48),
.B1(n_347),
.B2(n_349),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_64),
.C(n_71),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_49),
.A2(n_50),
.B1(n_71),
.B2(n_72),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_60),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_52),
.A2(n_61),
.B(n_224),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_53),
.A2(n_162),
.B1(n_165),
.B2(n_166),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_53),
.A2(n_60),
.B(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_53)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_56),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_55),
.B(n_58),
.Y(n_173)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_56),
.A2(n_77),
.B(n_105),
.C(n_111),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_59),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_59),
.A2(n_165),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_61),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_61),
.A2(n_89),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_61),
.A2(n_89),
.B1(n_188),
.B2(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_61),
.A2(n_89),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_61),
.A2(n_297),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_63),
.B(n_89),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_64),
.B(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_71),
.A2(n_72),
.B1(n_326),
.B2(n_328),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_72),
.B(n_324),
.C(n_326),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_82),
.B(n_83),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_73),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_73),
.A2(n_82),
.B1(n_108),
.B2(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_73),
.A2(n_82),
.B1(n_117),
.B2(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_73),
.A2(n_83),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_73),
.B(n_251),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_75),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_78),
.B(n_105),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_78),
.B(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_78),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_78),
.A2(n_106),
.B1(n_249),
.B2(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_79),
.B(n_151),
.Y(n_150)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_82),
.B(n_83),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_84),
.A2(n_87),
.B1(n_88),
.B2(n_348),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_84),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_345),
.B(n_351),
.Y(n_92)
);

OAI321xp33_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_320),
.A3(n_338),
.B1(n_343),
.B2(n_344),
.C(n_353),
.Y(n_93)
);

AOI311xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_273),
.A3(n_311),
.B(n_314),
.C(n_315),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_232),
.C(n_268),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_205),
.B(n_231),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_181),
.B(n_204),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_157),
.B(n_180),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_131),
.B(n_156),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_112),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_101),
.B(n_112),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_110),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_103),
.B1(n_110),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_106),
.A2(n_200),
.B(n_201),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_106),
.A2(n_266),
.B(n_281),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_120),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_119),
.C(n_120),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_125),
.B(n_127),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_130),
.B1(n_135),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_121),
.A2(n_175),
.B(n_176),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_121),
.A2(n_176),
.B(n_247),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_121),
.A2(n_175),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_122),
.B(n_177),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_122),
.A2(n_129),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_124),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_124),
.A2(n_194),
.B(n_195),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_127),
.B(n_195),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_128),
.Y(n_175)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_140),
.B(n_155),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_133),
.B(n_138),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_145),
.B(n_154),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_142),
.B(n_143),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_158),
.B(n_159),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_171),
.B1(n_178),
.B2(n_179),
.Y(n_159)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_166),
.Y(n_187)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_170),
.C(n_178),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_174),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_182),
.B(n_183),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_196),
.B2(n_197),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_199),
.C(n_202),
.Y(n_206)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_191),
.C(n_192),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_202),
.B2(n_203),
.Y(n_197)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_199),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_201),
.B(n_250),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_206),
.B(n_207),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_221),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_208)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_209),
.B(n_220),
.C(n_221),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_213),
.B1(n_216),
.B2(n_217),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_210),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_216),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_213),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_228),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_225),
.C(n_228),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_226),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_227),
.Y(n_251)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI21xp33_ASAP7_75t_L g316 ( 
.A1(n_233),
.A2(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_252),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_234),
.B(n_252),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_244),
.C(n_245),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_235),
.A2(n_236),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_239),
.C(n_240),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_244),
.B(n_245),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_248),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_252),
.Y(n_313)
);

FAx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_263),
.CI(n_267),
.CON(n_252),
.SN(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_262),
.Y(n_253)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_254),
.Y(n_262)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_260),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_257),
.B(n_260),
.C(n_262),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_261),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_265),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_269),
.B(n_270),
.Y(n_317)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

O2A1O1Ixp33_ASAP7_75t_SL g315 ( 
.A1(n_274),
.A2(n_312),
.B(n_316),
.C(n_319),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_292),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_275),
.B(n_313),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_292),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_275),
.B(n_313),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_283),
.CI(n_291),
.CON(n_275),
.SN(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_279),
.B1(n_280),
.B2(n_282),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_277),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_280),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_282),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_282),
.A2(n_301),
.B(n_305),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_290),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_287),
.C(n_288),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_286),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_289),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_310),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_300),
.B1(n_308),
.B2(n_309),
.Y(n_293)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_298),
.B(n_299),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_295),
.B(n_298),
.Y(n_299)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_299),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_299),
.A2(n_322),
.B1(n_330),
.B2(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_300),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_300),
.B(n_308),
.C(n_310),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_307),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_303),
.Y(n_307)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_332),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_321),
.B(n_332),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_330),
.C(n_331),
.Y(n_321)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_322),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_324),
.B1(n_325),
.B2(n_329),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_323),
.A2(n_324),
.B1(n_334),
.B2(n_336),
.Y(n_333)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_324),
.B(n_336),
.C(n_337),
.Y(n_350)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_325),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_326),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_337),
.Y(n_332)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_334),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_339),
.B(n_340),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_350),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_346),
.B(n_350),
.Y(n_351)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_347),
.Y(n_349)
);


endmodule