module real_aes_2311_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_0), .B(n_499), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_1), .A2(n_501), .B(n_502), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_2), .B(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g800 ( .A(n_3), .Y(n_800) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_4), .B(n_177), .Y(n_535) );
INVx1_ASAP7_75t_L g132 ( .A(n_5), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_6), .B(n_141), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_7), .B(n_177), .Y(n_523) );
INVx1_ASAP7_75t_L g187 ( .A(n_8), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g835 ( .A(n_9), .Y(n_835) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_10), .Y(n_203) );
NAND2xp33_ASAP7_75t_L g556 ( .A(n_11), .B(n_174), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_12), .A2(n_38), .B1(n_823), .B2(n_824), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_12), .Y(n_824) );
INVx2_ASAP7_75t_L g140 ( .A(n_13), .Y(n_140) );
AOI221x1_ASAP7_75t_L g580 ( .A1(n_14), .A2(n_28), .B1(n_499), .B2(n_501), .C(n_581), .Y(n_580) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_15), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_16), .B(n_499), .Y(n_552) );
INVx1_ASAP7_75t_L g175 ( .A(n_17), .Y(n_175) );
AO21x2_ASAP7_75t_L g550 ( .A1(n_18), .A2(n_163), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_19), .B(n_217), .Y(n_584) );
XOR2xp5_ASAP7_75t_L g790 ( .A(n_20), .B(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_21), .B(n_177), .Y(n_512) );
AO21x1_ASAP7_75t_L g530 ( .A1(n_22), .A2(n_499), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g115 ( .A(n_23), .Y(n_115) );
NOR2xp33_ASAP7_75t_SL g832 ( .A(n_23), .B(n_116), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_24), .A2(n_59), .B1(n_792), .B2(n_793), .Y(n_791) );
CKINVDCx16_ASAP7_75t_R g793 ( .A(n_24), .Y(n_793) );
INVx1_ASAP7_75t_L g172 ( .A(n_25), .Y(n_172) );
INVx1_ASAP7_75t_SL g247 ( .A(n_26), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_27), .B(n_152), .Y(n_151) );
AOI33xp33_ASAP7_75t_L g224 ( .A1(n_29), .A2(n_55), .A3(n_129), .B1(n_147), .B2(n_225), .B3(n_226), .Y(n_224) );
NAND2x1_ASAP7_75t_L g573 ( .A(n_30), .B(n_177), .Y(n_573) );
NAND2x1_ASAP7_75t_L g522 ( .A(n_31), .B(n_174), .Y(n_522) );
INVx1_ASAP7_75t_L g196 ( .A(n_32), .Y(n_196) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_33), .A2(n_90), .B(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g142 ( .A(n_33), .B(n_90), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_34), .B(n_185), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_35), .B(n_174), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_36), .B(n_177), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_37), .B(n_174), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_38), .Y(n_823) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_39), .A2(n_501), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g135 ( .A(n_40), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g146 ( .A(n_40), .Y(n_146) );
AND2x2_ASAP7_75t_L g161 ( .A(n_40), .B(n_132), .Y(n_161) );
OR2x6_ASAP7_75t_L g113 ( .A(n_41), .B(n_114), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g833 ( .A(n_41), .B(n_111), .C(n_834), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_42), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_43), .B(n_499), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_44), .B(n_185), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_45), .A2(n_126), .B1(n_138), .B2(n_141), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_46), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_47), .B(n_152), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_48), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_49), .B(n_174), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_50), .B(n_163), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_51), .B(n_152), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_52), .A2(n_501), .B(n_521), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_53), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_54), .B(n_174), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_56), .B(n_152), .Y(n_215) );
INVx1_ASAP7_75t_L g130 ( .A(n_57), .Y(n_130) );
INVx1_ASAP7_75t_L g154 ( .A(n_57), .Y(n_154) );
AND2x2_ASAP7_75t_L g216 ( .A(n_58), .B(n_217), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_59), .Y(n_792) );
AOI221xp5_ASAP7_75t_L g184 ( .A1(n_60), .A2(n_76), .B1(n_144), .B2(n_185), .C(n_186), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_61), .B(n_185), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_62), .B(n_177), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_63), .B(n_138), .Y(n_205) );
AOI21xp5_ASAP7_75t_SL g235 ( .A1(n_64), .A2(n_144), .B(n_236), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_65), .A2(n_501), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g168 ( .A(n_66), .Y(n_168) );
AO21x1_ASAP7_75t_L g532 ( .A1(n_67), .A2(n_501), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_68), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g214 ( .A(n_69), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_70), .B(n_499), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_71), .A2(n_144), .B(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g546 ( .A(n_72), .B(n_218), .Y(n_546) );
INVx1_ASAP7_75t_L g136 ( .A(n_73), .Y(n_136) );
INVx1_ASAP7_75t_L g156 ( .A(n_73), .Y(n_156) );
AND2x2_ASAP7_75t_L g525 ( .A(n_74), .B(n_192), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_75), .B(n_185), .Y(n_227) );
AND2x2_ASAP7_75t_L g249 ( .A(n_77), .B(n_192), .Y(n_249) );
INVx1_ASAP7_75t_L g169 ( .A(n_78), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_79), .A2(n_144), .B(n_246), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_80), .A2(n_144), .B(n_150), .C(n_162), .Y(n_143) );
INVx1_ASAP7_75t_L g116 ( .A(n_81), .Y(n_116) );
AND2x2_ASAP7_75t_L g496 ( .A(n_82), .B(n_192), .Y(n_496) );
AND2x2_ASAP7_75t_SL g233 ( .A(n_83), .B(n_192), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_84), .B(n_499), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_85), .A2(n_144), .B1(n_222), .B2(n_223), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_86), .B(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g531 ( .A(n_87), .B(n_141), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_88), .A2(n_821), .B1(n_825), .B2(n_826), .Y(n_820) );
CKINVDCx16_ASAP7_75t_R g826 ( .A(n_88), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_89), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_91), .B(n_174), .Y(n_513) );
AND2x2_ASAP7_75t_L g576 ( .A(n_92), .B(n_192), .Y(n_576) );
INVx1_ASAP7_75t_L g237 ( .A(n_93), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_94), .B(n_177), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_95), .A2(n_501), .B(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_96), .B(n_174), .Y(n_582) );
AND2x2_ASAP7_75t_L g228 ( .A(n_97), .B(n_192), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_98), .B(n_177), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_99), .A2(n_194), .B(n_195), .C(n_197), .Y(n_193) );
BUFx2_ASAP7_75t_L g812 ( .A(n_100), .Y(n_812) );
BUFx2_ASAP7_75t_SL g816 ( .A(n_100), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_101), .A2(n_501), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_102), .B(n_152), .Y(n_238) );
AOI21xp33_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_827), .B(n_836), .Y(n_103) );
AO22x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_808), .B1(n_813), .B2(n_817), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_804), .Y(n_105) );
AOI221xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_790), .B1(n_794), .B2(n_798), .C(n_799), .Y(n_106) );
OAI22xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_117), .B1(n_489), .B2(n_788), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
AOI22xp5_ASAP7_75t_L g795 ( .A1(n_109), .A2(n_117), .B1(n_489), .B2(n_796), .Y(n_795) );
CKINVDCx11_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
OR2x6_ASAP7_75t_SL g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AND2x6_ASAP7_75t_SL g789 ( .A(n_111), .B(n_113), .Y(n_789) );
OR2x2_ASAP7_75t_L g803 ( .A(n_111), .B(n_113), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_111), .B(n_112), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_423), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_346), .Y(n_118) );
NAND3xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_293), .C(n_326), .Y(n_119) );
AOI211xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_250), .B(n_259), .C(n_283), .Y(n_120) );
OAI21xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_179), .B(n_229), .Y(n_121) );
OR2x2_ASAP7_75t_L g303 ( .A(n_122), .B(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g458 ( .A(n_122), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AOI22xp33_ASAP7_75t_SL g348 ( .A1(n_123), .A2(n_349), .B1(n_353), .B2(n_355), .Y(n_348) );
AND2x2_ASAP7_75t_L g385 ( .A(n_123), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_164), .Y(n_123) );
INVx1_ASAP7_75t_L g282 ( .A(n_124), .Y(n_282) );
AND2x4_ASAP7_75t_L g299 ( .A(n_124), .B(n_280), .Y(n_299) );
INVx2_ASAP7_75t_L g321 ( .A(n_124), .Y(n_321) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_124), .Y(n_404) );
AND2x2_ASAP7_75t_L g475 ( .A(n_124), .B(n_232), .Y(n_475) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_143), .Y(n_124) );
NOR3xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_133), .C(n_137), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g185 ( .A(n_128), .B(n_134), .Y(n_185) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
OR2x6_ASAP7_75t_L g159 ( .A(n_129), .B(n_148), .Y(n_159) );
INVxp33_ASAP7_75t_L g225 ( .A(n_129), .Y(n_225) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g149 ( .A(n_130), .B(n_132), .Y(n_149) );
AND2x4_ASAP7_75t_L g177 ( .A(n_130), .B(n_155), .Y(n_177) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x6_ASAP7_75t_L g501 ( .A(n_135), .B(n_149), .Y(n_501) );
INVx2_ASAP7_75t_L g148 ( .A(n_136), .Y(n_148) );
AND2x6_ASAP7_75t_L g174 ( .A(n_136), .B(n_153), .Y(n_174) );
INVx4_ASAP7_75t_L g192 ( .A(n_138), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_138), .B(n_202), .Y(n_201) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx4f_ASAP7_75t_L g163 ( .A(n_139), .Y(n_163) );
AND2x4_ASAP7_75t_L g141 ( .A(n_140), .B(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_SL g218 ( .A(n_140), .B(n_142), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_141), .B(n_160), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_141), .A2(n_235), .B(n_239), .Y(n_234) );
INVx1_ASAP7_75t_SL g508 ( .A(n_141), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_141), .B(n_537), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_141), .A2(n_552), .B(n_553), .Y(n_551) );
INVxp67_ASAP7_75t_L g204 ( .A(n_144), .Y(n_204) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_149), .Y(n_144) );
NOR2x1p5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
INVx1_ASAP7_75t_L g226 ( .A(n_147), .Y(n_226) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_157), .B(n_160), .Y(n_150) );
INVx1_ASAP7_75t_L g170 ( .A(n_152), .Y(n_170) );
AND2x4_ASAP7_75t_L g499 ( .A(n_152), .B(n_161), .Y(n_499) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g167 ( .A1(n_159), .A2(n_168), .B1(n_169), .B2(n_170), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_SL g186 ( .A1(n_159), .A2(n_160), .B(n_187), .C(n_188), .Y(n_186) );
INVxp67_ASAP7_75t_L g194 ( .A(n_159), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_159), .A2(n_160), .B(n_214), .C(n_215), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_159), .A2(n_160), .B(n_237), .C(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_SL g246 ( .A1(n_159), .A2(n_160), .B(n_247), .C(n_248), .Y(n_246) );
INVx1_ASAP7_75t_L g222 ( .A(n_160), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_160), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_160), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_160), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_160), .A2(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_160), .A2(n_543), .B(n_544), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_160), .A2(n_555), .B(n_556), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_160), .A2(n_573), .B(n_574), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_160), .A2(n_582), .B(n_583), .Y(n_581) );
INVx5_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_161), .Y(n_197) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_162), .A2(n_220), .B(n_228), .Y(n_219) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_162), .A2(n_220), .B(n_228), .Y(n_264) );
INVx2_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
OA21x2_ASAP7_75t_L g183 ( .A1(n_163), .A2(n_184), .B(n_189), .Y(n_183) );
AND2x2_ASAP7_75t_L g240 ( .A(n_164), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g269 ( .A(n_164), .Y(n_269) );
INVx3_ASAP7_75t_L g280 ( .A(n_164), .Y(n_280) );
AND2x4_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_171), .B(n_178), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_170), .B(n_196), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B1(n_175), .B2(n_176), .Y(n_171) );
INVxp67_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVxp67_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_179), .A2(n_470), .B1(n_472), .B2(n_474), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_179), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_SL g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_207), .Y(n_180) );
INVx3_ASAP7_75t_L g253 ( .A(n_181), .Y(n_253) );
AND2x2_ASAP7_75t_L g261 ( .A(n_181), .B(n_262), .Y(n_261) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_181), .Y(n_291) );
NAND2x1_ASAP7_75t_SL g485 ( .A(n_181), .B(n_252), .Y(n_485) );
AND2x4_ASAP7_75t_L g181 ( .A(n_182), .B(n_190), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g258 ( .A(n_183), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_183), .B(n_264), .Y(n_276) );
AND2x2_ASAP7_75t_L g289 ( .A(n_183), .B(n_190), .Y(n_289) );
AND2x4_ASAP7_75t_L g296 ( .A(n_183), .B(n_297), .Y(n_296) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_183), .Y(n_345) );
INVxp67_ASAP7_75t_L g352 ( .A(n_183), .Y(n_352) );
INVx1_ASAP7_75t_L g357 ( .A(n_183), .Y(n_357) );
INVx1_ASAP7_75t_L g206 ( .A(n_185), .Y(n_206) );
INVx1_ASAP7_75t_L g256 ( .A(n_190), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_190), .B(n_266), .Y(n_275) );
INVx2_ASAP7_75t_L g343 ( .A(n_190), .Y(n_343) );
INVx1_ASAP7_75t_L g382 ( .A(n_190), .Y(n_382) );
OR2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_200), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B1(n_198), .B2(n_199), .Y(n_191) );
INVx3_ASAP7_75t_L g199 ( .A(n_192), .Y(n_199) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_199), .A2(n_210), .B(n_216), .Y(n_209) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_199), .A2(n_210), .B(n_216), .Y(n_266) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_199), .A2(n_540), .B(n_546), .Y(n_539) );
AO21x2_ASAP7_75t_L g561 ( .A1(n_199), .A2(n_540), .B(n_546), .Y(n_561) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_199), .A2(n_570), .B(n_576), .Y(n_569) );
AO21x2_ASAP7_75t_L g594 ( .A1(n_199), .A2(n_570), .B(n_576), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_204), .B1(n_205), .B2(n_206), .Y(n_200) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g312 ( .A(n_207), .B(n_289), .Y(n_312) );
AND2x2_ASAP7_75t_L g380 ( .A(n_207), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g394 ( .A(n_207), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_207), .B(n_409), .Y(n_408) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_219), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2x1_ASAP7_75t_L g257 ( .A(n_209), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g350 ( .A(n_209), .B(n_343), .Y(n_350) );
AND2x2_ASAP7_75t_L g441 ( .A(n_209), .B(n_263), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_217), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_217), .A2(n_498), .B(n_500), .Y(n_497) );
OA21x2_ASAP7_75t_L g579 ( .A1(n_217), .A2(n_580), .B(n_584), .Y(n_579) );
OA21x2_ASAP7_75t_L g624 ( .A1(n_217), .A2(n_580), .B(n_584), .Y(n_624) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g252 ( .A(n_219), .Y(n_252) );
INVx2_ASAP7_75t_L g297 ( .A(n_219), .Y(n_297) );
AND2x2_ASAP7_75t_L g342 ( .A(n_219), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_221), .B(n_227), .Y(n_220) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_240), .Y(n_230) );
AND2x2_ASAP7_75t_L g384 ( .A(n_231), .B(n_385), .Y(n_384) );
OR2x6_ASAP7_75t_L g443 ( .A(n_231), .B(n_444), .Y(n_443) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx4_ASAP7_75t_L g273 ( .A(n_232), .Y(n_273) );
AND2x4_ASAP7_75t_L g281 ( .A(n_232), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g316 ( .A(n_232), .B(n_241), .Y(n_316) );
INVx2_ASAP7_75t_L g365 ( .A(n_232), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_232), .B(n_339), .Y(n_414) );
AND2x2_ASAP7_75t_L g451 ( .A(n_232), .B(n_269), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_232), .B(n_334), .Y(n_459) );
OR2x6_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
AND2x2_ASAP7_75t_L g292 ( .A(n_240), .B(n_281), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_240), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_SL g431 ( .A(n_240), .B(n_319), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_240), .B(n_332), .Y(n_453) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_241), .Y(n_271) );
AND2x2_ASAP7_75t_L g279 ( .A(n_241), .B(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_241), .Y(n_302) );
INVx2_ASAP7_75t_L g305 ( .A(n_241), .Y(n_305) );
INVx1_ASAP7_75t_L g338 ( .A(n_241), .Y(n_338) );
INVx1_ASAP7_75t_L g386 ( .A(n_241), .Y(n_386) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_249), .Y(n_241) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_242), .A2(n_519), .B(n_525), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
NAND2xp33_ASAP7_75t_L g250 ( .A(n_251), .B(n_254), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_252), .B(n_255), .Y(n_328) );
OR2x2_ASAP7_75t_L g400 ( .A(n_252), .B(n_401), .Y(n_400) );
AND4x1_ASAP7_75t_SL g446 ( .A(n_252), .B(n_428), .C(n_447), .D(n_448), .Y(n_446) );
OR2x2_ASAP7_75t_L g470 ( .A(n_253), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
AND2x2_ASAP7_75t_L g307 ( .A(n_256), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_256), .B(n_265), .Y(n_457) );
AND2x2_ASAP7_75t_L g482 ( .A(n_257), .B(n_342), .Y(n_482) );
OAI32xp33_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_267), .A3(n_272), .B1(n_274), .B2(n_277), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g355 ( .A(n_262), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g455 ( .A(n_262), .B(n_409), .Y(n_455) );
AND2x4_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
AND2x2_ASAP7_75t_L g351 ( .A(n_263), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g437 ( .A(n_263), .Y(n_437) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_264), .B(n_266), .Y(n_471) );
INVx3_ASAP7_75t_L g288 ( .A(n_265), .Y(n_288) );
NAND2x1p5_ASAP7_75t_L g466 ( .A(n_265), .B(n_393), .Y(n_466) );
INVx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_266), .Y(n_325) );
AND2x2_ASAP7_75t_L g344 ( .A(n_266), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g478 ( .A(n_268), .Y(n_478) );
NAND2x1_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_L g318 ( .A(n_269), .Y(n_318) );
NOR2x1_ASAP7_75t_L g419 ( .A(n_269), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_272), .B(n_378), .Y(n_377) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g310 ( .A(n_273), .B(n_278), .Y(n_310) );
AND2x4_ASAP7_75t_L g332 ( .A(n_273), .B(n_282), .Y(n_332) );
AND2x4_ASAP7_75t_SL g403 ( .A(n_273), .B(n_404), .Y(n_403) );
NOR2x1_ASAP7_75t_L g429 ( .A(n_273), .B(n_354), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_274), .A2(n_397), .B1(n_400), .B2(n_402), .Y(n_396) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx2_ASAP7_75t_SL g416 ( .A(n_275), .Y(n_416) );
INVx2_ASAP7_75t_L g308 ( .A(n_276), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_279), .B(n_285), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_279), .A2(n_415), .B1(n_418), .B2(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g339 ( .A(n_280), .Y(n_339) );
AND2x2_ASAP7_75t_L g362 ( .A(n_280), .B(n_321), .Y(n_362) );
INVx2_ASAP7_75t_L g285 ( .A(n_281), .Y(n_285) );
OAI21xp5_ASAP7_75t_SL g283 ( .A1(n_284), .A2(n_286), .B(n_290), .Y(n_283) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_287), .A2(n_359), .B1(n_363), .B2(n_364), .Y(n_358) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_288), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_288), .B(n_356), .Y(n_372) );
INVx1_ASAP7_75t_L g376 ( .A(n_288), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
NOR3xp33_ASAP7_75t_L g293 ( .A(n_294), .B(n_309), .C(n_313), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_298), .B1(n_303), .B2(n_306), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g323 ( .A(n_296), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g363 ( .A(n_296), .B(n_350), .Y(n_363) );
AND2x2_ASAP7_75t_L g415 ( .A(n_296), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g432 ( .A(n_296), .B(n_382), .Y(n_432) );
AND2x2_ASAP7_75t_L g487 ( .A(n_296), .B(n_381), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx4_ASAP7_75t_L g354 ( .A(n_299), .Y(n_354) );
AND2x2_ASAP7_75t_L g364 ( .A(n_299), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx2_ASAP7_75t_L g369 ( .A(n_302), .Y(n_369) );
AND2x2_ASAP7_75t_L g378 ( .A(n_302), .B(n_362), .Y(n_378) );
INVx1_ASAP7_75t_L g413 ( .A(n_304), .Y(n_413) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g334 ( .A(n_305), .Y(n_334) );
INVxp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_307), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_308), .B(n_376), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_317), .B(n_322), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_315), .B(n_354), .Y(n_463) );
INVx2_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AOI21xp33_ASAP7_75t_SL g326 ( .A1(n_318), .A2(n_327), .B(n_329), .Y(n_326) );
AND2x2_ASAP7_75t_L g473 ( .A(n_318), .B(n_332), .Y(n_473) );
AND2x4_ASAP7_75t_L g336 ( .A(n_319), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_SL g370 ( .A(n_319), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_319), .B(n_386), .Y(n_452) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI21xp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_335), .B(n_340), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_332), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_332), .B(n_337), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_333), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g395 ( .A(n_333), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_333), .Y(n_399) );
AND2x2_ASAP7_75t_L g483 ( .A(n_333), .B(n_451), .Y(n_483) );
AND2x2_ASAP7_75t_L g486 ( .A(n_333), .B(n_403), .Y(n_486) );
INVx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x4_ASAP7_75t_SL g337 ( .A(n_338), .B(n_339), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_338), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
INVx1_ASAP7_75t_L g465 ( .A(n_342), .Y(n_465) );
AND2x2_ASAP7_75t_L g356 ( .A(n_343), .B(n_357), .Y(n_356) );
NAND4xp75_ASAP7_75t_L g346 ( .A(n_347), .B(n_366), .C(n_387), .D(n_405), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_358), .Y(n_347) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_350), .B(n_437), .Y(n_436) );
NAND2x1p5_ASAP7_75t_L g422 ( .A(n_351), .B(n_416), .Y(n_422) );
NAND2xp5_ASAP7_75t_R g438 ( .A(n_354), .B(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g488 ( .A(n_354), .Y(n_488) );
INVx2_ASAP7_75t_L g401 ( .A(n_356), .Y(n_401) );
BUFx3_ASAP7_75t_L g393 ( .A(n_357), .Y(n_393) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g444 ( .A(n_362), .Y(n_444) );
AND2x2_ASAP7_75t_L g398 ( .A(n_364), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g420 ( .A(n_365), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_371), .B(n_373), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_369), .B(n_403), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_370), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_372), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_377), .B1(n_379), .B2(n_383), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
OA21x2_ASAP7_75t_L g388 ( .A1(n_381), .A2(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g409 ( .A(n_381), .Y(n_409) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g440 ( .A(n_382), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g448 ( .A(n_382), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_383), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g418 ( .A(n_386), .B(n_419), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_394), .B(n_396), .Y(n_387) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g435 ( .A(n_392), .B(n_436), .Y(n_435) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_399), .Y(n_447) );
INVx2_ASAP7_75t_SL g439 ( .A(n_403), .Y(n_439) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_417), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_410), .B1(n_412), .B2(n_415), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g468 ( .A(n_412), .Y(n_468) );
NOR2x1_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
INVx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_460), .Y(n_423) );
NAND3xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_433), .C(n_445), .Y(n_424) );
NOR2x1_ASAP7_75t_L g425 ( .A(n_426), .B(n_430), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
AOI22xp33_ASAP7_75t_SL g433 ( .A1(n_434), .A2(n_438), .B1(n_440), .B2(n_442), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NOR3xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_449), .C(n_456), .Y(n_445) );
AOI21xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_453), .B(n_454), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_479), .Y(n_460) );
NOR3xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_469), .C(n_476), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B1(n_467), .B2(n_468), .Y(n_462) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g476 ( .A(n_470), .B(n_475), .C(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVxp67_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AOI222xp33_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_483), .B1(n_484), .B2(n_486), .C1(n_487), .C2(n_488), .Y(n_479) );
INVx1_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
XNOR2x1_ASAP7_75t_L g821 ( .A(n_489), .B(n_822), .Y(n_821) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_673), .Y(n_489) );
NOR3xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_628), .C(n_657), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_492), .B(n_601), .Y(n_491) );
AOI221xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_526), .B1(n_547), .B2(n_558), .C(n_562), .Y(n_492) );
INVx3_ASAP7_75t_SL g718 ( .A(n_493), .Y(n_718) );
AND2x2_ASAP7_75t_SL g493 ( .A(n_494), .B(n_505), .Y(n_493) );
NAND2x1p5_ASAP7_75t_L g564 ( .A(n_494), .B(n_517), .Y(n_564) );
INVx4_ASAP7_75t_L g599 ( .A(n_494), .Y(n_599) );
AND2x2_ASAP7_75t_L g621 ( .A(n_494), .B(n_518), .Y(n_621) );
AND2x2_ASAP7_75t_L g627 ( .A(n_494), .B(n_566), .Y(n_627) );
INVx5_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g596 ( .A(n_495), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_495), .B(n_517), .Y(n_672) );
AND2x2_ASAP7_75t_L g677 ( .A(n_495), .B(n_518), .Y(n_677) );
AND2x2_ASAP7_75t_L g689 ( .A(n_495), .B(n_550), .Y(n_689) );
NOR2x1_ASAP7_75t_SL g728 ( .A(n_495), .B(n_566), .Y(n_728) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g557 ( .A(n_505), .Y(n_557) );
AND2x2_ASAP7_75t_L g661 ( .A(n_505), .B(n_610), .Y(n_661) );
AND2x2_ASAP7_75t_L g758 ( .A(n_505), .B(n_689), .Y(n_758) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_517), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g590 ( .A(n_507), .Y(n_590) );
INVx2_ASAP7_75t_L g612 ( .A(n_507), .Y(n_612) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B(n_515), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_508), .B(n_516), .Y(n_515) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_508), .A2(n_509), .B(n_515), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_514), .Y(n_509) );
AND2x2_ASAP7_75t_L g587 ( .A(n_517), .B(n_549), .Y(n_587) );
INVx2_ASAP7_75t_L g591 ( .A(n_517), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_517), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g690 ( .A(n_517), .B(n_655), .Y(n_690) );
OR2x2_ASAP7_75t_L g737 ( .A(n_517), .B(n_550), .Y(n_737) );
INVx4_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_518), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_524), .Y(n_519) );
AND2x2_ASAP7_75t_L g734 ( .A(n_526), .B(n_615), .Y(n_734) );
AND2x2_ASAP7_75t_L g784 ( .A(n_526), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g660 ( .A(n_527), .B(n_604), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_538), .Y(n_527) );
AND2x2_ASAP7_75t_L g593 ( .A(n_528), .B(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g623 ( .A(n_528), .B(n_624), .Y(n_623) );
AND2x4_ASAP7_75t_L g644 ( .A(n_528), .B(n_624), .Y(n_644) );
AND2x4_ASAP7_75t_L g679 ( .A(n_528), .B(n_667), .Y(n_679) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g560 ( .A(n_529), .Y(n_560) );
OAI21x1_ASAP7_75t_SL g529 ( .A1(n_530), .A2(n_532), .B(n_536), .Y(n_529) );
INVx1_ASAP7_75t_L g537 ( .A(n_531), .Y(n_537) );
AND2x2_ASAP7_75t_L g606 ( .A(n_538), .B(n_559), .Y(n_606) );
AND2x2_ASAP7_75t_L g692 ( .A(n_538), .B(n_624), .Y(n_692) );
AND2x2_ASAP7_75t_L g703 ( .A(n_538), .B(n_568), .Y(n_703) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g567 ( .A(n_539), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g634 ( .A(n_539), .B(n_569), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_541), .B(n_545), .Y(n_540) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_557), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_549), .B(n_599), .Y(n_656) );
AND2x2_ASAP7_75t_L g700 ( .A(n_549), .B(n_566), .Y(n_700) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_550), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g610 ( .A(n_550), .Y(n_610) );
BUFx3_ASAP7_75t_L g619 ( .A(n_550), .Y(n_619) );
AND2x2_ASAP7_75t_L g642 ( .A(n_550), .B(n_612), .Y(n_642) );
OAI322xp33_ASAP7_75t_L g562 ( .A1(n_557), .A2(n_563), .A3(n_567), .B1(n_577), .B2(n_585), .C1(n_592), .C2(n_597), .Y(n_562) );
INVx1_ASAP7_75t_L g723 ( .A(n_557), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_558), .B(n_598), .Y(n_597) );
AND2x4_ASAP7_75t_L g636 ( .A(n_558), .B(n_578), .Y(n_636) );
INVx2_ASAP7_75t_L g681 ( .A(n_558), .Y(n_681) );
AND2x2_ASAP7_75t_L g697 ( .A(n_558), .B(n_639), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_558), .B(n_715), .Y(n_745) );
AND2x4_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
AND2x2_ASAP7_75t_SL g648 ( .A(n_559), .B(n_624), .Y(n_648) );
OR2x2_ASAP7_75t_L g669 ( .A(n_559), .B(n_586), .Y(n_669) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx2_ASAP7_75t_L g641 ( .A(n_560), .Y(n_641) );
INVx2_ASAP7_75t_L g586 ( .A(n_561), .Y(n_586) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_561), .Y(n_588) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g631 ( .A(n_564), .Y(n_631) );
INVxp67_ASAP7_75t_SL g651 ( .A(n_565), .Y(n_651) );
INVx1_ASAP7_75t_L g749 ( .A(n_565), .Y(n_749) );
INVxp67_ASAP7_75t_SL g764 ( .A(n_565), .Y(n_764) );
NAND2x1_ASAP7_75t_L g774 ( .A(n_567), .B(n_578), .Y(n_774) );
INVx1_ASAP7_75t_L g781 ( .A(n_567), .Y(n_781) );
BUFx2_ASAP7_75t_L g615 ( .A(n_568), .Y(n_615) );
AND2x2_ASAP7_75t_L g691 ( .A(n_568), .B(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx3_ASAP7_75t_L g600 ( .A(n_569), .Y(n_600) );
INVxp67_ASAP7_75t_L g604 ( .A(n_569), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_575), .Y(n_570) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_577), .B(n_593), .C(n_595), .Y(n_592) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_SL g613 ( .A(n_578), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_578), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g765 ( .A(n_578), .B(n_714), .Y(n_765) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g667 ( .A(n_579), .Y(n_667) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_579), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B1(n_588), .B2(n_589), .Y(n_585) );
AND2x4_ASAP7_75t_SL g714 ( .A(n_586), .B(n_594), .Y(n_714) );
AND2x2_ASAP7_75t_L g727 ( .A(n_587), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_588), .Y(n_729) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx2_ASAP7_75t_L g686 ( .A(n_590), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_590), .B(n_599), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_591), .B(n_609), .Y(n_608) );
AND3x2_ASAP7_75t_L g626 ( .A(n_591), .B(n_619), .C(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g650 ( .A(n_591), .Y(n_650) );
AND2x2_ASAP7_75t_L g763 ( .A(n_591), .B(n_764), .Y(n_763) );
BUFx2_ASAP7_75t_L g639 ( .A(n_594), .Y(n_639) );
INVx1_ASAP7_75t_L g717 ( .A(n_594), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_595), .B(n_618), .Y(n_756) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_596), .B(n_700), .Y(n_705) );
AND2x4_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AND2x2_ASAP7_75t_L g696 ( .A(n_599), .B(n_642), .Y(n_696) );
INVx1_ASAP7_75t_SL g647 ( .A(n_600), .Y(n_647) );
AND2x2_ASAP7_75t_L g755 ( .A(n_600), .B(n_667), .Y(n_755) );
AND2x2_ASAP7_75t_L g776 ( .A(n_600), .B(n_648), .Y(n_776) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_607), .B1(n_613), .B2(n_616), .C(n_622), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g768 ( .A(n_604), .Y(n_768) );
AOI21xp33_ASAP7_75t_SL g622 ( .A1(n_605), .A2(n_623), .B(n_625), .Y(n_622) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g614 ( .A(n_606), .B(n_615), .Y(n_614) );
AOI222xp33_ASAP7_75t_L g637 ( .A1(n_606), .A2(n_638), .B1(n_640), .B2(n_645), .C1(n_649), .C2(n_652), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_606), .B(n_755), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_607), .A2(n_636), .B1(n_659), .B2(n_661), .Y(n_658) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g643 ( .A(n_610), .Y(n_643) );
AND2x2_ASAP7_75t_L g762 ( .A(n_610), .B(n_728), .Y(n_762) );
OAI32xp33_ASAP7_75t_L g766 ( .A1(n_610), .A2(n_635), .A3(n_687), .B1(n_695), .B2(n_767), .Y(n_766) );
AND2x2_ASAP7_75t_L g771 ( .A(n_610), .B(n_621), .Y(n_771) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g655 ( .A(n_612), .Y(n_655) );
OAI21xp5_ASAP7_75t_SL g662 ( .A1(n_613), .A2(n_663), .B(n_670), .Y(n_662) );
INVx1_ASAP7_75t_L g726 ( .A(n_615), .Y(n_726) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
AND2x2_ASAP7_75t_L g630 ( .A(n_618), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g638 ( .A(n_621), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g711 ( .A(n_621), .B(n_642), .Y(n_711) );
INVx1_ASAP7_75t_SL g782 ( .A(n_623), .Y(n_782) );
AND2x2_ASAP7_75t_L g716 ( .A(n_624), .B(n_717), .Y(n_716) );
OAI222xp33_ASAP7_75t_L g769 ( .A1(n_625), .A2(n_678), .B1(n_757), .B2(n_770), .C1(n_772), .C2(n_774), .Y(n_769) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x4_ASAP7_75t_L g742 ( .A(n_627), .B(n_743), .Y(n_742) );
OAI21xp33_ASAP7_75t_SL g628 ( .A1(n_629), .A2(n_632), .B(n_637), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_631), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g710 ( .A(n_633), .Y(n_710) );
INVx1_ASAP7_75t_L g678 ( .A(n_634), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_634), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g732 ( .A(n_639), .Y(n_732) );
AO22x1_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_643), .B2(n_644), .Y(n_640) );
OAI322xp33_ASAP7_75t_L g752 ( .A1(n_641), .A2(n_702), .A3(n_705), .B1(n_753), .B2(n_754), .C1(n_756), .C2(n_757), .Y(n_752) );
AND2x2_ASAP7_75t_SL g676 ( .A(n_642), .B(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g671 ( .A(n_643), .B(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g731 ( .A(n_644), .B(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g773 ( .A(n_644), .B(n_703), .Y(n_773) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g753 ( .A(n_647), .Y(n_753) );
INVx1_ASAP7_75t_SL g682 ( .A(n_648), .Y(n_682) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .Y(n_653) );
OR2x2_ASAP7_75t_L g684 ( .A(n_656), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g722 ( .A(n_656), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_662), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_668), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g695 ( .A(n_666), .B(n_681), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_666), .B(n_703), .Y(n_702) );
BUFx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g725 ( .A(n_669), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NOR2x1_ASAP7_75t_L g673 ( .A(n_674), .B(n_738), .Y(n_673) );
NAND4xp25_ASAP7_75t_L g674 ( .A(n_675), .B(n_693), .C(n_706), .D(n_719), .Y(n_674) );
AOI322xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_678), .A3(n_679), .B1(n_680), .B2(n_683), .C1(n_688), .C2(n_691), .Y(n_675) );
AOI211xp5_ASAP7_75t_L g775 ( .A1(n_676), .A2(n_776), .B(n_777), .C(n_780), .Y(n_775) );
AND2x2_ASAP7_75t_L g787 ( .A(n_677), .B(n_764), .Y(n_787) );
INVx1_ASAP7_75t_L g709 ( .A(n_679), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_679), .B(n_714), .Y(n_751) );
NAND2xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_687), .B(n_700), .Y(n_767) );
AND2x4_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
AOI222xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B1(n_697), .B2(n_698), .C1(n_701), .C2(n_704), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_696), .A2(n_707), .B1(n_710), .B2(n_711), .C(n_712), .Y(n_706) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AOI21xp33_ASAP7_75t_SL g712 ( .A1(n_713), .A2(n_715), .B(n_718), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_724), .B1(n_727), .B2(n_729), .C(n_730), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g779 ( .A(n_728), .Y(n_779) );
AOI21xp33_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_733), .B(n_735), .Y(n_730) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx2_ASAP7_75t_L g743 ( .A(n_737), .Y(n_743) );
OR2x2_ASAP7_75t_L g778 ( .A(n_737), .B(n_779), .Y(n_778) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_759), .C(n_775), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_752), .Y(n_739) );
OAI21xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_744), .B(n_746), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_750), .Y(n_746) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AOI221xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_765), .B1(n_766), .B2(n_768), .C(n_769), .Y(n_759) );
INVxp67_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NOR2x1_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_774), .B(n_778), .Y(n_777) );
O2A1O1Ixp33_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_782), .B(n_783), .C(n_786), .Y(n_780) );
INVxp67_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
CKINVDCx11_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_789), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_790), .Y(n_798) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx3_ASAP7_75t_SL g796 ( .A(n_797), .Y(n_796) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx3_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
OAI21x1_ASAP7_75t_SL g817 ( .A1(n_804), .A2(n_818), .B(n_820), .Y(n_817) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
BUFx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
BUFx2_ASAP7_75t_R g819 ( .A(n_807), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
BUFx3_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
CKINVDCx11_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
CKINVDCx8_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx2_ASAP7_75t_L g825 ( .A(n_821), .Y(n_825) );
INVx2_ASAP7_75t_SL g827 ( .A(n_828), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_829), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_829), .B(n_837), .Y(n_836) );
INVx3_ASAP7_75t_R g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
AND2x2_ASAP7_75t_SL g831 ( .A(n_832), .B(n_833), .Y(n_831) );
endmodule