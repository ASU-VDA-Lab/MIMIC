module fake_jpeg_16163_n_239 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_239);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_239;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_2),
.B(n_4),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx5_ASAP7_75t_SL g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g91 ( 
.A(n_41),
.Y(n_91)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_62),
.B1(n_37),
.B2(n_34),
.Y(n_76)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_54),
.Y(n_67)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx5_ASAP7_75t_SL g54 ( 
.A(n_29),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_58),
.Y(n_79)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_61),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_7),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_33),
.B1(n_32),
.B2(n_17),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_71),
.A2(n_77),
.B1(n_11),
.B2(n_12),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_35),
.B(n_26),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_88),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_35),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_74),
.A2(n_18),
.B1(n_9),
.B2(n_10),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_76),
.B(n_95),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_51),
.A2(n_17),
.B1(n_32),
.B2(n_33),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_37),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_80),
.B(n_82),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_34),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_15),
.C(n_25),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_23),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_89),
.B(n_90),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_60),
.A2(n_25),
.B(n_23),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_26),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_96),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_19),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_46),
.B(n_28),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_39),
.B(n_7),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_97),
.B(n_12),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_40),
.B(n_14),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_28),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_103),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_28),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_38),
.Y(n_104)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_8),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_131),
.Y(n_136)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_81),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_112),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_66),
.Y(n_112)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_115),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_77),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_114),
.A2(n_123),
.B1(n_128),
.B2(n_109),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_14),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_66),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_121),
.Y(n_143)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_11),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_125),
.B(n_72),
.Y(n_149)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_71),
.A2(n_69),
.B1(n_78),
.B2(n_84),
.Y(n_128)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_133),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_74),
.B(n_79),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_65),
.B(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_65),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_72),
.B(n_86),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_78),
.A2(n_92),
.B1(n_87),
.B2(n_86),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_134),
.A2(n_102),
.B1(n_87),
.B2(n_99),
.Y(n_139)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_150),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_152),
.B1(n_161),
.B2(n_114),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_99),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_142),
.B(n_154),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_65),
.B(n_104),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_145),
.B(n_149),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_126),
.B(n_85),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_160),
.C(n_154),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_116),
.A2(n_102),
.B1(n_75),
.B2(n_85),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_75),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_158),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_81),
.B(n_70),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_111),
.B(n_125),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_124),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_110),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_70),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_70),
.C(n_116),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_165),
.C(n_166),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_139),
.B1(n_148),
.B2(n_129),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_106),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_123),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_105),
.C(n_107),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_141),
.C(n_143),
.Y(n_184)
);

AOI221xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_136),
.B1(n_155),
.B2(n_140),
.C(n_143),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_136),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_171),
.B(n_175),
.Y(n_185)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_173),
.B(n_178),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_118),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_110),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_176),
.B(n_177),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_149),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_120),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_180),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_112),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_119),
.B1(n_117),
.B2(n_129),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_181),
.A2(n_159),
.B1(n_138),
.B2(n_157),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_171),
.B(n_194),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_193),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_142),
.C(n_152),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_191),
.C(n_164),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_175),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_187),
.B(n_194),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_189),
.A2(n_197),
.B1(n_173),
.B2(n_172),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_146),
.C(n_159),
.Y(n_191)
);

NOR3xp33_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_177),
.C(n_141),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_164),
.A2(n_146),
.B(n_157),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_195),
.A2(n_169),
.B(n_170),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_200),
.C(n_181),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_199),
.A2(n_188),
.B(n_190),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_203),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_170),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_202),
.A2(n_185),
.B(n_187),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_165),
.C(n_167),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_208),
.C(n_195),
.Y(n_210)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_207),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_191),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_189),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_215),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_163),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_216),
.B(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_204),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_223),
.B(n_202),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_211),
.A2(n_203),
.B1(n_200),
.B2(n_205),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_225),
.A2(n_214),
.B1(n_202),
.B2(n_210),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_227),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_222),
.A2(n_215),
.B1(n_206),
.B2(n_212),
.Y(n_228)
);

AOI322xp5_ASAP7_75t_L g232 ( 
.A1(n_228),
.A2(n_230),
.A3(n_219),
.B1(n_224),
.B2(n_225),
.C1(n_108),
.C2(n_130),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_201),
.C(n_144),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_219),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_147),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_229),
.A2(n_221),
.B(n_224),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_231),
.A2(n_232),
.B(n_234),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_135),
.B1(n_147),
.B2(n_113),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_135),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_238),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);


endmodule