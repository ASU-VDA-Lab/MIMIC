module fake_jpeg_4929_n_129 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_24),
.Y(n_40)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_28),
.Y(n_33)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx6p67_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_23),
.A2(n_19),
.B1(n_22),
.B2(n_18),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_14),
.B1(n_18),
.B2(n_13),
.Y(n_53)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_11),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_50),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_48),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_44),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_26),
.B(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_53),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_20),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_52),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_39),
.B1(n_38),
.B2(n_35),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_63),
.B1(n_46),
.B2(n_36),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_39),
.B1(n_33),
.B2(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_53),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_39),
.B1(n_25),
.B2(n_45),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_56),
.B1(n_61),
.B2(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_50),
.C(n_43),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_69),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_64),
.C(n_65),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_30),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_36),
.B(n_55),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_60),
.B(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_77),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_19),
.B1(n_55),
.B2(n_11),
.Y(n_84)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_16),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_86),
.B(n_87),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_90),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_88),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_79),
.B1(n_71),
.B2(n_68),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_76),
.B(n_21),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_76),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_12),
.B(n_22),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_16),
.B(n_13),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_95),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_85),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_98),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_52),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_75),
.B(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_100),
.B(n_105),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_31),
.C(n_32),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_104),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_99),
.C(n_92),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_92),
.B(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_108),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_29),
.B1(n_30),
.B2(n_21),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_1),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_104),
.A2(n_30),
.B1(n_29),
.B2(n_32),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_113),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_102),
.A2(n_32),
.B1(n_52),
.B2(n_3),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_103),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_115),
.B(n_4),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_112),
.A2(n_106),
.B(n_7),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_120),
.C(n_115),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_106),
.C(n_7),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_113),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_122),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_R g125 ( 
.A1(n_123),
.A2(n_111),
.B1(n_114),
.B2(n_110),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_8),
.B(n_9),
.C(n_113),
.Y(n_126)
);

NAND2x1p5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_126),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_127),
.Y(n_129)
);


endmodule