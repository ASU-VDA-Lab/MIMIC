module fake_netlist_1_5318_n_526 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_526);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_526;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_420;
wire n_165;
wire n_195;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_SL g77 ( .A(n_46), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_47), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_2), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_60), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_24), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_41), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_2), .Y(n_83) );
NAND2xp5_ASAP7_75t_L g84 ( .A(n_29), .B(n_57), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_13), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_52), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_11), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_34), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_10), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_22), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_21), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_7), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_8), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_42), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_72), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_23), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_62), .Y(n_97) );
OR2x2_ASAP7_75t_L g98 ( .A(n_9), .B(n_48), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_18), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_54), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_45), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_27), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_40), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_70), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_43), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_4), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_56), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_30), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_4), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_68), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_17), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_82), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_82), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_86), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_89), .B(n_0), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_86), .Y(n_116) );
AND2x6_ASAP7_75t_L g117 ( .A(n_88), .B(n_36), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_89), .B(n_0), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_88), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_90), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_90), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_107), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_109), .B(n_1), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_107), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_109), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_98), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_100), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_78), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_94), .B(n_1), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_79), .B(n_3), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_83), .B(n_3), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_95), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_96), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_97), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_114), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_126), .B(n_83), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_114), .Y(n_137) );
INVx1_ASAP7_75t_SL g138 ( .A(n_126), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_117), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_126), .B(n_79), .Y(n_140) );
AND2x6_ASAP7_75t_L g141 ( .A(n_126), .B(n_101), .Y(n_141) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_131), .A2(n_87), .B1(n_85), .B2(n_106), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_112), .B(n_102), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_114), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_112), .B(n_80), .Y(n_145) );
INVxp67_ASAP7_75t_SL g146 ( .A(n_130), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_113), .B(n_103), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_113), .B(n_104), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_116), .B(n_80), .Y(n_149) );
INVx1_ASAP7_75t_SL g150 ( .A(n_127), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_114), .Y(n_151) );
AND2x6_ASAP7_75t_L g152 ( .A(n_131), .B(n_85), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_114), .Y(n_153) );
INVx5_ASAP7_75t_L g154 ( .A(n_117), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_117), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_114), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_122), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_122), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_116), .B(n_87), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_122), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_146), .B(n_115), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_150), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_139), .Y(n_163) );
AOI22xp33_ASAP7_75t_L g164 ( .A1(n_152), .A2(n_117), .B1(n_115), .B2(n_118), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_138), .Y(n_165) );
AOI22xp5_ASAP7_75t_L g166 ( .A1(n_152), .A2(n_123), .B1(n_118), .B2(n_132), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_144), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_138), .B(n_120), .Y(n_169) );
INVx1_ASAP7_75t_SL g170 ( .A(n_140), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_159), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_150), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_141), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_159), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_140), .B(n_123), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_159), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_144), .Y(n_178) );
BUFx12f_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_136), .B(n_120), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_159), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_136), .B(n_128), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g183 ( .A1(n_142), .A2(n_105), .B1(n_111), .B2(n_132), .Y(n_183) );
INVx5_ASAP7_75t_L g184 ( .A(n_141), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_136), .B(n_128), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_136), .B(n_124), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_145), .B(n_133), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_152), .A2(n_134), .B1(n_133), .B2(n_124), .Y(n_188) );
NAND2xp33_ASAP7_75t_L g189 ( .A(n_139), .B(n_117), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_152), .B(n_134), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_139), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_141), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_152), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_163), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_167), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_189), .A2(n_154), .B(n_139), .Y(n_197) );
BUFx2_ASAP7_75t_SL g198 ( .A(n_184), .Y(n_198) );
INVx1_ASAP7_75t_SL g199 ( .A(n_162), .Y(n_199) );
BUFx2_ASAP7_75t_L g200 ( .A(n_179), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_179), .Y(n_201) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_173), .Y(n_202) );
OR2x2_ASAP7_75t_L g203 ( .A(n_183), .B(n_143), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_163), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_167), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_191), .B(n_152), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_184), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_171), .Y(n_208) );
OR2x6_ASAP7_75t_SL g209 ( .A(n_180), .B(n_106), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_170), .A2(n_152), .B1(n_141), .B2(n_149), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_163), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_168), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_165), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_171), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_167), .Y(n_215) );
OR2x6_ASAP7_75t_L g216 ( .A(n_182), .B(n_139), .Y(n_216) );
BUFx12f_ASAP7_75t_L g217 ( .A(n_161), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_175), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_175), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_177), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_163), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_166), .A2(n_139), .B1(n_155), .B2(n_147), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_177), .A2(n_148), .B(n_147), .C(n_143), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_163), .Y(n_224) );
BUFx8_ASAP7_75t_L g225 ( .A(n_191), .Y(n_225) );
NAND2x1_ASAP7_75t_SL g226 ( .A(n_188), .B(n_119), .Y(n_226) );
INVx3_ASAP7_75t_L g227 ( .A(n_168), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_217), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_196), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_196), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_203), .B(n_161), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_205), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_208), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_203), .B(n_161), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_208), .Y(n_235) );
OAI22xp33_ASAP7_75t_L g236 ( .A1(n_199), .A2(n_166), .B1(n_188), .B2(n_165), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_205), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_223), .A2(n_169), .B(n_186), .C(n_176), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_213), .A2(n_164), .B(n_181), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_213), .A2(n_181), .B1(n_182), .B2(n_185), .Y(n_240) );
OR2x2_ASAP7_75t_L g241 ( .A(n_202), .B(n_161), .Y(n_241) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_217), .Y(n_242) );
CKINVDCx6p67_ASAP7_75t_R g243 ( .A(n_209), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_209), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_222), .A2(n_182), .B1(n_185), .B2(n_148), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_206), .B(n_176), .Y(n_246) );
AND2x4_ASAP7_75t_L g247 ( .A(n_206), .B(n_194), .Y(n_247) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_225), .Y(n_248) );
BUFx2_ASAP7_75t_SL g249 ( .A(n_201), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_225), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_214), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_206), .A2(n_141), .B1(n_182), .B2(n_185), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_206), .A2(n_141), .B1(n_185), .B2(n_194), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_225), .A2(n_141), .B1(n_187), .B2(n_193), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_234), .A2(n_210), .B1(n_216), .B2(n_220), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_241), .B(n_92), .Y(n_256) );
AOI222xp33_ASAP7_75t_L g257 ( .A1(n_231), .A2(n_93), .B1(n_218), .B2(n_220), .C1(n_219), .C2(n_214), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_231), .B(n_225), .Y(n_258) );
OAI221xp5_ASAP7_75t_L g259 ( .A1(n_241), .A2(n_226), .B1(n_129), .B2(n_219), .C(n_218), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_243), .A2(n_200), .B1(n_201), .B2(n_216), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_243), .A2(n_201), .B1(n_200), .B2(n_117), .Y(n_261) );
AOI211xp5_ASAP7_75t_L g262 ( .A1(n_244), .A2(n_98), .B(n_121), .C(n_119), .Y(n_262) );
NOR3xp33_ASAP7_75t_L g263 ( .A(n_236), .B(n_125), .C(n_99), .Y(n_263) );
OR2x6_ASAP7_75t_L g264 ( .A(n_250), .B(n_216), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_228), .B(n_226), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_248), .Y(n_266) );
AOI22xp33_ASAP7_75t_SL g267 ( .A1(n_250), .A2(n_125), .B1(n_198), .B2(n_119), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_234), .A2(n_216), .B1(n_215), .B2(n_184), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_240), .A2(n_216), .B1(n_215), .B2(n_184), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_240), .A2(n_184), .B1(n_193), .B2(n_168), .Y(n_270) );
AOI22xp33_ASAP7_75t_SL g271 ( .A1(n_245), .A2(n_125), .B1(n_198), .B2(n_121), .Y(n_271) );
INVxp67_ASAP7_75t_L g272 ( .A(n_242), .Y(n_272) );
AOI321xp33_ASAP7_75t_L g273 ( .A1(n_246), .A2(n_125), .A3(n_121), .B1(n_108), .B2(n_84), .C(n_9), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_243), .B(n_212), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_245), .A2(n_117), .B1(n_227), .B2(n_212), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_229), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_276), .Y(n_277) );
AOI21xp33_ASAP7_75t_L g278 ( .A1(n_259), .A2(n_238), .B(n_235), .Y(n_278) );
INVx2_ASAP7_75t_SL g279 ( .A(n_264), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_255), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_271), .A2(n_247), .B1(n_249), .B2(n_251), .Y(n_281) );
OAI21xp33_ASAP7_75t_SL g282 ( .A1(n_275), .A2(n_233), .B(n_235), .Y(n_282) );
AOI211xp5_ASAP7_75t_SL g283 ( .A1(n_262), .A2(n_91), .B(n_239), .C(n_233), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_271), .A2(n_247), .B1(n_249), .B2(n_251), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_265), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_266), .B(n_229), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_256), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_257), .A2(n_252), .B1(n_247), .B2(n_254), .Y(n_288) );
OAI21xp5_ASAP7_75t_L g289 ( .A1(n_263), .A2(n_238), .B(n_239), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_258), .A2(n_247), .B1(n_117), .B2(n_253), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_264), .Y(n_291) );
NOR2xp33_ASAP7_75t_R g292 ( .A(n_274), .B(n_81), .Y(n_292) );
OAI322xp33_ASAP7_75t_L g293 ( .A1(n_272), .A2(n_122), .A3(n_77), .B1(n_81), .B2(n_110), .C1(n_160), .C2(n_158), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_264), .Y(n_294) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_273), .A2(n_122), .B1(n_232), .B2(n_230), .C(n_229), .Y(n_295) );
OR2x6_ASAP7_75t_L g296 ( .A(n_269), .B(n_230), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_260), .Y(n_297) );
NAND4xp25_ASAP7_75t_L g298 ( .A(n_261), .B(n_160), .C(n_137), .D(n_151), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_291), .B(n_230), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_277), .Y(n_300) );
AOI22xp33_ASAP7_75t_SL g301 ( .A1(n_297), .A2(n_268), .B1(n_237), .B2(n_232), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_285), .B(n_232), .Y(n_302) );
INVxp67_ASAP7_75t_SL g303 ( .A(n_286), .Y(n_303) );
AND4x1_ASAP7_75t_L g304 ( .A(n_283), .B(n_267), .C(n_6), .D(n_7), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_277), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_280), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_285), .B(n_237), .Y(n_307) );
AOI211x1_ASAP7_75t_SL g308 ( .A1(n_278), .A2(n_122), .B(n_237), .C(n_270), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_291), .B(n_19), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_280), .B(n_267), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_295), .A2(n_110), .B1(n_227), .B2(n_212), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_286), .B(n_5), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_296), .Y(n_313) );
NOR2x1_ASAP7_75t_L g314 ( .A(n_296), .B(n_207), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_296), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_294), .Y(n_316) );
AOI322xp5_ASAP7_75t_L g317 ( .A1(n_287), .A2(n_5), .A3(n_6), .B1(n_8), .B2(n_10), .C1(n_11), .C2(n_12), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_296), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_297), .B(n_12), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_279), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_279), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_282), .Y(n_322) );
NOR3xp33_ASAP7_75t_L g323 ( .A(n_289), .B(n_137), .C(n_151), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_292), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_288), .B(n_13), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_284), .B(n_14), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_290), .B(n_71), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_303), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_306), .Y(n_330) );
OAI21x1_ASAP7_75t_L g331 ( .A1(n_314), .A2(n_298), .B(n_221), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_306), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_325), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_314), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_300), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_306), .B(n_14), .Y(n_336) );
AOI211xp5_ASAP7_75t_L g337 ( .A1(n_326), .A2(n_293), .B(n_158), .C(n_157), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_302), .B(n_15), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_302), .B(n_15), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_316), .B(n_300), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_307), .B(n_16), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_305), .Y(n_342) );
OAI221xp5_ASAP7_75t_L g343 ( .A1(n_304), .A2(n_317), .B1(n_319), .B2(n_327), .C(n_301), .Y(n_343) );
AND4x1_ASAP7_75t_L g344 ( .A(n_319), .B(n_16), .C(n_20), .D(n_25), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_307), .B(n_312), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_304), .B(n_26), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_305), .B(n_157), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_312), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_299), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_320), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_322), .B(n_157), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_322), .B(n_156), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_310), .B(n_156), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_315), .B(n_28), .Y(n_354) );
AOI211xp5_ASAP7_75t_SL g355 ( .A1(n_328), .A2(n_193), .B(n_168), .C(n_174), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_310), .B(n_31), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_321), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_299), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_320), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_315), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_313), .B(n_32), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_313), .B(n_33), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_299), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_327), .B(n_35), .Y(n_364) );
AOI32xp33_ASAP7_75t_L g365 ( .A1(n_328), .A2(n_174), .A3(n_193), .B1(n_135), .B2(n_153), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_318), .B(n_37), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_317), .B(n_38), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_299), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_324), .B(n_39), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_318), .B(n_135), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_324), .B(n_44), .Y(n_371) );
NOR2x1_ASAP7_75t_L g372 ( .A(n_328), .B(n_207), .Y(n_372) );
OAI311xp33_ASAP7_75t_L g373 ( .A1(n_311), .A2(n_153), .A3(n_135), .B1(n_51), .C1(n_53), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_348), .B(n_324), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_329), .Y(n_375) );
OR2x2_ASAP7_75t_SL g376 ( .A(n_340), .B(n_324), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_360), .B(n_324), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_350), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_350), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_357), .B(n_324), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_359), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_334), .B(n_309), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_359), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_345), .B(n_309), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_333), .B(n_328), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_340), .B(n_309), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_357), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_360), .B(n_309), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_336), .Y(n_389) );
NOR3xp33_ASAP7_75t_L g390 ( .A(n_343), .B(n_323), .C(n_311), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_344), .B(n_49), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_342), .B(n_50), .Y(n_392) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_372), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_349), .B(n_55), .Y(n_394) );
OAI221xp5_ASAP7_75t_L g395 ( .A1(n_346), .A2(n_308), .B1(n_135), .B2(n_153), .C(n_174), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_330), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_342), .B(n_58), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_330), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_335), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_332), .B(n_308), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_349), .B(n_59), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_367), .A2(n_221), .B1(n_204), .B2(n_227), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_334), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_335), .B(n_153), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_338), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_363), .B(n_61), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_363), .B(n_368), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_368), .B(n_63), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_351), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_351), .B(n_64), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_358), .B(n_65), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_352), .Y(n_412) );
AND2x2_ASAP7_75t_SL g413 ( .A(n_354), .B(n_155), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_352), .B(n_66), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_354), .B(n_67), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_353), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_370), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_339), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_361), .B(n_69), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_341), .B(n_73), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_390), .A2(n_356), .B1(n_364), .B2(n_373), .C(n_371), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_375), .Y(n_422) );
OAI32xp33_ASAP7_75t_L g423 ( .A1(n_385), .A2(n_369), .A3(n_366), .B1(n_362), .B2(n_361), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_378), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_379), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_381), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_387), .B(n_366), .Y(n_427) );
OAI21xp5_ASAP7_75t_L g428 ( .A1(n_391), .A2(n_355), .B(n_331), .Y(n_428) );
NOR2x1_ASAP7_75t_L g429 ( .A(n_403), .B(n_362), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_383), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_405), .A2(n_337), .B1(n_331), .B2(n_347), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_418), .B(n_347), .Y(n_432) );
XOR2xp5_ASAP7_75t_L g433 ( .A(n_384), .B(n_74), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_396), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_380), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_417), .B(n_365), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_398), .Y(n_437) );
INVxp67_ASAP7_75t_L g438 ( .A(n_374), .Y(n_438) );
OAI321xp33_ASAP7_75t_L g439 ( .A1(n_393), .A2(n_75), .A3(n_76), .B1(n_204), .B2(n_221), .C(n_211), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_407), .Y(n_440) );
INVx2_ASAP7_75t_SL g441 ( .A(n_386), .Y(n_441) );
NOR2x1_ASAP7_75t_SL g442 ( .A(n_388), .B(n_207), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_377), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_416), .A2(n_227), .B1(n_212), .B2(n_174), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_399), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_409), .Y(n_446) );
XNOR2x1_ASAP7_75t_L g447 ( .A(n_415), .B(n_155), .Y(n_447) );
NAND2x1_ASAP7_75t_SL g448 ( .A(n_403), .B(n_190), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_412), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_420), .B(n_224), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_389), .B(n_190), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g452 ( .A1(n_376), .A2(n_184), .B1(n_155), .B2(n_211), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_400), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_400), .Y(n_454) );
XNOR2xp5_ASAP7_75t_L g455 ( .A(n_413), .B(n_197), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_382), .Y(n_456) );
XNOR2xp5_ASAP7_75t_L g457 ( .A(n_402), .B(n_178), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_419), .Y(n_458) );
CKINVDCx14_ASAP7_75t_R g459 ( .A(n_408), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_406), .B(n_178), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_404), .Y(n_461) );
XNOR2x1_ASAP7_75t_L g462 ( .A(n_406), .B(n_155), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_404), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_392), .Y(n_464) );
NAND2xp33_ASAP7_75t_L g465 ( .A(n_397), .B(n_224), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_394), .B(n_401), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_420), .A2(n_195), .B1(n_211), .B2(n_172), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_411), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_414), .Y(n_469) );
INVx2_ASAP7_75t_SL g470 ( .A(n_410), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_414), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_395), .A2(n_195), .B(n_154), .C(n_172), .Y(n_472) );
NOR3xp33_ASAP7_75t_L g473 ( .A(n_395), .B(n_195), .C(n_154), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_413), .A2(n_195), .B(n_154), .Y(n_474) );
NAND3xp33_ASAP7_75t_L g475 ( .A(n_387), .B(n_195), .C(n_154), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_375), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_375), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_413), .B(n_154), .Y(n_478) );
NOR2x1_ASAP7_75t_L g479 ( .A(n_375), .B(n_163), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_375), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_375), .B(n_154), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g482 ( .A1(n_390), .A2(n_192), .B1(n_343), .B2(n_244), .C(n_326), .Y(n_482) );
INVx1_ASAP7_75t_SL g483 ( .A(n_405), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_405), .B(n_192), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_375), .B(n_192), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_459), .A2(n_458), .B1(n_483), .B2(n_453), .Y(n_486) );
AOI221xp5_ASAP7_75t_L g487 ( .A1(n_482), .A2(n_454), .B1(n_422), .B2(n_476), .C(n_480), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_421), .A2(n_431), .B1(n_470), .B2(n_436), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_440), .B(n_443), .Y(n_489) );
AOI21xp33_ASAP7_75t_L g490 ( .A1(n_484), .A2(n_471), .B(n_469), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_452), .A2(n_442), .B(n_478), .Y(n_491) );
INVx2_ASAP7_75t_SL g492 ( .A(n_448), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_479), .Y(n_493) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_477), .A2(n_449), .B1(n_446), .B2(n_432), .C(n_438), .Y(n_494) );
AOI221xp5_ASAP7_75t_L g495 ( .A1(n_424), .A2(n_425), .B1(n_426), .B2(n_430), .C(n_441), .Y(n_495) );
OAI31xp33_ASAP7_75t_L g496 ( .A1(n_462), .A2(n_433), .A3(n_447), .B(n_472), .Y(n_496) );
BUFx2_ASAP7_75t_L g497 ( .A(n_429), .Y(n_497) );
XOR2xp5_ASAP7_75t_L g498 ( .A(n_466), .B(n_455), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_437), .Y(n_499) );
AOI21xp33_ASAP7_75t_L g500 ( .A1(n_428), .A2(n_481), .B(n_463), .Y(n_500) );
INVxp67_ASAP7_75t_L g501 ( .A(n_434), .Y(n_501) );
NAND4xp25_ASAP7_75t_L g502 ( .A(n_428), .B(n_473), .C(n_461), .D(n_423), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_489), .Y(n_503) );
NAND3xp33_ASAP7_75t_L g504 ( .A(n_488), .B(n_475), .C(n_457), .Y(n_504) );
AOI31xp33_ASAP7_75t_L g505 ( .A1(n_491), .A2(n_474), .A3(n_435), .B(n_464), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_499), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_501), .Y(n_507) );
INVx2_ASAP7_75t_SL g508 ( .A(n_486), .Y(n_508) );
OAI211xp5_ASAP7_75t_SL g509 ( .A1(n_487), .A2(n_435), .B(n_465), .C(n_456), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_497), .B(n_445), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_495), .B(n_468), .Y(n_511) );
AND4x1_ASAP7_75t_L g512 ( .A(n_504), .B(n_496), .C(n_494), .D(n_498), .Y(n_512) );
AOI211xp5_ASAP7_75t_L g513 ( .A1(n_508), .A2(n_502), .B(n_500), .C(n_496), .Y(n_513) );
NAND4xp25_ASAP7_75t_L g514 ( .A(n_504), .B(n_490), .C(n_493), .D(n_450), .Y(n_514) );
NAND3xp33_ASAP7_75t_SL g515 ( .A(n_511), .B(n_467), .C(n_460), .Y(n_515) );
NOR3xp33_ASAP7_75t_L g516 ( .A(n_505), .B(n_439), .C(n_492), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_514), .B(n_503), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_513), .A2(n_507), .B1(n_506), .B2(n_510), .Y(n_518) );
OR4x2_ASAP7_75t_L g519 ( .A(n_512), .B(n_509), .C(n_466), .D(n_439), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_517), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_518), .Y(n_521) );
OAI21x1_ASAP7_75t_L g522 ( .A1(n_520), .A2(n_519), .B(n_515), .Y(n_522) );
XNOR2xp5_ASAP7_75t_L g523 ( .A(n_521), .B(n_516), .Y(n_523) );
XOR2xp5_ASAP7_75t_L g524 ( .A(n_523), .B(n_444), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_524), .A2(n_522), .B1(n_427), .B2(n_485), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_525), .A2(n_522), .B(n_451), .Y(n_526) );
endmodule