module fake_ariane_279_n_71 (n_8, n_3, n_2, n_11, n_7, n_16, n_5, n_14, n_1, n_0, n_12, n_15, n_6, n_13, n_9, n_17, n_4, n_10, n_71);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_16;
input n_5;
input n_14;
input n_1;
input n_0;
input n_12;
input n_15;
input n_6;
input n_13;
input n_9;
input n_17;
input n_4;
input n_10;

output n_71;

wire n_66;
wire n_56;
wire n_60;
wire n_24;
wire n_22;
wire n_43;
wire n_49;
wire n_20;
wire n_27;
wire n_48;
wire n_29;
wire n_64;
wire n_41;
wire n_50;
wire n_38;
wire n_55;
wire n_62;
wire n_47;
wire n_18;
wire n_32;
wire n_28;
wire n_37;
wire n_58;
wire n_65;
wire n_51;
wire n_67;
wire n_45;
wire n_34;
wire n_69;
wire n_26;
wire n_46;
wire n_52;
wire n_36;
wire n_68;
wire n_33;
wire n_44;
wire n_19;
wire n_30;
wire n_39;
wire n_40;
wire n_59;
wire n_31;
wire n_42;
wire n_57;
wire n_63;
wire n_53;
wire n_21;
wire n_70;
wire n_23;
wire n_61;
wire n_35;
wire n_54;
wire n_25;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_6),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

AND2x4_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

AND2x4_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_20),
.A2(n_5),
.B(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

OAI21x1_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_19),
.B(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_28),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_36),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_19),
.B(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_22),
.Y(n_41)
);

OAI21x1_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_31),
.B(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_21),
.B1(n_29),
.B2(n_22),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_21),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_23),
.Y(n_51)
);

AND2x4_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_23),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_48),
.Y(n_56)
);

NOR2x1p5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_49),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_51),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_54),
.B(n_52),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_48),
.B(n_53),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NOR4xp25_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_58),
.C(n_57),
.D(n_53),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

NAND3x2_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_52),
.C(n_61),
.Y(n_65)
);

OAI22x1_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_62),
.B1(n_53),
.B2(n_4),
.Y(n_66)
);

AND4x1_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_60),
.C(n_25),
.D(n_27),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_67),
.B(n_25),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_65),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

OR2x6_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_68),
.Y(n_71)
);


endmodule