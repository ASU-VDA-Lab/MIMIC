module fake_jpeg_21506_n_249 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_249);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_10),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

FAx1_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_30),
.CI(n_27),
.CON(n_42),
.SN(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_21),
.B1(n_11),
.B2(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_21),
.B1(n_11),
.B2(n_23),
.Y(n_49)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_31),
.B1(n_38),
.B2(n_27),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_53),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_27),
.B(n_31),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_40),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_14),
.Y(n_71)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_65),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_34),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_17),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_18),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_78),
.B(n_79),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_75),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_54),
.C(n_26),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_63),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_31),
.B1(n_38),
.B2(n_57),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_82),
.B1(n_87),
.B2(n_91),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_28),
.B1(n_53),
.B2(n_43),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_86),
.B(n_89),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_28),
.B1(n_26),
.B2(n_37),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_28),
.B1(n_24),
.B2(n_26),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_73),
.B1(n_35),
.B2(n_24),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_63),
.A2(n_67),
.B1(n_60),
.B2(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_92),
.B(n_17),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_93),
.B(n_102),
.Y(n_120)
);

INVxp67_ASAP7_75t_SL g94 ( 
.A(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_94),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_76),
.A2(n_73),
.B(n_71),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_108),
.B(n_109),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_89),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_107),
.B(n_12),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_84),
.B(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_112),
.B(n_133),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_93),
.A2(n_85),
.B1(n_88),
.B2(n_79),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_134),
.B1(n_101),
.B2(n_103),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_85),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_124),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_129),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_105),
.A2(n_92),
.B(n_87),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_92),
.B1(n_28),
.B2(n_62),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_122),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_69),
.C(n_68),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_128),
.C(n_36),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_62),
.B1(n_26),
.B2(n_69),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_96),
.A2(n_33),
.B1(n_48),
.B2(n_46),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_72),
.B1(n_45),
.B2(n_52),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_68),
.C(n_33),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_95),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_59),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_55),
.Y(n_131)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_132),
.B(n_99),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_24),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_35),
.B1(n_33),
.B2(n_72),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_142),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_141),
.A2(n_123),
.B1(n_122),
.B2(n_119),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_100),
.B1(n_107),
.B2(n_33),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_143),
.A2(n_150),
.B1(n_121),
.B2(n_36),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_25),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_152),
.B1(n_40),
.B2(n_36),
.Y(n_167)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_24),
.B1(n_72),
.B2(n_40),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_120),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_113),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_40),
.B1(n_45),
.B2(n_29),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_12),
.Y(n_157)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_158),
.Y(n_170)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_162),
.A2(n_168),
.B1(n_148),
.B2(n_144),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_112),
.C(n_115),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_176),
.C(n_159),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_116),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_169),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_167),
.A2(n_141),
.B1(n_150),
.B2(n_137),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_138),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_172),
.B(n_154),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_13),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_173),
.B(n_159),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_32),
.C(n_29),
.Y(n_176)
);

NAND2xp33_ASAP7_75t_SL g178 ( 
.A(n_144),
.B(n_22),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_25),
.B(n_40),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_181),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_136),
.Y(n_180)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_189),
.B1(n_191),
.B2(n_194),
.Y(n_200)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_185),
.B(n_188),
.Y(n_206)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_186),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_187),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_143),
.C(n_152),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_140),
.B1(n_9),
.B2(n_10),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_140),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_13),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_193),
.A2(n_176),
.B1(n_174),
.B2(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_193),
.Y(n_196)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_202),
.Y(n_211)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_179),
.B(n_165),
.CI(n_170),
.CON(n_202),
.SN(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_182),
.A2(n_171),
.B1(n_170),
.B2(n_169),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_190),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_167),
.B(n_9),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_204),
.A2(n_8),
.B(n_10),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_181),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_210),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g209 ( 
.A(n_196),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_209),
.B(n_212),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_192),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_190),
.C(n_32),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_213),
.B(n_215),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_7),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_197),
.B(n_7),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_216),
.B(n_218),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_217),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_199),
.B(n_16),
.Y(n_218)
);

AOI211xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_200),
.B(n_202),
.C(n_201),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_219),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_207),
.B1(n_198),
.B2(n_32),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_220),
.A2(n_225),
.B1(n_226),
.B2(n_3),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_211),
.A2(n_198),
.B1(n_8),
.B2(n_2),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_0),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_32),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_221),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_229),
.B(n_230),
.Y(n_236)
);

INVxp67_ASAP7_75t_SL g231 ( 
.A(n_223),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_231),
.B(n_232),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_16),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_224),
.B(n_3),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_234),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_225),
.A2(n_25),
.B(n_16),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_235),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_SL g238 ( 
.A1(n_228),
.A2(n_22),
.B(n_4),
.C(n_5),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_238),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_242)
);

NOR2x1_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_230),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_241),
.A2(n_242),
.B(n_243),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_29),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_241),
.A2(n_239),
.B(n_237),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_245),
.A2(n_29),
.B(n_5),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_246),
.A2(n_244),
.B(n_5),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_3),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_6),
.B(n_236),
.Y(n_249)
);


endmodule