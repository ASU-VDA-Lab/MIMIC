module fake_ariane_206_n_189 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_189);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_189;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_156;
wire n_96;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_178;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_188;
wire n_185;
wire n_32;
wire n_58;
wire n_37;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_29;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_146;
wire n_80;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVxp67_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVxp67_ASAP7_75t_SL g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

INVxp67_ASAP7_75t_SL g37 ( 
.A(n_15),
.Y(n_37)
);

INVxp33_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_3),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2x1p5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

OAI221xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_35),
.B1(n_30),
.B2(n_33),
.C(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_49),
.Y(n_82)
);

OAI221xp5_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_47),
.B1(n_29),
.B2(n_37),
.C(n_36),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_38),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_47),
.B1(n_44),
.B2(n_8),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_57),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_63),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_84),
.B(n_56),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_64),
.B1(n_56),
.B2(n_69),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_63),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_70),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_72),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_70),
.B1(n_68),
.B2(n_65),
.Y(n_100)
);

AND2x4_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_82),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_75),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_63),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_98),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_83),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_91),
.Y(n_111)
);

OR2x6_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_97),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_90),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

NAND2xp33_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_107),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_102),
.B(n_103),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_93),
.B1(n_110),
.B2(n_113),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_90),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

AND2x4_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_112),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_93),
.C(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_124),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_108),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_121),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_112),
.B1(n_101),
.B2(n_68),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_130),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_125),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_122),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_138),
.Y(n_147)
);

NAND2x1p5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_115),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_77),
.B(n_60),
.C(n_61),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_53),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_52),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_51),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_112),
.B1(n_101),
.B2(n_105),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_145),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_62),
.C(n_66),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_144),
.B1(n_148),
.B2(n_97),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_154),
.A2(n_144),
.B1(n_148),
.B2(n_97),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_96),
.C(n_102),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_115),
.B(n_109),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_153),
.C(n_155),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_8),
.Y(n_168)
);

AOI221xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_150),
.B1(n_81),
.B2(n_78),
.C(n_79),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_9),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_75),
.B1(n_128),
.B2(n_87),
.Y(n_171)
);

OAI22x1_ASAP7_75t_SL g172 ( 
.A1(n_163),
.A2(n_80),
.B1(n_105),
.B2(n_94),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_96),
.C(n_89),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_SL g174 ( 
.A(n_164),
.B(n_100),
.C(n_94),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_166),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_170),
.Y(n_176)
);

AO22x2_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_101),
.B1(n_109),
.B2(n_86),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_174),
.A2(n_101),
.B1(n_88),
.B2(n_128),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_88),
.B1(n_104),
.B2(n_106),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_175),
.B(n_106),
.Y(n_180)
);

AOI211xp5_ASAP7_75t_L g181 ( 
.A1(n_167),
.A2(n_99),
.B(n_106),
.C(n_104),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_176),
.A2(n_171),
.B(n_173),
.C(n_169),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_177),
.A2(n_106),
.B1(n_99),
.B2(n_13),
.Y(n_183)
);

OAI22x1_ASAP7_75t_L g184 ( 
.A1(n_179),
.A2(n_10),
.B1(n_12),
.B2(n_17),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_180),
.A2(n_99),
.B1(n_20),
.B2(n_22),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_181),
.B1(n_178),
.B2(n_99),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_99),
.C(n_26),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_186),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_187),
.B1(n_184),
.B2(n_185),
.Y(n_189)
);


endmodule