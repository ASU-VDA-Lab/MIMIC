module real_jpeg_9436_n_18 (n_17, n_8, n_0, n_2, n_284, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_284;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_80;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_1),
.A2(n_46),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_1),
.B(n_46),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_1),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_1),
.A2(n_73),
.B1(n_76),
.B2(n_135),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_1),
.A2(n_32),
.B(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_1),
.B(n_32),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_1),
.B(n_181),
.Y(n_180)
);

AOI21xp33_ASAP7_75t_L g200 ( 
.A1(n_1),
.A2(n_29),
.B(n_33),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_1),
.A2(n_26),
.B1(n_35),
.B2(n_137),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_2),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_2),
.A2(n_58),
.B1(n_59),
.B2(n_126),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_126),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_2),
.A2(n_26),
.B1(n_35),
.B2(n_126),
.Y(n_222)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_5),
.A2(n_50),
.B1(n_58),
.B2(n_59),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_7),
.A2(n_26),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_7),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_7),
.A2(n_38),
.B1(n_58),
.B2(n_59),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_SL g55 ( 
.A1(n_8),
.A2(n_46),
.B(n_56),
.C(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_8),
.B(n_46),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_52),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_11),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_13),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_117),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_117),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_13),
.A2(n_26),
.B1(n_35),
.B2(n_117),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_14),
.A2(n_26),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_14),
.A2(n_36),
.B1(n_58),
.B2(n_59),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_14),
.A2(n_36),
.B1(n_46),
.B2(n_47),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_16),
.A2(n_26),
.B1(n_35),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_16),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_16),
.A2(n_58),
.B1(n_59),
.B2(n_100),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_16),
.A2(n_46),
.B1(n_47),
.B2(n_100),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_100),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_17),
.A2(n_26),
.B1(n_35),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_17),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_17),
.A2(n_58),
.B1(n_59),
.B2(n_83),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_17),
.A2(n_46),
.B1(n_47),
.B2(n_83),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_83),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_84),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_21),
.B(n_84),
.Y(n_105)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_21),
.Y(n_283)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_64),
.CI(n_69),
.CON(n_21),
.SN(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_39),
.B2(n_40),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_25),
.A2(n_31),
.B1(n_34),
.B2(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_25),
.A2(n_31),
.B1(n_82),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_25),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_25),
.A2(n_31),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_25),
.A2(n_31),
.B1(n_99),
.B2(n_234),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_28),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_26),
.A2(n_28),
.B(n_137),
.C(n_200),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_31),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_43),
.Y(n_44)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_53),
.B1(n_54),
.B2(n_63),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_45),
.B1(n_49),
.B2(n_51),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_45),
.B1(n_49),
.B2(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_42),
.A2(n_45),
.B1(n_66),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_42),
.A2(n_45),
.B1(n_159),
.B2(n_161),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_42),
.A2(n_45),
.B1(n_161),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_42),
.A2(n_45),
.B1(n_177),
.B2(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_42),
.A2(n_45),
.B1(n_218),
.B2(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_42),
.A2(n_45),
.B1(n_103),
.B2(n_230),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_44),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_45),
.B(n_137),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_46),
.B(n_48),
.Y(n_165)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_47),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_57),
.B(n_61),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_55),
.A2(n_57),
.B1(n_61),
.B2(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_55),
.A2(n_57),
.B1(n_68),
.B2(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_55),
.A2(n_57),
.B1(n_79),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_55),
.A2(n_57),
.B1(n_123),
.B2(n_125),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_55),
.A2(n_57),
.B1(n_125),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_55),
.A2(n_57),
.B1(n_150),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_55),
.A2(n_57),
.B1(n_157),
.B2(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_55),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_55),
.A2(n_57),
.B1(n_96),
.B2(n_240),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_57),
.B(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_57),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_58),
.B(n_60),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_58),
.B(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_59),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_65),
.B(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_80),
.B(n_81),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_71),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_72),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_80),
.B1(n_81),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_72),
.A2(n_78),
.B1(n_80),
.B2(n_265),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_76),
.B(n_77),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_76),
.B1(n_77),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_73),
.A2(n_76),
.B1(n_116),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_73),
.A2(n_76),
.B1(n_119),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_73),
.A2(n_76),
.B1(n_152),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_73),
.A2(n_76),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_73),
.A2(n_76),
.B1(n_94),
.B2(n_204),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_74),
.A2(n_75),
.B1(n_115),
.B2(n_118),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_74),
.A2(n_75),
.B1(n_169),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_76),
.B(n_137),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_78),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.C(n_90),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_85),
.B(n_89),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_90),
.A2(n_91),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.C(n_101),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_92),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_93),
.B(n_95),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_102),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI321xp33_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_259),
.A3(n_270),
.B1(n_276),
.B2(n_281),
.C(n_284),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_224),
.C(n_255),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_193),
.B(n_223),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_171),
.B(n_192),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_154),
.B(n_170),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_144),
.B(n_153),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_132),
.B(n_143),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_120),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_114),
.B(n_120),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_127),
.B2(n_131),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_121),
.B(n_131),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_124),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_127),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_138),
.B(n_142),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_136),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_145),
.B(n_146),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_147),
.B(n_155),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_149),
.CI(n_151),
.CON(n_147),
.SN(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_155),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_158),
.CI(n_162),
.CON(n_155),
.SN(n_155)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_160),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_167),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_172),
.B(n_173),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_185),
.B2(n_186),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_188),
.C(n_190),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_178),
.B1(n_179),
.B2(n_184),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_176),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_182),
.C(n_184),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_181),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_183),
.Y(n_203)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_187),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_188),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_189),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_194),
.B(n_195),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_208),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_197),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_197),
.B(n_207),
.C(n_208),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_202),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_205),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_219),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_216),
.B2(n_217),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_216),
.C(n_219),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_214),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_222),
.Y(n_233)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g277 ( 
.A1(n_225),
.A2(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_242),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_226),
.B(n_242),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_237),
.C(n_241),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_236),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_231),
.B1(n_232),
.B2(n_235),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_229),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_SL g253 ( 
.A(n_231),
.B(n_235),
.C(n_236),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_241),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_239),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_253),
.B2(n_254),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_246),
.C(n_254),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_250),
.C(n_252),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_249),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_253),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_257),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_260),
.B(n_267),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.C(n_266),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_264),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_271),
.A2(n_277),
.B(n_280),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_272),
.B(n_273),
.Y(n_280)
);


endmodule