module fake_jpeg_7899_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_6),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_19),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_0),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_47),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_24),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_47),
.A2(n_26),
.B1(n_33),
.B2(n_23),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_53),
.B1(n_71),
.B2(n_74),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_33),
.B1(n_16),
.B2(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_62),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_66),
.Y(n_99)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_19),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_72),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_70),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_33),
.B1(n_26),
.B2(n_23),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_18),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_16),
.B1(n_23),
.B2(n_26),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_16),
.B1(n_24),
.B2(n_17),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_17),
.B1(n_24),
.B2(n_16),
.Y(n_101)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_77),
.Y(n_104)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_72),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_78),
.B(n_79),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_38),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_81),
.Y(n_123)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_85),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_41),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_87),
.B(n_88),
.Y(n_137)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_50),
.A2(n_41),
.B(n_20),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_93),
.A2(n_94),
.B(n_100),
.C(n_21),
.Y(n_142)
);

OR2x4_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_48),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_54),
.B(n_28),
.Y(n_95)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_30),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_22),
.B(n_27),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_34),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_110),
.Y(n_126)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_30),
.B(n_48),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_101),
.A2(n_113),
.B1(n_116),
.B2(n_46),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_24),
.B1(n_17),
.B2(n_30),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_103),
.A2(n_17),
.B1(n_22),
.B2(n_27),
.Y(n_133)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_55),
.B(n_32),
.Y(n_109)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_34),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_48),
.C(n_44),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_46),
.C(n_36),
.Y(n_127)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_40),
.Y(n_132)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

FAx1_ASAP7_75t_SL g117 ( 
.A(n_89),
.B(n_60),
.CI(n_48),
.CON(n_117),
.SN(n_117)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_117),
.B(n_96),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_118),
.A2(n_144),
.B1(n_112),
.B2(n_108),
.Y(n_170)
);

NOR2x1_ASAP7_75t_R g119 ( 
.A(n_94),
.B(n_48),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_111),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_104),
.B1(n_82),
.B2(n_115),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_131),
.B1(n_135),
.B2(n_142),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_147),
.C(n_46),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_80),
.A2(n_40),
.B1(n_27),
.B2(n_34),
.Y(n_131)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_143),
.B1(n_25),
.B2(n_107),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_88),
.A2(n_22),
.B1(n_31),
.B2(n_29),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_97),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_145),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_99),
.A2(n_31),
.B1(n_32),
.B2(n_28),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_31),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_31),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_114),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_93),
.B(n_44),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_123),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_148),
.B(n_155),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_149),
.A2(n_153),
.B(n_146),
.Y(n_191)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_152),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_151),
.A2(n_170),
.B1(n_14),
.B2(n_7),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_141),
.B(n_25),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_100),
.B1(n_98),
.B2(n_105),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_156),
.A2(n_167),
.B1(n_172),
.B2(n_176),
.Y(n_192)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_163),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_159),
.C(n_165),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_106),
.C(n_55),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_55),
.C(n_92),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_166),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_112),
.B1(n_108),
.B2(n_84),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_122),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_168),
.B(n_169),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_129),
.B(n_85),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_126),
.B(n_86),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g208 ( 
.A(n_171),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_84),
.B1(n_113),
.B2(n_25),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_122),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_173),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_0),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_178),
.Y(n_183)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_175),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_92),
.B1(n_2),
.B2(n_4),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_177),
.A2(n_143),
.B1(n_120),
.B2(n_135),
.Y(n_196)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_8),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_179),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_14),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_181),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_147),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_202),
.C(n_212),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_189),
.B(n_198),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_117),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_190),
.B(n_11),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_191),
.A2(n_201),
.B(n_149),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_137),
.Y(n_194)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_196),
.A2(n_209),
.B1(n_211),
.B2(n_185),
.Y(n_242)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_161),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_200),
.B(n_204),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_178),
.A2(n_127),
.B1(n_118),
.B2(n_121),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_133),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_156),
.A2(n_130),
.B1(n_121),
.B2(n_124),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_124),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_211),
.Y(n_217)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_7),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_6),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_177),
.C(n_151),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_226),
.C(n_240),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_201),
.A2(n_154),
.B1(n_149),
.B2(n_166),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_219),
.A2(n_224),
.B1(n_184),
.B2(n_206),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_193),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_220),
.B(n_228),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_216),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_176),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_223),
.A2(n_237),
.B(n_183),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_189),
.A2(n_175),
.B1(n_150),
.B2(n_4),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_1),
.C(n_2),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_188),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_227),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_210),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_222),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_231),
.A2(n_234),
.B1(n_241),
.B2(n_242),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_207),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_232),
.Y(n_263)
);

AO22x1_ASAP7_75t_SL g233 ( 
.A1(n_192),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_233),
.A2(n_194),
.B1(n_185),
.B2(n_191),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_198),
.A2(n_5),
.B1(n_11),
.B2(n_12),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_199),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_236),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_4),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_215),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_12),
.C(n_13),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_192),
.A2(n_13),
.B1(n_183),
.B2(n_196),
.Y(n_241)
);

INVxp33_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_243),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_246),
.B(n_254),
.Y(n_280)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_248),
.A2(n_251),
.B(n_260),
.Y(n_268)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_195),
.C(n_190),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_235),
.C(n_240),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_230),
.A2(n_187),
.B1(n_212),
.B2(n_184),
.Y(n_257)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_233),
.A2(n_186),
.B1(n_214),
.B2(n_208),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_261),
.B(n_218),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_219),
.A2(n_203),
.B(n_186),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_223),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_221),
.Y(n_270)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_223),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_243),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_258),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_272),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_247),
.Y(n_269)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_274),
.C(n_275),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_238),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_235),
.C(n_226),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_254),
.C(n_246),
.Y(n_278)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_229),
.C(n_237),
.Y(n_279)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_263),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_229),
.C(n_237),
.Y(n_284)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_268),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_301),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_265),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_261),
.B(n_266),
.Y(n_296)
);

NAND2xp33_ASAP7_75t_SL g306 ( 
.A(n_296),
.B(n_272),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_285),
.A2(n_242),
.B1(n_245),
.B2(n_233),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_302),
.B1(n_252),
.B2(n_280),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_281),
.A2(n_245),
.B(n_251),
.Y(n_299)
);

MAJx2_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_296),
.C(n_273),
.Y(n_303)
);

BUFx12_ASAP7_75t_L g301 ( 
.A(n_269),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_276),
.A2(n_260),
.B1(n_248),
.B2(n_259),
.Y(n_302)
);

AO21x1_ASAP7_75t_L g318 ( 
.A1(n_303),
.A2(n_306),
.B(n_300),
.Y(n_318)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_299),
.B(n_284),
.CI(n_280),
.CON(n_304),
.SN(n_304)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_309),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_282),
.Y(n_305)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_305),
.Y(n_316)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_278),
.C(n_275),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_310),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_301),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_244),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_314),
.Y(n_317)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_315),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_302),
.B(n_274),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_298),
.B(n_264),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_320),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_303),
.A2(n_291),
.B1(n_297),
.B2(n_294),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_270),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_293),
.C(n_288),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_288),
.C(n_277),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_326),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_322),
.A2(n_305),
.B(n_301),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_316),
.A2(n_304),
.B1(n_244),
.B2(n_311),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_327),
.B(n_321),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_279),
.C(n_319),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_SL g330 ( 
.A(n_318),
.B(n_317),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_330),
.B(n_331),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_324),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_337),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_317),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_338),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_332),
.C(n_333),
.Y(n_340)
);

INVxp33_ASAP7_75t_L g341 ( 
.A(n_340),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_328),
.Y(n_342)
);


endmodule