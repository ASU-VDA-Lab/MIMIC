module real_jpeg_23012_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_0),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_0),
.B(n_17),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_0),
.B(n_93),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_0),
.B(n_51),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_0),
.B(n_54),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_0),
.B(n_37),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_0),
.B(n_30),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_0),
.B(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_2),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_3),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_3),
.B(n_86),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_3),
.B(n_93),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_3),
.B(n_51),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_3),
.B(n_54),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_3),
.B(n_37),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_3),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_3),
.B(n_196),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_4),
.B(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_4),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_4),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_4),
.B(n_93),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_5),
.B(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_30),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_5),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_5),
.B(n_86),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_5),
.B(n_93),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_5),
.B(n_51),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_5),
.B(n_54),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_5),
.B(n_37),
.Y(n_366)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_8),
.B(n_51),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_8),
.B(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_8),
.B(n_54),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_8),
.B(n_37),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_8),
.B(n_30),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_9),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_9),
.B(n_86),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_9),
.B(n_93),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_9),
.B(n_51),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_9),
.B(n_54),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_9),
.B(n_37),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_9),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_9),
.B(n_253),
.Y(n_325)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_11),
.B(n_24),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_11),
.B(n_117),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_11),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_11),
.B(n_93),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_11),
.B(n_51),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_11),
.B(n_54),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_11),
.B(n_37),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_11),
.B(n_30),
.Y(n_365)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_13),
.B(n_17),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_13),
.B(n_86),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_13),
.B(n_93),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_13),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_13),
.B(n_37),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_13),
.B(n_30),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_13),
.B(n_253),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_15),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_15),
.B(n_86),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_15),
.B(n_93),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_15),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_15),
.B(n_54),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_15),
.B(n_37),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_16),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_16),
.B(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_16),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_16),
.B(n_51),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_16),
.B(n_54),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_16),
.B(n_37),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_16),
.B(n_30),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_16),
.B(n_24),
.Y(n_235)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_17),
.Y(n_108)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_17),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_65),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_41),
.B2(n_42),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_35),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_27),
.Y(n_196)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_27),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_36),
.C(n_40),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_28),
.A2(n_34),
.B1(n_36),
.B2(n_59),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_29),
.B(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_29),
.B(n_281),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_29),
.B(n_244),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_32),
.B(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_32),
.B(n_232),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_62),
.C(n_63),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_43),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_43),
.B(n_382),
.Y(n_381)
);

FAx1_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_45),
.CI(n_55),
.CON(n_43),
.SN(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.C(n_53),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_46),
.A2(n_47),
.B1(n_371),
.B2(n_372),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_49),
.A2(n_311),
.B1(n_312),
.B2(n_339),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_49),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_SL g369 ( 
.A(n_49),
.B(n_312),
.C(n_337),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_49),
.A2(n_53),
.B1(n_58),
.B2(n_339),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_50),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_50),
.B(n_244),
.Y(n_243)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_53),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_59),
.C(n_61),
.Y(n_62)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_54),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_60),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_62),
.B(n_63),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_381),
.C(n_383),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_376),
.C(n_377),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_358),
.C(n_359),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_329),
.C(n_330),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_304),
.C(n_305),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_273),
.C(n_274),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_237),
.C(n_238),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_202),
.C(n_203),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_170),
.C(n_171),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_148),
.C(n_149),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_130),
.C(n_131),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_109),
.C(n_110),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_95),
.C(n_100),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_89),
.B2(n_90),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_91),
.C(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_84),
.B1(n_85),
.B2(n_88),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_86),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.C(n_104),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_103),
.B(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_108),
.B(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_121),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_115),
.C(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_116),
.Y(n_120)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_117),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_118),
.B(n_120),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_129),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_122),
.Y(n_129)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_125),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_128),
.C(n_129),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_139),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_134),
.C(n_139),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_137),
.C(n_138),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_142),
.C(n_143),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_147),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_164),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_165),
.C(n_169),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_160),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_159),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_159),
.C(n_160),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_153),
.Y(n_158)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_158),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g386 ( 
.A(n_160),
.Y(n_386)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_162),
.CI(n_163),
.CON(n_160),
.SN(n_160)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_162),
.C(n_163),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_165),
.Y(n_187)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_167),
.CI(n_168),
.CON(n_165),
.SN(n_165)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_186),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_175),
.C(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_182),
.C(n_185),
.Y(n_206)
);

BUFx24_ASAP7_75t_SL g385 ( 
.A(n_177),
.Y(n_385)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_179),
.CI(n_180),
.CON(n_177),
.SN(n_177)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_179),
.C(n_180),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_193),
.C(n_200),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_193),
.B1(n_200),
.B2(n_201),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_189),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B(n_192),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_191),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_192),
.B(n_227),
.C(n_228),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_193),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_198),
.C(n_199),
.Y(n_222)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_223),
.B2(n_236),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_224),
.C(n_225),
.Y(n_237)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_208),
.C(n_216),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_216),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_212),
.C(n_215),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_214),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_221),
.C(n_222),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_220),
.Y(n_221)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_235),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_233),
.C(n_235),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_271),
.B2(n_272),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_239),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_262),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_262),
.C(n_271),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_249),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_242),
.B(n_250),
.C(n_251),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g389 ( 
.A(n_242),
.Y(n_389)
);

FAx1_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_245),
.CI(n_247),
.CON(n_242),
.SN(n_242)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_243),
.B(n_245),
.C(n_247),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_254),
.B1(n_255),
.B2(n_261),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_252),
.Y(n_261)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_256),
.A2(n_257),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_260),
.C(n_261),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_256),
.B(n_280),
.C(n_283),
.Y(n_327)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_265),
.C(n_266),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_269),
.C(n_270),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_277),
.C(n_303),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_291),
.B2(n_303),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_285),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_279),
.B(n_286),
.C(n_287),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_283),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_283),
.A2(n_284),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_SL g343 ( 
.A(n_283),
.B(n_309),
.C(n_312),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g388 ( 
.A(n_287),
.Y(n_388)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_289),
.CI(n_290),
.CON(n_287),
.SN(n_287)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_289),
.C(n_290),
.Y(n_314)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g387 ( 
.A(n_291),
.Y(n_387)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.CI(n_294),
.CON(n_291),
.SN(n_291)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_293),
.C(n_294),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_302),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_295),
.B(n_298),
.C(n_300),
.Y(n_322)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_297),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_298),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_299),
.A2(n_300),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_326),
.C(n_327),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_328),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_319),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_319),
.C(n_328),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_308),
.B(n_314),
.C(n_315),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g384 ( 
.A(n_315),
.Y(n_384)
);

FAx1_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_317),
.CI(n_318),
.CON(n_315),
.SN(n_315)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_317),
.C(n_318),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_322),
.C(n_323),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_327),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_325),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_331),
.B(n_333),
.C(n_345),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_344),
.B2(n_345),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_336),
.B1(n_340),
.B2(n_341),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_335),
.B(n_342),
.C(n_343),
.Y(n_361)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_346),
.B(n_348),
.C(n_351),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_348),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_351),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_354),
.C(n_357),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_355),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_356),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_373),
.B1(n_374),
.B2(n_375),
.Y(n_359)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_360),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_361),
.B(n_362),
.C(n_375),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_368),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_363),
.B(n_369),
.C(n_370),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_364),
.B(n_380),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_364),
.B(n_378),
.C(n_380),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g364 ( 
.A(n_365),
.B(n_366),
.CI(n_367),
.CON(n_364),
.SN(n_364)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_371),
.Y(n_372)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_373),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);


endmodule