module fake_netlist_5_1605_n_184 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_30, n_20, n_5, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_184);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;

output n_184;

wire n_137;
wire n_168;
wire n_164;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_176;
wire n_140;
wire n_124;
wire n_86;
wire n_136;
wire n_146;
wire n_182;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_180;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_179;
wire n_125;
wire n_35;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_151;
wire n_131;
wire n_47;
wire n_173;
wire n_53;
wire n_160;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_154;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_183;
wire n_175;
wire n_169;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_181;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_178;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_162;
wire n_170;
wire n_64;
wire n_102;
wire n_77;
wire n_106;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_174;
wire n_134;
wire n_32;
wire n_41;
wire n_104;
wire n_172;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_141;
wire n_166;
wire n_171;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVxp67_ASAP7_75t_SL g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_0),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_1),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_1),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_7),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_32),
.B(n_7),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NAND2x1p5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_51),
.Y(n_78)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_55),
.B1(n_60),
.B2(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

AO22x2_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_53),
.B1(n_47),
.B2(n_44),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_39),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_52),
.B(n_49),
.C(n_37),
.Y(n_86)
);

AND2x4_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_49),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_8),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_37),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_87),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_46),
.C(n_64),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_67),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_63),
.B1(n_66),
.B2(n_74),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_73),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_79),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_75),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_79),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_82),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_77),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_109),
.A2(n_100),
.B(n_99),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_82),
.Y(n_114)
);

NOR2x1_ASAP7_75t_SL g115 ( 
.A(n_109),
.B(n_102),
.Y(n_115)
);

NOR2x1_ASAP7_75t_SL g116 ( 
.A(n_106),
.B(n_97),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_97),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_108),
.B(n_104),
.C(n_111),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

AO21x2_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_110),
.B(n_105),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_121),
.A2(n_112),
.B1(n_117),
.B2(n_104),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_114),
.B1(n_107),
.B2(n_82),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_115),
.B(n_116),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_122),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_77),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_130),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_114),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_114),
.B1(n_89),
.B2(n_96),
.Y(n_139)
);

NOR2x1_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_118),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_129),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_87),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_125),
.B1(n_96),
.B2(n_101),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_126),
.Y(n_144)
);

NAND2x1_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_126),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_139),
.B(n_128),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_133),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_131),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_143),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_101),
.C(n_94),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_153),
.A2(n_127),
.B(n_131),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_115),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_90),
.B(n_110),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_155),
.A2(n_61),
.B(n_9),
.Y(n_167)
);

XNOR2x1_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_8),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_160),
.C(n_157),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_156),
.Y(n_170)
);

OAI221xp5_ASAP7_75t_L g171 ( 
.A1(n_162),
.A2(n_61),
.B1(n_73),
.B2(n_71),
.C(n_69),
.Y(n_171)
);

OA211x2_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_9),
.B(n_116),
.C(n_11),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_71),
.Y(n_173)
);

NAND4xp75_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_163),
.C(n_103),
.D(n_91),
.Y(n_174)
);

OAI211xp5_ASAP7_75t_SL g175 ( 
.A1(n_169),
.A2(n_61),
.B(n_103),
.C(n_85),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_59),
.C(n_118),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_173),
.A2(n_59),
.B1(n_12),
.B2(n_14),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_10),
.B(n_16),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_171),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_21),
.Y(n_180)
);

NAND4xp25_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_24),
.C(n_26),
.D(n_59),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_180),
.A2(n_178),
.B1(n_174),
.B2(n_59),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_179),
.B1(n_181),
.B2(n_59),
.Y(n_184)
);


endmodule