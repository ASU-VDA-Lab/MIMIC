module real_jpeg_4584_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_487;
wire n_242;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx5_ASAP7_75t_L g185 ( 
.A(n_0),
.Y(n_185)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_0),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_0),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_0),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_0),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g324 ( 
.A(n_1),
.Y(n_324)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_1),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_1),
.Y(n_399)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_2),
.A2(n_175),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_2),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_2),
.A2(n_178),
.B1(n_259),
.B2(n_261),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_2),
.A2(n_100),
.B1(n_178),
.B2(n_360),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_2),
.A2(n_178),
.B1(n_323),
.B2(n_399),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_3),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_3),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_3),
.A2(n_209),
.B1(n_228),
.B2(n_232),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_3),
.A2(n_91),
.B1(n_209),
.B2(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_3),
.A2(n_65),
.B1(n_209),
.B2(n_419),
.Y(n_418)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g328 ( 
.A(n_4),
.Y(n_328)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_6),
.A2(n_91),
.B1(n_93),
.B2(n_95),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_6),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_6),
.A2(n_60),
.B1(n_95),
.B2(n_134),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_6),
.A2(n_95),
.B1(n_229),
.B2(n_378),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_6),
.A2(n_95),
.B1(n_404),
.B2(n_405),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_7),
.A2(n_86),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_7),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_7),
.A2(n_161),
.B1(n_195),
.B2(n_199),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_7),
.A2(n_93),
.B1(n_161),
.B2(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_7),
.A2(n_161),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_8),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_8),
.Y(n_117)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_8),
.Y(n_122)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_9),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_10),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_10),
.Y(n_127)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_10),
.Y(n_189)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_13),
.A2(n_153),
.B1(n_156),
.B2(n_158),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_13),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_13),
.B(n_117),
.C(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_13),
.B(n_81),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_13),
.B(n_185),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_13),
.B(n_165),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_13),
.B(n_94),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_14),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_14),
.A2(n_56),
.B1(n_220),
.B2(n_308),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_14),
.A2(n_56),
.B1(n_283),
.B2(n_386),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_14),
.A2(n_56),
.B1(n_395),
.B2(n_396),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_15),
.A2(n_98),
.B1(n_100),
.B2(n_104),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_15),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_15),
.A2(n_104),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_15),
.A2(n_104),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_15),
.A2(n_104),
.B1(n_382),
.B2(n_383),
.Y(n_381)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_17),
.A2(n_176),
.B1(n_228),
.B2(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_17),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_17),
.A2(n_277),
.B1(n_365),
.B2(n_367),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_17),
.A2(n_277),
.B1(n_391),
.B2(n_393),
.Y(n_390)
);

OAI22xp33_ASAP7_75t_L g446 ( 
.A1(n_17),
.A2(n_65),
.B1(n_140),
.B2(n_277),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_18),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_18),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_18),
.A2(n_66),
.B1(n_123),
.B2(n_340),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_18),
.A2(n_66),
.B1(n_154),
.B2(n_365),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_18),
.A2(n_66),
.B1(n_265),
.B2(n_433),
.Y(n_432)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_522),
.B(n_525),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_142),
.B(n_521),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_138),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_27),
.B(n_138),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_132),
.C(n_135),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_28),
.A2(n_29),
.B1(n_517),
.B2(n_518),
.Y(n_516)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_67),
.C(n_105),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g508 ( 
.A(n_30),
.B(n_509),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_51),
.B1(n_57),
.B2(n_59),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_31),
.A2(n_57),
.B1(n_59),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_31),
.A2(n_57),
.B1(n_133),
.B2(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_31),
.A2(n_351),
.B(n_398),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_31),
.A2(n_57),
.B1(n_398),
.B2(n_418),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_31),
.A2(n_51),
.B1(n_57),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_32),
.A2(n_347),
.B(n_350),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_32),
.B(n_352),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_32),
.A2(n_58),
.B(n_524),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_42),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_35),
.Y(n_325)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_36),
.Y(n_134)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_38),
.Y(n_353)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_50),
.Y(n_42)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_45),
.Y(n_322)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_46),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_46),
.Y(n_395)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_49),
.Y(n_331)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_54),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_57),
.B(n_158),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_57),
.A2(n_418),
.B(n_447),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_58),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_58),
.B(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_64),
.Y(n_356)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_65),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_65),
.B(n_158),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_67),
.A2(n_105),
.B1(n_106),
.B2(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_67),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_90),
.B1(n_96),
.B2(n_97),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_68),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_68),
.A2(n_96),
.B1(n_298),
.B2(n_359),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_68),
.A2(n_96),
.B1(n_390),
.B2(n_394),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_68),
.A2(n_90),
.B1(n_96),
.B2(n_498),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_81),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_74),
.B1(n_76),
.B2(n_79),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_72),
.Y(n_281)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g362 ( 
.A(n_75),
.Y(n_362)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_78),
.Y(n_287)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_81),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_81),
.A2(n_136),
.B(n_137),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_81),
.A2(n_136),
.B1(n_303),
.B2(n_423),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_81),
.A2(n_136),
.B1(n_431),
.B2(n_432),
.Y(n_430)
);

AO22x2_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_88),
.Y(n_81)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_83),
.Y(n_168)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_83),
.Y(n_208)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_84),
.Y(n_260)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_85),
.Y(n_164)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_85),
.Y(n_406)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_87),
.Y(n_212)
);

INVx6_ASAP7_75t_L g368 ( 
.A(n_87),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_87),
.Y(n_404)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_91),
.Y(n_434)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_96),
.B(n_271),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_96),
.A2(n_298),
.B(n_302),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_98),
.Y(n_393)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_100),
.Y(n_272)
);

AOI32xp33_ASAP7_75t_L g278 ( 
.A1(n_100),
.A2(n_259),
.A3(n_269),
.B1(n_279),
.B2(n_282),
.Y(n_278)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_103),
.Y(n_267)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_103),
.Y(n_392)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_103),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_105),
.A2(n_106),
.B1(n_496),
.B2(n_497),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_105),
.B(n_493),
.C(n_496),
.Y(n_504)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_119),
.B(n_128),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_152),
.B(n_159),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_107),
.A2(n_119),
.B1(n_206),
.B2(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_107),
.A2(n_159),
.B(n_258),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_107),
.A2(n_119),
.B1(n_364),
.B2(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_108),
.B(n_160),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_108),
.A2(n_165),
.B1(n_385),
.B2(n_387),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_108),
.A2(n_165),
.B1(n_387),
.B2(n_403),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_108),
.A2(n_165),
.B1(n_403),
.B2(n_437),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_119),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B1(n_116),
.B2(n_118),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_112),
.Y(n_261)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22x1_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_120),
.B1(n_123),
.B2(n_126),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_119),
.A2(n_206),
.B(n_213),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_119),
.A2(n_213),
.B(n_364),
.Y(n_363)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

BUFx8_ASAP7_75t_L g222 ( 
.A(n_125),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_127),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_127),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_127),
.Y(n_382)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_128),
.Y(n_437)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_131),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_132),
.B(n_135),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_136),
.A2(n_264),
.B(n_270),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_136),
.B(n_303),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_136),
.A2(n_270),
.B(n_460),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_138),
.B(n_523),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_138),
.B(n_523),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_139),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_515),
.B(n_520),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_487),
.B(n_512),
.Y(n_143)
);

OAI311xp33_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_371),
.A3(n_463),
.B1(n_481),
.C1(n_486),
.Y(n_144)
);

AOI21x1_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_313),
.B(n_370),
.Y(n_145)
);

AO21x1_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_289),
.B(n_312),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_252),
.B(n_288),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_216),
.B(n_251),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_172),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_150),
.B(n_172),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_166),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_151),
.A2(n_166),
.B1(n_167),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_151),
.Y(n_249)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_155),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_155),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_158),
.A2(n_183),
.B(n_190),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_SL g264 ( 
.A1(n_158),
.A2(n_265),
.B(n_268),
.Y(n_264)
);

OAI21xp33_ASAP7_75t_SL g347 ( 
.A1(n_158),
.A2(n_332),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_165),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_203),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_173),
.B(n_204),
.C(n_215),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_183),
.B(n_190),
.Y(n_173)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_182),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_183),
.A2(n_335),
.B1(n_336),
.B2(n_338),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_183),
.A2(n_246),
.B1(n_377),
.B2(n_381),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_183),
.A2(n_192),
.B(n_381),
.Y(n_407)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_184),
.B(n_194),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_184),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_184),
.A2(n_276),
.B1(n_307),
.B2(n_309),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_184),
.A2(n_339),
.B1(n_414),
.B2(n_415),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_196),
.Y(n_308)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_214),
.B2(n_215),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_240),
.B(n_250),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_225),
.B(n_239),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_224),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_238),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_238),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_234),
.B(n_237),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_237),
.A2(n_246),
.B(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_248),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_248),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_246),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_247),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_253),
.B(n_254),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_273),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_262),
.B2(n_263),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_262),
.C(n_273),
.Y(n_290)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVxp33_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_271),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_278),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_278),
.Y(n_295)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp33_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_290),
.B(n_291),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_296),
.B2(n_311),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_295),
.C(n_311),
.Y(n_314)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_304),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_297),
.B(n_305),
.C(n_306),
.Y(n_341)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_307),
.Y(n_335)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_314),
.B(n_315),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_344),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.Y(n_316)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_317),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_333),
.B2(n_334),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_319),
.B(n_333),
.Y(n_458)
);

OAI32xp33_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_323),
.A3(n_325),
.B1(n_326),
.B2(n_332),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx12f_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx5_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_341),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_341),
.B(n_342),
.C(n_344),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_346),
.B1(n_357),
.B2(n_369),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_345),
.B(n_358),
.C(n_363),
.Y(n_472)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_357),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_363),
.Y(n_357)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_359),
.Y(n_460)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx6_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx8_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_448),
.Y(n_371)
);

A2O1A1Ixp33_ASAP7_75t_SL g481 ( 
.A1(n_372),
.A2(n_448),
.B(n_482),
.C(n_485),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_424),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_373),
.B(n_424),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_400),
.C(n_409),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_374),
.B(n_400),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_388),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_389),
.C(n_397),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_384),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_376),
.B(n_384),
.Y(n_454)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_377),
.Y(n_414)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_385),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_397),
.Y(n_388)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_390),
.Y(n_423)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_394),
.Y(n_431)
);

INVx8_ASAP7_75t_L g421 ( 
.A(n_399),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_401),
.A2(n_402),
.B1(n_407),
.B2(n_408),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_402),
.B(n_407),
.Y(n_441)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_407),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_407),
.A2(n_408),
.B1(n_443),
.B2(n_444),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_407),
.A2(n_441),
.B(n_444),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_409),
.B(n_462),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_416),
.C(n_422),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_410),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_413),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_411),
.B(n_413),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_416),
.A2(n_417),
.B1(n_422),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_422),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_425),
.B(n_428),
.C(n_439),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_428),
.B1(n_439),
.B2(n_440),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_435),
.B(n_438),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_430),
.B(n_436),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_432),
.Y(n_498)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

FAx1_ASAP7_75t_SL g489 ( 
.A(n_438),
.B(n_490),
.CI(n_491),
.CON(n_489),
.SN(n_489)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_438),
.B(n_490),
.C(n_491),
.Y(n_511)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_447),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_446),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_461),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_449),
.B(n_461),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_454),
.C(n_455),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_450),
.A2(n_451),
.B1(n_454),
.B2(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_454),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_455),
.B(n_474),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_458),
.C(n_459),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_456),
.A2(n_457),
.B1(n_459),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_458),
.B(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_459),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_476),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_465),
.A2(n_483),
.B(n_484),
.Y(n_482)
);

NOR2x1_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_473),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_473),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_470),
.C(n_472),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_479),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_470),
.A2(n_471),
.B1(n_472),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_472),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_477),
.B(n_478),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_501),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_500),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_489),
.B(n_500),
.Y(n_513)
);

BUFx24_ASAP7_75t_SL g527 ( 
.A(n_489),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_493),
.B1(n_495),
.B2(n_499),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_492),
.A2(n_493),
.B1(n_507),
.B2(n_508),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_503),
.C(n_507),
.Y(n_519)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_495),
.Y(n_499)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_501),
.A2(n_513),
.B(n_514),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_511),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_502),
.B(n_511),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_504),
.B1(n_505),
.B2(n_506),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_519),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_516),
.B(n_519),
.Y(n_520)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

CKINVDCx14_ASAP7_75t_R g525 ( 
.A(n_526),
.Y(n_525)
);


endmodule