module real_jpeg_9468_n_18 (n_17, n_8, n_0, n_84, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_86, n_85, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_84;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_86;
input n_85;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_68;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_61;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_43;
wire n_57;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_0),
.A2(n_24),
.B(n_30),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_0),
.B(n_4),
.Y(n_30)
);

OAI221xp5_ASAP7_75t_L g32 ( 
.A1(n_0),
.A2(n_7),
.B1(n_33),
.B2(n_34),
.C(n_35),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_0),
.A2(n_5),
.B1(n_33),
.B2(n_36),
.Y(n_35)
);

NAND3xp33_ASAP7_75t_SL g44 ( 
.A(n_0),
.B(n_41),
.C(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_0),
.A2(n_27),
.B1(n_33),
.B2(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_1),
.B(n_84),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_3),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_2),
.B(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_6),
.A2(n_52),
.B1(n_55),
.B2(n_66),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_6),
.B(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_9),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_10),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_11),
.B(n_85),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_11),
.B(n_86),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_12),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_12),
.B(n_15),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_20),
.B1(n_21),
.B2(n_50),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_13),
.A2(n_50),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

AOI221xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_51),
.B1(n_67),
.B2(n_77),
.C(n_82),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_37),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_22),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_31),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_40),
.B(n_41),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_26),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_29),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_43),
.Y(n_42)
);

OAI221xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.C(n_47),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_41),
.A2(n_42),
.B(n_47),
.Y(n_76)
);

OAI221xp5_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_44),
.B1(n_71),
.B2(n_74),
.C(n_75),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_56),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_62),
.B(n_65),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B(n_61),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_64),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_73),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);


endmodule