module real_aes_14717_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_139;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
INVx2_ASAP7_75t_SL g261 ( .A(n_0), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_1), .Y(n_124) );
OA21x2_ASAP7_75t_L g110 ( .A1(n_2), .A2(n_39), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g163 ( .A(n_2), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_3), .B(n_93), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_4), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g562 ( .A(n_5), .Y(n_562) );
AND2x2_ASAP7_75t_L g165 ( .A(n_6), .B(n_135), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_7), .B(n_296), .Y(n_295) );
BUFx3_ASAP7_75t_L g531 ( .A(n_8), .Y(n_531) );
INVx1_ASAP7_75t_L g577 ( .A(n_9), .Y(n_577) );
INVx3_ASAP7_75t_L g608 ( .A(n_10), .Y(n_608) );
INVx1_ASAP7_75t_L g528 ( .A(n_11), .Y(n_528) );
INVx2_ASAP7_75t_L g537 ( .A(n_11), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_12), .B(n_130), .Y(n_201) );
INVx1_ASAP7_75t_L g95 ( .A(n_13), .Y(n_95) );
BUFx3_ASAP7_75t_L g117 ( .A(n_13), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_14), .B(n_134), .Y(n_212) );
AOI21xp33_ASAP7_75t_L g570 ( .A1(n_15), .A2(n_571), .B(n_574), .Y(n_570) );
INVxp33_ASAP7_75t_SL g627 ( .A(n_15), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_16), .A2(n_48), .B1(n_569), .B2(n_582), .Y(n_581) );
INVxp67_ASAP7_75t_L g644 ( .A(n_16), .Y(n_644) );
INVx1_ASAP7_75t_L g599 ( .A(n_17), .Y(n_599) );
INVx1_ASAP7_75t_L g604 ( .A(n_18), .Y(n_604) );
BUFx10_ASAP7_75t_L g711 ( .A(n_19), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_20), .A2(n_32), .B1(n_691), .B2(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_20), .Y(n_691) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_21), .Y(n_195) );
NAND3xp33_ASAP7_75t_L g277 ( .A(n_22), .B(n_115), .C(n_275), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_23), .B(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g620 ( .A(n_24), .B(n_621), .Y(n_620) );
INVxp33_ASAP7_75t_L g654 ( .A(n_24), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_24), .Y(n_657) );
AND2x2_ASAP7_75t_L g669 ( .A(n_24), .B(n_31), .Y(n_669) );
INVx1_ASAP7_75t_L g85 ( .A(n_25), .Y(n_85) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_26), .A2(n_52), .B1(n_524), .B2(n_532), .Y(n_523) );
INVx1_ASAP7_75t_L g661 ( .A(n_26), .Y(n_661) );
INVx2_ASAP7_75t_L g617 ( .A(n_27), .Y(n_617) );
AOI21xp33_ASAP7_75t_L g583 ( .A1(n_28), .A2(n_584), .B(n_586), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_28), .A2(n_74), .B1(n_646), .B2(n_648), .Y(n_645) );
OAI22xp33_ASAP7_75t_L g540 ( .A1(n_29), .A2(n_75), .B1(n_541), .B2(n_547), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_29), .A2(n_47), .B1(n_614), .B2(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_30), .B(n_255), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_30), .A2(n_730), .B1(n_736), .B2(n_738), .Y(n_729) );
INVx2_ASAP7_75t_L g621 ( .A(n_31), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_31), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_32), .B(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g692 ( .A(n_32), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g127 ( .A(n_33), .B(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g84 ( .A(n_34), .B(n_85), .Y(n_84) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_34), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_35), .B(n_134), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_36), .B(n_229), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_37), .B(n_134), .Y(n_291) );
INVx1_ASAP7_75t_L g527 ( .A(n_38), .Y(n_527) );
INVx1_ASAP7_75t_L g539 ( .A(n_38), .Y(n_539) );
INVx1_ASAP7_75t_L g162 ( .A(n_39), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_40), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_41), .A2(n_92), .B(n_259), .C(n_262), .Y(n_258) );
INVx1_ASAP7_75t_L g111 ( .A(n_42), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_43), .B(n_134), .Y(n_133) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_44), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_44), .Y(n_696) );
INVx3_ASAP7_75t_L g192 ( .A(n_45), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_46), .A2(n_74), .B1(n_568), .B2(n_569), .Y(n_567) );
INVxp67_ASAP7_75t_L g641 ( .A(n_46), .Y(n_641) );
INVxp67_ASAP7_75t_SL g553 ( .A(n_47), .Y(n_553) );
INVxp33_ASAP7_75t_SL g612 ( .A(n_48), .Y(n_612) );
BUFx3_ASAP7_75t_L g697 ( .A(n_49), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_50), .B(n_188), .Y(n_302) );
INVx1_ASAP7_75t_L g204 ( .A(n_51), .Y(n_204) );
INVx1_ASAP7_75t_L g678 ( .A(n_52), .Y(n_678) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_53), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_54), .B(n_119), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g114 ( .A(n_55), .B(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_56), .B(n_245), .Y(n_244) );
BUFx2_ASAP7_75t_L g688 ( .A(n_57), .Y(n_688) );
INVx1_ASAP7_75t_L g253 ( .A(n_58), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_59), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_60), .B(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_61), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g89 ( .A(n_62), .Y(n_89) );
BUFx3_ASAP7_75t_L g130 ( .A(n_62), .Y(n_130) );
INVx1_ASAP7_75t_L g158 ( .A(n_62), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_63), .B(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g190 ( .A(n_64), .Y(n_190) );
INVx2_ASAP7_75t_L g618 ( .A(n_65), .Y(n_618) );
INVxp67_ASAP7_75t_SL g630 ( .A(n_65), .Y(n_630) );
AND2x2_ASAP7_75t_L g634 ( .A(n_65), .B(n_617), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_66), .B(n_146), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_67), .B(n_135), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_68), .A2(n_521), .B1(n_700), .B2(n_719), .Y(n_718) );
CKINVDCx5p33_ASAP7_75t_R g719 ( .A(n_68), .Y(n_719) );
INVx2_ASAP7_75t_L g530 ( .A(n_69), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_70), .B(n_300), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_71), .Y(n_182) );
INVx1_ASAP7_75t_L g177 ( .A(n_72), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_73), .Y(n_149) );
OAI21xp33_ASAP7_75t_L g671 ( .A1(n_75), .A2(n_672), .B(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_76), .B(n_188), .Y(n_294) );
AOI21xp33_ASAP7_75t_SL g77 ( .A1(n_78), .A2(n_96), .B(n_519), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_86), .Y(n_80) );
AO31x2_ASAP7_75t_L g138 ( .A1(n_81), .A2(n_139), .A3(n_159), .B(n_165), .Y(n_138) );
AO31x2_ASAP7_75t_L g337 ( .A1(n_81), .A2(n_139), .A3(n_159), .B(n_165), .Y(n_337) );
BUFx2_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
OAI21xp33_ASAP7_75t_L g263 ( .A1(n_83), .A2(n_160), .B(n_257), .Y(n_263) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx2_ASAP7_75t_L g132 ( .A(n_84), .Y(n_132) );
INVx3_ASAP7_75t_L g180 ( .A(n_84), .Y(n_180) );
BUFx6f_ASAP7_75t_SL g211 ( .A(n_84), .Y(n_211) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_85), .Y(n_707) );
INVxp67_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AO21x2_ASAP7_75t_L g738 ( .A1(n_87), .A2(n_727), .B(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g87 ( .A(n_88), .B(n_90), .Y(n_87) );
AOI22x1_ASAP7_75t_L g140 ( .A1(n_88), .A2(n_141), .B1(n_150), .B2(n_155), .Y(n_140) );
INVx1_ASAP7_75t_L g262 ( .A(n_88), .Y(n_262) );
AOI21x1_ASAP7_75t_L g269 ( .A1(n_88), .A2(n_270), .B(n_271), .Y(n_269) );
BUFx3_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g122 ( .A(n_89), .Y(n_122) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
OAI22xp5_ASAP7_75t_L g150 ( .A1(n_92), .A2(n_151), .B1(n_153), .B2(n_154), .Y(n_150) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx2_ASAP7_75t_L g128 ( .A(n_94), .Y(n_128) );
INVx2_ASAP7_75t_L g297 ( .A(n_94), .Y(n_297) );
INVx1_ASAP7_75t_L g301 ( .A(n_94), .Y(n_301) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx2_ASAP7_75t_L g148 ( .A(n_95), .Y(n_148) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x4_ASAP7_75t_L g99 ( .A(n_100), .B(n_417), .Y(n_99) );
NOR3xp33_ASAP7_75t_L g100 ( .A(n_101), .B(n_339), .C(n_390), .Y(n_100) );
OAI221xp5_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_231), .B1(n_279), .B2(n_284), .C(n_308), .Y(n_101) );
AOI211xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_166), .B(n_213), .C(n_221), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g514 ( .A(n_104), .B(n_217), .Y(n_514) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_137), .Y(n_104) );
INVx1_ASAP7_75t_L g215 ( .A(n_105), .Y(n_215) );
AND2x2_ASAP7_75t_L g369 ( .A(n_105), .B(n_315), .Y(n_369) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_105), .Y(n_414) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g224 ( .A(n_106), .Y(n_224) );
INVx3_ASAP7_75t_L g317 ( .A(n_106), .Y(n_317) );
AND2x2_ASAP7_75t_L g345 ( .A(n_106), .B(n_226), .Y(n_345) );
AND2x2_ASAP7_75t_L g352 ( .A(n_106), .B(n_353), .Y(n_352) );
INVx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OAI21x1_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_112), .B(n_133), .Y(n_107) );
OAI21x1_ASAP7_75t_L g197 ( .A1(n_108), .A2(n_198), .B(n_212), .Y(n_197) );
BUFx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g136 ( .A(n_110), .Y(n_136) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_110), .Y(n_229) );
INVx1_ASAP7_75t_L g164 ( .A(n_111), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_123), .B(n_131), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B(n_121), .Y(n_113) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g206 ( .A(n_116), .Y(n_206) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_117), .Y(n_120) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_117), .Y(n_184) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g126 ( .A(n_120), .Y(n_126) );
INVx3_ASAP7_75t_L g143 ( .A(n_120), .Y(n_143) );
INVx2_ASAP7_75t_L g152 ( .A(n_120), .Y(n_152) );
INVx2_ASAP7_75t_L g238 ( .A(n_120), .Y(n_238) );
INVx3_ASAP7_75t_L g252 ( .A(n_120), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_121), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_121), .A2(n_243), .B(n_244), .Y(n_242) );
BUFx10_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g275 ( .A(n_122), .Y(n_275) );
O2A1O1Ixp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B(n_127), .C(n_129), .Y(n_123) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_130), .B(n_180), .Y(n_179) );
NOR3xp33_ASAP7_75t_L g189 ( .A(n_130), .B(n_180), .C(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g205 ( .A(n_130), .Y(n_205) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_131), .A2(n_269), .B(n_273), .Y(n_268) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_SL g306 ( .A(n_132), .Y(n_306) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_134), .Y(n_267) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OR2x2_ASAP7_75t_L g326 ( .A(n_138), .B(n_283), .Y(n_326) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_140), .A2(n_227), .B(n_230), .Y(n_226) );
OAI22x1_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_144), .B1(n_145), .B2(n_149), .Y(n_141) );
INVxp67_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g240 ( .A(n_147), .Y(n_240) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_147), .Y(n_255) );
INVx2_ASAP7_75t_L g272 ( .A(n_147), .Y(n_272) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_148), .Y(n_178) );
INVxp67_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVxp67_ASAP7_75t_L g200 ( .A(n_152), .Y(n_200) );
AOI21x1_ASAP7_75t_SL g250 ( .A1(n_155), .A2(n_251), .B(n_254), .Y(n_250) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_156), .A2(n_294), .B(n_295), .Y(n_293) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g186 ( .A(n_157), .Y(n_186) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx3_ASAP7_75t_L g241 ( .A(n_158), .Y(n_241) );
INVxp67_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AO21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_164), .Y(n_161) );
AOI21x1_ASAP7_75t_L g173 ( .A1(n_162), .A2(n_163), .B(n_164), .Y(n_173) );
INVx1_ASAP7_75t_L g230 ( .A(n_165), .Y(n_230) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI322xp5_ASAP7_75t_L g340 ( .A1(n_167), .A2(n_341), .A3(n_345), .B1(n_346), .B2(n_349), .C1(n_356), .C2(n_364), .Y(n_340) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g364 ( .A(n_169), .B(n_316), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_169), .B(n_316), .Y(n_379) );
AND2x2_ASAP7_75t_L g432 ( .A(n_169), .B(n_345), .Y(n_432) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_196), .Y(n_169) );
INVx3_ASAP7_75t_L g219 ( .A(n_170), .Y(n_219) );
AO21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_174), .B(n_194), .Y(n_170) );
AO21x1_ASAP7_75t_L g354 ( .A1(n_171), .A2(n_174), .B(n_194), .Y(n_354) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_SL g194 ( .A(n_172), .B(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_187), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_179), .B1(n_181), .B2(n_185), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
INVx1_ASAP7_75t_L g193 ( .A(n_178), .Y(n_193) );
INVx2_ASAP7_75t_L g245 ( .A(n_178), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_180), .B(n_186), .Y(n_185) );
NOR3xp33_ASAP7_75t_L g191 ( .A(n_180), .B(n_186), .C(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
INVx2_ASAP7_75t_L g188 ( .A(n_183), .Y(n_188) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g210 ( .A(n_184), .Y(n_210) );
INVx2_ASAP7_75t_L g260 ( .A(n_184), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B1(n_191), .B2(n_193), .Y(n_187) );
INVx1_ASAP7_75t_L g220 ( .A(n_196), .Y(n_220) );
AND2x2_ASAP7_75t_L g225 ( .A(n_196), .B(n_226), .Y(n_225) );
INVx3_ASAP7_75t_L g283 ( .A(n_196), .Y(n_283) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_196), .Y(n_374) );
INVx2_ASAP7_75t_L g387 ( .A(n_196), .Y(n_387) );
AND2x2_ASAP7_75t_L g397 ( .A(n_196), .B(n_219), .Y(n_397) );
INVx1_ASAP7_75t_L g458 ( .A(n_196), .Y(n_458) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OAI21x1_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_207), .B(n_211), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_202), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_206), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
OAI21x1_ASAP7_75t_L g235 ( .A1(n_211), .A2(n_236), .B(n_242), .Y(n_235) );
NOR2xp67_ASAP7_75t_L g213 ( .A(n_214), .B(n_216), .Y(n_213) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g475 ( .A(n_215), .Y(n_475) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
OR2x2_ASAP7_75t_L g501 ( .A(n_218), .B(n_336), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
INVx1_ASAP7_75t_L g315 ( .A(n_219), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_219), .B(n_317), .Y(n_338) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_223), .B(n_225), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_223), .B(n_423), .Y(n_447) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NOR2xp67_ASAP7_75t_L g281 ( .A(n_224), .B(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g406 ( .A(n_225), .B(n_407), .Y(n_406) );
AND2x4_ASAP7_75t_L g316 ( .A(n_226), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g425 ( .A(n_226), .Y(n_425) );
OAI21x1_ASAP7_75t_L g234 ( .A1(n_227), .A2(n_235), .B(n_246), .Y(n_234) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_227), .A2(n_235), .B(n_246), .Y(n_287) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NOR2x1_ASAP7_75t_SL g304 ( .A(n_228), .B(n_305), .Y(n_304) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g324 ( .A(n_229), .Y(n_324) );
OR2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_247), .Y(n_231) );
AND2x2_ASAP7_75t_L g331 ( .A(n_232), .B(n_289), .Y(n_331) );
OR2x2_ASAP7_75t_L g498 ( .A(n_232), .B(n_329), .Y(n_498) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g311 ( .A(n_233), .B(n_312), .Y(n_311) );
BUFx3_ASAP7_75t_L g343 ( .A(n_233), .Y(n_343) );
AND2x2_ASAP7_75t_L g470 ( .A(n_233), .B(n_248), .Y(n_470) );
AND2x4_ASAP7_75t_L g486 ( .A(n_233), .B(n_383), .Y(n_486) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_234), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_239), .B(n_241), .Y(n_236) );
INVx2_ASAP7_75t_L g303 ( .A(n_241), .Y(n_303) );
INVxp67_ASAP7_75t_L g276 ( .A(n_245), .Y(n_276) );
OR2x2_ASAP7_75t_L g347 ( .A(n_247), .B(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g394 ( .A(n_247), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_264), .Y(n_247) );
AND2x4_ASAP7_75t_L g286 ( .A(n_248), .B(n_287), .Y(n_286) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_248), .Y(n_333) );
INVx1_ASAP7_75t_L g359 ( .A(n_248), .Y(n_359) );
AND2x2_ASAP7_75t_L g402 ( .A(n_248), .B(n_322), .Y(n_402) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g321 ( .A(n_249), .Y(n_321) );
OAI21x1_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_256), .B(n_263), .Y(n_249) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_261), .A2(n_521), .B1(n_700), .B2(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_261), .Y(n_737) );
AND2x4_ASAP7_75t_L g363 ( .A(n_264), .B(n_289), .Y(n_363) );
INVx1_ASAP7_75t_L g377 ( .A(n_264), .Y(n_377) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVxp67_ASAP7_75t_SL g307 ( .A(n_265), .Y(n_307) );
INVx2_ASAP7_75t_L g330 ( .A(n_265), .Y(n_330) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OAI21x1_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_268), .B(n_278), .Y(n_266) );
OA21x2_ASAP7_75t_L g322 ( .A1(n_268), .A2(n_278), .B(n_323), .Y(n_322) );
OAI21xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_276), .B(n_277), .Y(n_273) );
INVxp67_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g444 ( .A(n_282), .B(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g465 ( .A(n_282), .Y(n_465) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_283), .B(n_454), .Y(n_468) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g375 ( .A(n_286), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g438 ( .A(n_286), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g463 ( .A(n_286), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g507 ( .A(n_286), .Y(n_507) );
AND2x2_ASAP7_75t_L g360 ( .A(n_287), .B(n_330), .Y(n_360) );
AND2x4_ASAP7_75t_L g362 ( .A(n_287), .B(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g367 ( .A(n_287), .B(n_320), .Y(n_367) );
AND2x4_ASAP7_75t_L g382 ( .A(n_287), .B(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_307), .Y(n_288) );
INVx2_ASAP7_75t_L g312 ( .A(n_289), .Y(n_312) );
INVx2_ASAP7_75t_L g334 ( .A(n_289), .Y(n_334) );
BUFx2_ASAP7_75t_L g348 ( .A(n_289), .Y(n_348) );
INVx1_ASAP7_75t_L g404 ( .A(n_289), .Y(n_404) );
AND2x2_ASAP7_75t_L g464 ( .A(n_289), .B(n_322), .Y(n_464) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2x1_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
OAI21x1_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_298), .B(n_304), .Y(n_292) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_302), .B(n_303), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g344 ( .A(n_307), .B(n_312), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_318), .B(n_325), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_311), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g487 ( .A(n_311), .Y(n_487) );
AND2x2_ASAP7_75t_L g499 ( .A(n_311), .B(n_319), .Y(n_499) );
BUFx2_ASAP7_75t_L g439 ( .A(n_312), .Y(n_439) );
INVx1_ASAP7_75t_L g513 ( .A(n_312), .Y(n_513) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_316), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g388 ( .A(n_316), .Y(n_388) );
INVx2_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_319), .A2(n_510), .B1(n_512), .B2(n_514), .Y(n_509) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_SL g320 ( .A(n_321), .B(n_322), .Y(n_320) );
OR2x6_ASAP7_75t_L g329 ( .A(n_321), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g383 ( .A(n_321), .Y(n_383) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B1(n_332), .B2(n_335), .Y(n_325) );
INVx2_ASAP7_75t_SL g370 ( .A(n_326), .Y(n_370) );
OR2x2_ASAP7_75t_L g399 ( .A(n_326), .B(n_338), .Y(n_399) );
INVx2_ASAP7_75t_L g436 ( .A(n_327), .Y(n_436) );
NAND2x1p5_ASAP7_75t_L g327 ( .A(n_328), .B(n_331), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g484 ( .A(n_329), .B(n_334), .Y(n_484) );
OR2x2_ASAP7_75t_L g517 ( .A(n_329), .B(n_343), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AND2x2_ASAP7_75t_L g405 ( .A(n_333), .B(n_360), .Y(n_405) );
INVx1_ASAP7_75t_L g381 ( .A(n_334), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_334), .B(n_358), .Y(n_421) );
OR2x2_ASAP7_75t_L g457 ( .A(n_334), .B(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx1_ASAP7_75t_L g454 ( .A(n_336), .Y(n_454) );
BUFx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g355 ( .A(n_337), .Y(n_355) );
INVx1_ASAP7_75t_L g407 ( .A(n_338), .Y(n_407) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_338), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_365), .Y(n_339) );
INVx2_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx2_ASAP7_75t_L g411 ( .A(n_343), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_343), .B(n_363), .Y(n_416) );
AND2x2_ASAP7_75t_L g429 ( .A(n_344), .B(n_430), .Y(n_429) );
BUFx3_ASAP7_75t_L g489 ( .A(n_344), .Y(n_489) );
INVx1_ASAP7_75t_L g491 ( .A(n_345), .Y(n_491) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g469 ( .A(n_348), .B(n_470), .Y(n_469) );
NAND2x1_ASAP7_75t_L g455 ( .A(n_349), .B(n_456), .Y(n_455) );
INVx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g482 ( .A(n_350), .Y(n_482) );
OR2x6_ASAP7_75t_L g350 ( .A(n_351), .B(n_355), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g445 ( .A(n_352), .Y(n_445) );
AND2x2_ASAP7_75t_L g505 ( .A(n_352), .B(n_355), .Y(n_505) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g386 ( .A(n_354), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_354), .B(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_355), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g496 ( .A(n_355), .Y(n_496) );
NAND2x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_361), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_358), .Y(n_459) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AOI221x1_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_368), .B1(n_371), .B2(n_375), .C(n_378), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_368), .A2(n_401), .B1(n_405), .B2(n_406), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_368), .A2(n_409), .B1(n_412), .B2(n_415), .Y(n_408) );
INVxp67_ASAP7_75t_SL g506 ( .A(n_368), .Y(n_506) );
AND2x4_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g446 ( .A(n_373), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVxp67_ASAP7_75t_SL g389 ( .A(n_376), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_376), .B(n_411), .Y(n_410) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_384), .B2(n_389), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
AND2x4_ASAP7_75t_L g449 ( .A(n_381), .B(n_394), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_382), .A2(n_392), .B1(n_395), .B2(n_398), .Y(n_391) );
AND2x2_ASAP7_75t_L g472 ( .A(n_382), .B(n_439), .Y(n_472) );
OR2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_388), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g453 ( .A(n_386), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g474 ( .A(n_386), .Y(n_474) );
AND2x2_ASAP7_75t_L g495 ( .A(n_386), .B(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g512 ( .A(n_386), .B(n_513), .Y(n_512) );
NAND3xp33_ASAP7_75t_SL g390 ( .A(n_391), .B(n_400), .C(n_408), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_397), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g443 ( .A(n_405), .Y(n_443) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_406), .A2(n_467), .B(n_469), .Y(n_466) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVxp67_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g511 ( .A(n_414), .Y(n_511) );
INVx1_ASAP7_75t_L g427 ( .A(n_415), .Y(n_427) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NOR2x1_ASAP7_75t_L g417 ( .A(n_418), .B(n_476), .Y(n_417) );
NAND3xp33_ASAP7_75t_SL g418 ( .A(n_419), .B(n_433), .C(n_450), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_422), .B(n_426), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B(n_431), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI22xp5_ASAP7_75t_SL g510 ( .A1(n_430), .A2(n_485), .B1(n_496), .B2(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g518 ( .A(n_430), .Y(n_518) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_440), .B(n_442), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
INVx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_446), .B2(n_448), .Y(n_442) );
INVx1_ASAP7_75t_L g462 ( .A(n_445), .Y(n_462) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_449), .A2(n_473), .B(n_493), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_459), .B(n_460), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_455), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_456), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g481 ( .A(n_458), .Y(n_481) );
NAND3xp33_ASAP7_75t_SL g460 ( .A(n_461), .B(n_466), .C(n_471), .Y(n_460) );
NAND3xp33_ASAP7_75t_SL g461 ( .A(n_462), .B(n_463), .C(n_465), .Y(n_461) );
AND2x2_ASAP7_75t_L g493 ( .A(n_464), .B(n_486), .Y(n_493) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .C(n_475), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_502), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_483), .B(n_490), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2x1p5_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND4xp25_ASAP7_75t_SL g483 ( .A(n_484), .B(n_485), .C(n_487), .D(n_488), .Y(n_483) );
INVx3_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OAI21xp5_ASAP7_75t_SL g490 ( .A1(n_491), .A2(n_492), .B(n_494), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_497), .B1(n_499), .B2(n_500), .Y(n_494) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_503), .B(n_508), .Y(n_502) );
AOI21xp5_ASAP7_75t_SL g503 ( .A1(n_504), .A2(n_506), .B(n_507), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_505), .A2(n_514), .B1(n_516), .B2(n_518), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_509), .B(n_515), .Y(n_508) );
INVx2_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
OAI221xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_701), .B1(n_718), .B2(n_720), .C(n_729), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_685), .B1(n_686), .B2(n_700), .Y(n_520) );
INVx1_ASAP7_75t_L g700 ( .A(n_521), .Y(n_700) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_609), .Y(n_521) );
OAI31xp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_540), .A3(n_551), .B(n_605), .Y(n_522) );
OR2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_529), .Y(n_524) );
INVx8_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
AND2x4_ASAP7_75t_L g550 ( .A(n_527), .B(n_536), .Y(n_550) );
INVx1_ASAP7_75t_L g596 ( .A(n_528), .Y(n_596) );
OR2x6_ASAP7_75t_SL g533 ( .A(n_529), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g543 ( .A(n_529), .Y(n_543) );
OR2x6_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g560 ( .A(n_530), .Y(n_560) );
BUFx2_ASAP7_75t_L g588 ( .A(n_530), .Y(n_588) );
AND2x2_ASAP7_75t_L g559 ( .A(n_531), .B(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g575 ( .A(n_531), .B(n_560), .Y(n_575) );
AND2x4_ASAP7_75t_L g587 ( .A(n_531), .B(n_588), .Y(n_587) );
BUFx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_535), .Y(n_566) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_535), .Y(n_580) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g546 ( .A(n_537), .B(n_538), .Y(n_546) );
AND2x2_ASAP7_75t_L g557 ( .A(n_537), .B(n_539), .Y(n_557) );
INVx1_ASAP7_75t_L g602 ( .A(n_538), .Y(n_602) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
NAND2x1_ASAP7_75t_L g547 ( .A(n_543), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx5_ASAP7_75t_L g569 ( .A(n_545), .Y(n_569) );
INVx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx4_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_550), .Y(n_573) );
NAND5xp2_ASAP7_75t_L g551 ( .A(n_552), .B(n_561), .C(n_576), .D(n_589), .E(n_592), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
AND2x4_ASAP7_75t_L g554 ( .A(n_555), .B(n_558), .Y(n_554) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_555), .Y(n_568) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_557), .Y(n_585) );
INVx3_ASAP7_75t_L g590 ( .A(n_558), .Y(n_590) );
BUFx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g598 ( .A(n_559), .Y(n_598) );
OAI211xp5_ASAP7_75t_SL g561 ( .A1(n_562), .A2(n_563), .B(n_567), .C(n_570), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_562), .A2(n_627), .B1(n_628), .B2(n_632), .Y(n_626) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx5_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g591 ( .A(n_566), .Y(n_591) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
BUFx2_ASAP7_75t_L g582 ( .A(n_573), .Y(n_582) );
BUFx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx6f_ASAP7_75t_L g712 ( .A(n_575), .Y(n_712) );
OAI211xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B(n_581), .C(n_583), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_577), .A2(n_612), .B1(n_613), .B2(n_622), .Y(n_611) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
BUFx4f_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x6_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_599), .B1(n_600), .B2(n_604), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_SL g717 ( .A(n_595), .Y(n_717) );
AND2x4_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_596), .B(n_710), .C(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g603 ( .A(n_598), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_599), .A2(n_674), .B1(n_678), .B2(n_679), .Y(n_673) );
AND2x4_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVx3_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI221xp5_ASAP7_75t_SL g658 ( .A1(n_604), .A2(n_659), .B1(n_661), .B2(n_662), .C(n_663), .Y(n_658) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x6_ASAP7_75t_L g655 ( .A(n_607), .B(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x4_ASAP7_75t_L g619 ( .A(n_608), .B(n_620), .Y(n_619) );
AND3x2_ASAP7_75t_SL g651 ( .A(n_608), .B(n_652), .C(n_654), .Y(n_651) );
NAND2x1p5_ASAP7_75t_L g668 ( .A(n_608), .B(n_669), .Y(n_668) );
AND2x4_ASAP7_75t_SL g684 ( .A(n_608), .B(n_669), .Y(n_684) );
NOR3xp33_ASAP7_75t_SL g609 ( .A(n_610), .B(n_635), .C(n_671), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_626), .Y(n_610) );
AND2x4_ASAP7_75t_L g613 ( .A(n_614), .B(n_619), .Y(n_613) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_615), .Y(n_649) );
AND2x4_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx1_ASAP7_75t_L g631 ( .A(n_616), .Y(n_631) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_616), .Y(n_677) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g624 ( .A(n_617), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_617), .B(n_618), .Y(n_640) );
INVx2_ASAP7_75t_L g625 ( .A(n_618), .Y(n_625) );
AND2x2_ASAP7_75t_L g622 ( .A(n_619), .B(n_623), .Y(n_622) );
AND2x6_ASAP7_75t_L g628 ( .A(n_619), .B(n_629), .Y(n_628) );
AND2x4_ASAP7_75t_L g632 ( .A(n_619), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g653 ( .A(n_621), .Y(n_653) );
AND2x4_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g643 ( .A(n_624), .B(n_625), .Y(n_643) );
AND2x4_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g683 ( .A(n_630), .Y(n_683) );
INVx3_ASAP7_75t_L g647 ( .A(n_633), .Y(n_647) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx4f_ASAP7_75t_L g665 ( .A(n_634), .Y(n_665) );
OAI221xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_650), .B1(n_655), .B2(n_658), .C(n_666), .Y(n_635) );
OAI221xp5_ASAP7_75t_SL g636 ( .A1(n_637), .A2(n_641), .B1(n_642), .B2(n_644), .C(n_645), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g660 ( .A(n_639), .Y(n_660) );
OR2x4_ASAP7_75t_L g672 ( .A(n_639), .B(n_668), .Y(n_672) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
BUFx3_ASAP7_75t_L g662 ( .A(n_642), .Y(n_662) );
BUFx12f_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_643), .Y(n_670) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
BUFx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
BUFx3_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OR2x6_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
OR2x6_ASAP7_75t_L g675 ( .A(n_668), .B(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
BUFx4f_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AND2x4_ASAP7_75t_L g680 ( .A(n_681), .B(n_684), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_694), .B1(n_695), .B2(n_699), .Y(n_686) );
CKINVDCx5p33_ASAP7_75t_R g699 ( .A(n_687), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B1(n_690), .B2(n_693), .Y(n_687) );
INVx1_ASAP7_75t_SL g693 ( .A(n_688), .Y(n_693) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
CKINVDCx5p33_ASAP7_75t_R g698 ( .A(n_697), .Y(n_698) );
INVx3_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x6_ASAP7_75t_L g702 ( .A(n_703), .B(n_713), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_708), .Y(n_703) );
INVxp67_ASAP7_75t_L g734 ( .A(n_704), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g728 ( .A(n_705), .Y(n_728) );
INVx1_ASAP7_75t_L g740 ( .A(n_706), .Y(n_740) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
BUFx2_ASAP7_75t_L g727 ( .A(n_707), .Y(n_727) );
INVxp67_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_709), .B(n_717), .Y(n_735) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
CKINVDCx11_ASAP7_75t_R g715 ( .A(n_711), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .Y(n_713) );
CKINVDCx5p33_ASAP7_75t_R g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_721), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_722), .Y(n_721) );
INVx3_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_724), .Y(n_723) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g739 ( .A(n_728), .B(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
BUFx4f_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx4_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
endmodule