module fake_netlist_6_2342_n_1516 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_350, n_78, n_84, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1516);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1516;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_1413;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1504;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_1437;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_1485;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_1408;
wire n_1196;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_1028;
wire n_576;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1109;
wire n_712;
wire n_1276;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_859;
wire n_570;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_629;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

INVx1_ASAP7_75t_L g392 ( 
.A(n_61),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_236),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_323),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_379),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_256),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_81),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_167),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_357),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_77),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_382),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_341),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_47),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_13),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_122),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_87),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_23),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_186),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_252),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_29),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_60),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_306),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_54),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_266),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_28),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_171),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_109),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_170),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_374),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_367),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_218),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_372),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_51),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_50),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_349),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_230),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_100),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_177),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_146),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_376),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_378),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_14),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_36),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_365),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_83),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_106),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_384),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_35),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_327),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_169),
.Y(n_440)
);

BUFx5_ASAP7_75t_L g441 ( 
.A(n_324),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_30),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_40),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_112),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_155),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_42),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_55),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_14),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_287),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_41),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_334),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_316),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_114),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_339),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_320),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_352),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_91),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_102),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_273),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_117),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_11),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_107),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_380),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_261),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_131),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_34),
.Y(n_466)
);

BUFx10_ASAP7_75t_L g467 ( 
.A(n_233),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_326),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_149),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_333),
.Y(n_470)
);

BUFx10_ASAP7_75t_L g471 ( 
.A(n_31),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_97),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_257),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_68),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_258),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_370),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_160),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_383),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_191),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_205),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_299),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_98),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_189),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_45),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_262),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_309),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_342),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_172),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_204),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_202),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_165),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_7),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_78),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_371),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_190),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_329),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_156),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_119),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_274),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_222),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_168),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_8),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_187),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_161),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_152),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_179),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_260),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_174),
.Y(n_508)
);

BUFx10_ASAP7_75t_L g509 ( 
.A(n_16),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_34),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_246),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_20),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_360),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_344),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_35),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_29),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_79),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_243),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_377),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_4),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_270),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_354),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_249),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_196),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_181),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_234),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_113),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_121),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_366),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_303),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_36),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_137),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_239),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_294),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_198),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_185),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_126),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_381),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_238),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_123),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_118),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_364),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_105),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_1),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_340),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_59),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_69),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_373),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_206),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_289),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_368),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_244),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_242),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_17),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_312),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_145),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_86),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_45),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_103),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_53),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_237),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_162),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_369),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_330),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_42),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_183),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_166),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_180),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_245),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_297),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_296),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_52),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_355),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_325),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_38),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_16),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_322),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_31),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_277),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_197),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_84),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_375),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_175),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_193),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_184),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_321),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_32),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_73),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_151),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_247),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_127),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_426),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_554),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_554),
.Y(n_594)
);

CKINVDCx14_ASAP7_75t_R g595 ( 
.A(n_400),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_R g596 ( 
.A(n_430),
.B(n_0),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_441),
.Y(n_597)
);

INVxp33_ASAP7_75t_SL g598 ( 
.A(n_459),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_435),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_404),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_459),
.B(n_0),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_464),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_398),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_401),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_443),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_402),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_481),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_578),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_587),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_408),
.Y(n_610)
);

CKINVDCx16_ASAP7_75t_R g611 ( 
.A(n_454),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_397),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_556),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_411),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_556),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_392),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_393),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_394),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_395),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_412),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_396),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_413),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_414),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_483),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_416),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_417),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_405),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_409),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_534),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_419),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_423),
.Y(n_631)
);

INVxp67_ASAP7_75t_SL g632 ( 
.A(n_581),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_422),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_428),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_441),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_541),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_437),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_586),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_420),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_453),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_446),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_407),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_455),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_471),
.Y(n_644)
);

INVxp67_ASAP7_75t_SL g645 ( 
.A(n_420),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_424),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_425),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_456),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_457),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_458),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_427),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_460),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g653 ( 
.A(n_399),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_474),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_410),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_429),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_431),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_434),
.Y(n_658)
);

NOR2xp67_ASAP7_75t_L g659 ( 
.A(n_512),
.B(n_1),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_501),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_403),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_504),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_469),
.B(n_2),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_506),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_439),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_445),
.B(n_2),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_440),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_471),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_444),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_517),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_452),
.B(n_3),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_524),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_529),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_495),
.B(n_3),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_447),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_449),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_406),
.B(n_4),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_451),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_462),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_463),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_472),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_473),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_475),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_415),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_530),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_533),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_535),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_539),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_477),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_441),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_542),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_478),
.Y(n_692)
);

INVxp67_ASAP7_75t_SL g693 ( 
.A(n_485),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_479),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_480),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_612),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_612),
.Y(n_697)
);

OA21x2_ASAP7_75t_L g698 ( 
.A1(n_677),
.A2(n_549),
.B(n_548),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_616),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_617),
.Y(n_700)
);

NOR3xp33_ASAP7_75t_L g701 ( 
.A(n_601),
.B(n_433),
.C(n_432),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_612),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_612),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_655),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_600),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_598),
.B(n_467),
.Y(n_706)
);

OA21x2_ASAP7_75t_L g707 ( 
.A1(n_671),
.A2(n_552),
.B(n_551),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_605),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_618),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_684),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_608),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_619),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_609),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_684),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_621),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_597),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_641),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_655),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_627),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_628),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_674),
.B(n_639),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_635),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_690),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_630),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_633),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_634),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_645),
.B(n_482),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_593),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_637),
.B(n_640),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_594),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_643),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_648),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_649),
.B(n_591),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_603),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_604),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_650),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_652),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_654),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_660),
.B(n_487),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_662),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_661),
.B(n_438),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_664),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_642),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_647),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_670),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_672),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_673),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_685),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_686),
.Y(n_749)
);

INVx1_ASAP7_75t_SL g750 ( 
.A(n_596),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_687),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_688),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_691),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_642),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_653),
.B(n_693),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_613),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_615),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_666),
.B(n_467),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_663),
.B(n_632),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_606),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_663),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_659),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_666),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_610),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_614),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_620),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_622),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_623),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_625),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_626),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_611),
.B(n_470),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_631),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_646),
.B(n_590),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_651),
.B(n_470),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_656),
.Y(n_775)
);

NAND2xp33_ASAP7_75t_L g776 ( 
.A(n_665),
.B(n_442),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_669),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_675),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_676),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_679),
.A2(n_421),
.B(n_418),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_681),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_595),
.B(n_476),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_716),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_750),
.B(n_595),
.Y(n_784)
);

INVx8_ASAP7_75t_L g785 ( 
.A(n_735),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_773),
.B(n_683),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_773),
.B(n_689),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_750),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_722),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_696),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_728),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_721),
.A2(n_694),
.B(n_692),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_770),
.B(n_657),
.Y(n_793)
);

INVx4_ASAP7_75t_L g794 ( 
.A(n_770),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_697),
.Y(n_795)
);

INVx8_ASAP7_75t_L g796 ( 
.A(n_770),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_721),
.B(n_489),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_717),
.B(n_644),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_755),
.B(n_500),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_699),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_696),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_697),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_697),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_700),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_709),
.Y(n_805)
);

INVx4_ASAP7_75t_L g806 ( 
.A(n_778),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_702),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_L g808 ( 
.A(n_759),
.B(n_397),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_761),
.A2(n_436),
.B1(n_465),
.B2(n_397),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_703),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_712),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_755),
.B(n_559),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_723),
.Y(n_813)
);

OAI21xp33_ASAP7_75t_L g814 ( 
.A1(n_763),
.A2(n_450),
.B(n_448),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_715),
.Y(n_815)
);

INVx5_ASAP7_75t_L g816 ( 
.A(n_705),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_727),
.B(n_488),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_719),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_720),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_734),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_726),
.Y(n_821)
);

NOR2x1p5_ASAP7_75t_L g822 ( 
.A(n_782),
.B(n_461),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_714),
.B(n_743),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_731),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_737),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_738),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_778),
.Y(n_827)
);

NAND2x1p5_ASAP7_75t_L g828 ( 
.A(n_778),
.B(n_397),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_744),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_745),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_727),
.B(n_658),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_764),
.B(n_667),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_728),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_728),
.Y(n_834)
);

BUFx4f_ASAP7_75t_L g835 ( 
.A(n_730),
.Y(n_835)
);

INVx4_ASAP7_75t_L g836 ( 
.A(n_730),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_730),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_746),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_740),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_740),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_749),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_780),
.A2(n_680),
.B(n_678),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_760),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_766),
.B(n_682),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_740),
.Y(n_845)
);

OR2x6_ASAP7_75t_L g846 ( 
.A(n_771),
.B(n_668),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_714),
.B(n_695),
.Y(n_847)
);

INVx8_ASAP7_75t_L g848 ( 
.A(n_705),
.Y(n_848)
);

NAND2x1p5_ASAP7_75t_L g849 ( 
.A(n_760),
.B(n_436),
.Y(n_849)
);

OAI22xp33_ASAP7_75t_L g850 ( 
.A1(n_759),
.A2(n_484),
.B1(n_492),
.B2(n_466),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_758),
.B(n_706),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_742),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_751),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_753),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_743),
.B(n_596),
.Y(n_855)
);

AND2x6_ASAP7_75t_L g856 ( 
.A(n_765),
.B(n_436),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_762),
.B(n_710),
.Y(n_857)
);

INVx4_ASAP7_75t_L g858 ( 
.A(n_742),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_724),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_757),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_742),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_768),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_747),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_747),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_733),
.B(n_490),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_747),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_710),
.B(n_754),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_725),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_767),
.B(n_592),
.Y(n_869)
);

OAI22xp33_ASAP7_75t_SL g870 ( 
.A1(n_758),
.A2(n_706),
.B1(n_774),
.B2(n_771),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_774),
.B(n_476),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_752),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_769),
.B(n_562),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_775),
.B(n_563),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_772),
.B(n_599),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_748),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_786),
.B(n_777),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_851),
.A2(n_779),
.B1(n_781),
.B2(n_701),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_830),
.Y(n_879)
);

AO22x2_ASAP7_75t_L g880 ( 
.A1(n_871),
.A2(n_823),
.B1(n_870),
.B2(n_847),
.Y(n_880)
);

AO22x2_ASAP7_75t_L g881 ( 
.A1(n_857),
.A2(n_741),
.B1(n_701),
.B2(n_580),
.Y(n_881)
);

AO22x2_ASAP7_75t_L g882 ( 
.A1(n_867),
.A2(n_585),
.B1(n_589),
.B2(n_566),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_830),
.Y(n_883)
);

AO22x2_ASAP7_75t_L g884 ( 
.A1(n_793),
.A2(n_486),
.B1(n_527),
.B2(n_468),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_792),
.B(n_733),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_838),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_838),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_800),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_840),
.Y(n_889)
);

CKINVDCx16_ASAP7_75t_R g890 ( 
.A(n_829),
.Y(n_890)
);

BUFx8_ASAP7_75t_L g891 ( 
.A(n_798),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_797),
.A2(n_707),
.B1(n_698),
.B2(n_540),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_813),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_788),
.B(n_717),
.Y(n_894)
);

AND2x6_ASAP7_75t_L g895 ( 
.A(n_784),
.B(n_436),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_804),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_855),
.B(n_756),
.Y(n_897)
);

AO22x2_ASAP7_75t_L g898 ( 
.A1(n_842),
.A2(n_536),
.B1(n_553),
.B2(n_739),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_805),
.Y(n_899)
);

OR2x6_ASAP7_75t_L g900 ( 
.A(n_796),
.B(n_729),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_785),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_787),
.B(n_739),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_811),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_815),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_827),
.B(n_756),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_859),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_799),
.A2(n_607),
.B1(n_624),
.B2(n_602),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_843),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_850),
.A2(n_707),
.B1(n_698),
.B2(n_441),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_796),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_818),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_819),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_817),
.B(n_776),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_821),
.Y(n_914)
);

INVx6_ASAP7_75t_L g915 ( 
.A(n_794),
.Y(n_915)
);

AO22x2_ASAP7_75t_L g916 ( 
.A1(n_812),
.A2(n_509),
.B1(n_7),
.B2(n_5),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_824),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_825),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_831),
.A2(n_636),
.B1(n_638),
.B2(n_629),
.Y(n_919)
);

AO22x2_ASAP7_75t_L g920 ( 
.A1(n_812),
.A2(n_509),
.B1(n_8),
.B2(n_5),
.Y(n_920)
);

NAND2x1p5_ASAP7_75t_L g921 ( 
.A(n_794),
.B(n_806),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_868),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_865),
.B(n_732),
.Y(n_923)
);

AO22x2_ASAP7_75t_L g924 ( 
.A1(n_873),
.A2(n_10),
.B1(n_6),
.B2(n_9),
.Y(n_924)
);

NAND2x1p5_ASAP7_75t_L g925 ( 
.A(n_806),
.B(n_704),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_873),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_826),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_841),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_783),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_853),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_854),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_840),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_872),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_783),
.B(n_732),
.Y(n_934)
);

AO22x2_ASAP7_75t_L g935 ( 
.A1(n_874),
.A2(n_10),
.B1(n_6),
.B2(n_9),
.Y(n_935)
);

NOR2xp67_ASAP7_75t_L g936 ( 
.A(n_832),
.B(n_736),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_785),
.B(n_729),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_862),
.B(n_748),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_872),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_860),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_789),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_820),
.B(n_704),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_874),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_789),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_846),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_844),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_807),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_810),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_790),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_801),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_861),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_SL g952 ( 
.A1(n_846),
.A2(n_875),
.B1(n_869),
.B2(n_510),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_864),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_828),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_822),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_866),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_834),
.Y(n_957)
);

NAND2x1p5_ASAP7_75t_L g958 ( 
.A(n_858),
.B(n_718),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_839),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_845),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_863),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_852),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_852),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_876),
.Y(n_964)
);

OAI21xp33_ASAP7_75t_L g965 ( 
.A1(n_814),
.A2(n_515),
.B(n_502),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_834),
.Y(n_966)
);

AO22x2_ASAP7_75t_L g967 ( 
.A1(n_808),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_967)
);

AO22x2_ASAP7_75t_L g968 ( 
.A1(n_858),
.A2(n_17),
.B1(n_12),
.B2(n_15),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_876),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_791),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_833),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_837),
.B(n_708),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_837),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_848),
.Y(n_974)
);

AO22x2_ASAP7_75t_L g975 ( 
.A1(n_836),
.A2(n_19),
.B1(n_15),
.B2(n_18),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_835),
.B(n_748),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_877),
.B(n_902),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_936),
.B(n_849),
.Y(n_978)
);

NAND2xp33_ASAP7_75t_SL g979 ( 
.A(n_908),
.B(n_491),
.Y(n_979)
);

NAND2xp33_ASAP7_75t_SL g980 ( 
.A(n_910),
.B(n_493),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_897),
.B(n_885),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_878),
.B(n_836),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_946),
.B(n_816),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_938),
.B(n_816),
.Y(n_984)
);

NAND2xp33_ASAP7_75t_SL g985 ( 
.A(n_955),
.B(n_494),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_894),
.B(n_816),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_942),
.B(n_718),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_943),
.B(n_848),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_913),
.B(n_736),
.Y(n_989)
);

NAND2xp33_ASAP7_75t_SL g990 ( 
.A(n_952),
.B(n_496),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_921),
.B(n_795),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_905),
.B(n_795),
.Y(n_992)
);

NAND2xp33_ASAP7_75t_SL g993 ( 
.A(n_926),
.B(n_945),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_923),
.B(n_809),
.Y(n_994)
);

NAND2xp33_ASAP7_75t_SL g995 ( 
.A(n_954),
.B(n_497),
.Y(n_995)
);

NAND2xp33_ASAP7_75t_SL g996 ( 
.A(n_901),
.B(n_498),
.Y(n_996)
);

NAND2xp33_ASAP7_75t_SL g997 ( 
.A(n_976),
.B(n_499),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_879),
.B(n_802),
.Y(n_998)
);

NAND2xp33_ASAP7_75t_SL g999 ( 
.A(n_883),
.B(n_503),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_886),
.B(n_802),
.Y(n_1000)
);

NAND2xp33_ASAP7_75t_SL g1001 ( 
.A(n_887),
.B(n_962),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_888),
.B(n_803),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_896),
.B(n_803),
.Y(n_1003)
);

NAND2xp33_ASAP7_75t_SL g1004 ( 
.A(n_963),
.B(n_505),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_899),
.B(n_705),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_903),
.B(n_904),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_911),
.B(n_856),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_912),
.B(n_856),
.Y(n_1008)
);

NAND2xp33_ASAP7_75t_SL g1009 ( 
.A(n_964),
.B(n_507),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_914),
.B(n_713),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_917),
.B(n_713),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_918),
.B(n_711),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_927),
.B(n_713),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_928),
.B(n_508),
.Y(n_1014)
);

NAND2xp33_ASAP7_75t_SL g1015 ( 
.A(n_957),
.B(n_511),
.Y(n_1015)
);

NAND2xp33_ASAP7_75t_SL g1016 ( 
.A(n_966),
.B(n_513),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_930),
.B(n_514),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_931),
.B(n_518),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_940),
.B(n_519),
.Y(n_1019)
);

NAND2xp33_ASAP7_75t_SL g1020 ( 
.A(n_907),
.B(n_521),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_929),
.B(n_522),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_937),
.B(n_516),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_944),
.B(n_523),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_941),
.B(n_856),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_933),
.B(n_525),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_939),
.B(n_526),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_972),
.B(n_528),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_934),
.B(n_532),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_915),
.B(n_537),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_906),
.B(n_922),
.Y(n_1030)
);

NAND2xp33_ASAP7_75t_SL g1031 ( 
.A(n_889),
.B(n_932),
.Y(n_1031)
);

NAND2xp33_ASAP7_75t_SL g1032 ( 
.A(n_959),
.B(n_538),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_974),
.B(n_543),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_SL g1034 ( 
.A(n_960),
.B(n_545),
.Y(n_1034)
);

NAND2xp33_ASAP7_75t_SL g1035 ( 
.A(n_961),
.B(n_970),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_893),
.B(n_546),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_919),
.B(n_547),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_925),
.B(n_550),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_965),
.B(n_555),
.Y(n_1039)
);

NAND2xp33_ASAP7_75t_SL g1040 ( 
.A(n_971),
.B(n_557),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_951),
.B(n_560),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_953),
.B(n_561),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_956),
.B(n_564),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_949),
.B(n_567),
.Y(n_1044)
);

AND2x6_ASAP7_75t_SL g1045 ( 
.A(n_937),
.B(n_520),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_950),
.B(n_568),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_958),
.B(n_569),
.Y(n_1047)
);

NAND2xp33_ASAP7_75t_SL g1048 ( 
.A(n_909),
.B(n_570),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_915),
.B(n_571),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_947),
.B(n_948),
.Y(n_1050)
);

NAND2xp33_ASAP7_75t_SL g1051 ( 
.A(n_892),
.B(n_572),
.Y(n_1051)
);

NAND2xp33_ASAP7_75t_SL g1052 ( 
.A(n_880),
.B(n_573),
.Y(n_1052)
);

INVxp67_ASAP7_75t_L g1053 ( 
.A(n_1022),
.Y(n_1053)
);

INVxp67_ASAP7_75t_SL g1054 ( 
.A(n_998),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_977),
.A2(n_898),
.B(n_880),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1012),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_981),
.B(n_884),
.Y(n_1057)
);

AO31x2_ASAP7_75t_L g1058 ( 
.A1(n_994),
.A2(n_898),
.A3(n_884),
.B(n_881),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_982),
.A2(n_900),
.B(n_969),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_987),
.B(n_881),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_1012),
.Y(n_1061)
);

INVx5_ASAP7_75t_L g1062 ( 
.A(n_1045),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_1012),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_1052),
.A2(n_1048),
.B(n_1001),
.C(n_1020),
.Y(n_1064)
);

NOR4xp25_ASAP7_75t_L g1065 ( 
.A(n_1037),
.B(n_935),
.C(n_924),
.D(n_968),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_989),
.A2(n_1050),
.B(n_1024),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_1030),
.A2(n_1006),
.B(n_1007),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_978),
.A2(n_900),
.B(n_973),
.Y(n_1068)
);

NAND3xp33_ASAP7_75t_SL g1069 ( 
.A(n_990),
.B(n_544),
.C(n_531),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_1039),
.A2(n_895),
.B(n_577),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_SL g1071 ( 
.A1(n_1029),
.A2(n_465),
.B(n_574),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_1051),
.A2(n_882),
.B(n_465),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_1008),
.A2(n_895),
.B(n_441),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1000),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_986),
.Y(n_1075)
);

BUFx12f_ASAP7_75t_L g1076 ( 
.A(n_993),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_992),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1005),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_991),
.A2(n_895),
.B(n_441),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1025),
.B(n_1026),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1049),
.A2(n_882),
.B(n_465),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1010),
.Y(n_1082)
);

CKINVDCx6p67_ASAP7_75t_R g1083 ( 
.A(n_1033),
.Y(n_1083)
);

NAND3xp33_ASAP7_75t_L g1084 ( 
.A(n_979),
.B(n_891),
.C(n_890),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_1035),
.A2(n_967),
.A3(n_975),
.B(n_968),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1028),
.A2(n_967),
.B(n_582),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1014),
.A2(n_583),
.B(n_579),
.Y(n_1087)
);

O2A1O1Ixp5_ASAP7_75t_L g1088 ( 
.A1(n_1038),
.A2(n_975),
.B(n_935),
.C(n_924),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_1011),
.A2(n_56),
.B(n_49),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1017),
.A2(n_588),
.B(n_584),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1018),
.B(n_916),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1019),
.A2(n_565),
.B(n_558),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1047),
.A2(n_920),
.B(n_916),
.Y(n_1093)
);

NAND3xp33_ASAP7_75t_SL g1094 ( 
.A(n_996),
.B(n_576),
.C(n_575),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1013),
.Y(n_1095)
);

OA21x2_ASAP7_75t_L g1096 ( 
.A1(n_1021),
.A2(n_920),
.B(n_58),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_984),
.A2(n_62),
.B(n_57),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1002),
.A2(n_64),
.B(n_63),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_1003),
.A2(n_66),
.B(n_65),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_988),
.A2(n_70),
.B(n_67),
.Y(n_1100)
);

NAND2x1_ASAP7_75t_L g1101 ( 
.A(n_1031),
.B(n_71),
.Y(n_1101)
);

AND2x6_ASAP7_75t_L g1102 ( 
.A(n_983),
.B(n_72),
.Y(n_1102)
);

OR2x2_ASAP7_75t_L g1103 ( 
.A(n_1027),
.B(n_18),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_995),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_1036),
.A2(n_75),
.B(n_74),
.Y(n_1105)
);

AO31x2_ASAP7_75t_L g1106 ( 
.A1(n_999),
.A2(n_80),
.A3(n_82),
.B(n_76),
.Y(n_1106)
);

AO21x2_ASAP7_75t_L g1107 ( 
.A1(n_1023),
.A2(n_88),
.B(n_85),
.Y(n_1107)
);

AO31x2_ASAP7_75t_L g1108 ( 
.A1(n_997),
.A2(n_90),
.A3(n_92),
.B(n_89),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1044),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1046),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1041),
.A2(n_1043),
.B(n_1042),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1015),
.A2(n_94),
.B(n_93),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1004),
.B(n_19),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1032),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1034),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_1077),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1093),
.A2(n_985),
.B1(n_1009),
.B2(n_1040),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_1083),
.Y(n_1118)
);

OAI221xp5_ASAP7_75t_L g1119 ( 
.A1(n_1092),
.A2(n_980),
.B1(n_1016),
.B2(n_22),
.C(n_23),
.Y(n_1119)
);

OA21x2_ASAP7_75t_L g1120 ( 
.A1(n_1055),
.A2(n_1073),
.B(n_1066),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_1076),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_1063),
.Y(n_1122)
);

AO31x2_ASAP7_75t_L g1123 ( 
.A1(n_1072),
.A2(n_20),
.A3(n_21),
.B(n_22),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_1061),
.B(n_95),
.Y(n_1124)
);

NOR2xp67_ASAP7_75t_L g1125 ( 
.A(n_1053),
.B(n_391),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1067),
.A2(n_99),
.B(n_96),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1091),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1054),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_1128)
);

OA21x2_ASAP7_75t_L g1129 ( 
.A1(n_1057),
.A2(n_104),
.B(n_101),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1081),
.A2(n_26),
.A3(n_27),
.B(n_28),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1079),
.A2(n_110),
.B(n_108),
.Y(n_1131)
);

NOR2x1_ASAP7_75t_R g1132 ( 
.A(n_1062),
.B(n_111),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1097),
.A2(n_1099),
.B(n_1098),
.Y(n_1133)
);

AO31x2_ASAP7_75t_L g1134 ( 
.A1(n_1064),
.A2(n_27),
.A3(n_30),
.B(n_32),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_1103),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_1063),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1056),
.B(n_33),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1089),
.A2(n_1100),
.B(n_1105),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1074),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1060),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_1140)
);

BUFx2_ASAP7_75t_SL g1141 ( 
.A(n_1075),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1112),
.A2(n_116),
.B(n_115),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1078),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1095),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1082),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1069),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1080),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_1147)
);

NAND2x1_ASAP7_75t_L g1148 ( 
.A(n_1071),
.B(n_120),
.Y(n_1148)
);

INVx1_ASAP7_75t_SL g1149 ( 
.A(n_1109),
.Y(n_1149)
);

AO21x2_ASAP7_75t_L g1150 ( 
.A1(n_1070),
.A2(n_125),
.B(n_124),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1059),
.A2(n_129),
.B(n_128),
.Y(n_1151)
);

OAI211xp5_ASAP7_75t_L g1152 ( 
.A1(n_1065),
.A2(n_43),
.B(n_44),
.C(n_46),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_1104),
.B(n_44),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_1102),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1085),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1085),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1101),
.A2(n_132),
.B(n_130),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1110),
.B(n_46),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_1062),
.Y(n_1159)
);

OR2x6_ASAP7_75t_L g1160 ( 
.A(n_1068),
.B(n_133),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1101),
.A2(n_135),
.B(n_134),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1111),
.A2(n_138),
.B(n_136),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1058),
.Y(n_1163)
);

BUFx4_ASAP7_75t_SL g1164 ( 
.A(n_1084),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1058),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1115),
.B(n_139),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_SL g1167 ( 
.A1(n_1062),
.A2(n_47),
.B1(n_48),
.B2(n_140),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1102),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1085),
.Y(n_1169)
);

AO32x2_ASAP7_75t_L g1170 ( 
.A1(n_1058),
.A2(n_48),
.A3(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1086),
.A2(n_144),
.B(n_147),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_1094),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1102),
.Y(n_1173)
);

AOI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1114),
.A2(n_148),
.B(n_150),
.Y(n_1174)
);

INVx6_ASAP7_75t_L g1175 ( 
.A(n_1113),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1155),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1163),
.A2(n_1106),
.A3(n_1108),
.B(n_1096),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1124),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1124),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1145),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1165),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1144),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1136),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1139),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1143),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1156),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1169),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1117),
.B(n_1096),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1116),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1149),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1166),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1135),
.B(n_1166),
.Y(n_1192)
);

BUFx2_ASAP7_75t_SL g1193 ( 
.A(n_1118),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1152),
.B(n_1108),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1138),
.A2(n_1088),
.B(n_1087),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1168),
.B(n_1106),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1137),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1158),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_1122),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1160),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1134),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1120),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1134),
.Y(n_1203)
);

BUFx2_ASAP7_75t_SL g1204 ( 
.A(n_1159),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1172),
.A2(n_1175),
.B1(n_1173),
.B2(n_1119),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_1153),
.B(n_1090),
.Y(n_1206)
);

AOI221xp5_ASAP7_75t_L g1207 ( 
.A1(n_1147),
.A2(n_1140),
.B1(n_1128),
.B2(n_1146),
.C(n_1127),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1134),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1133),
.A2(n_1107),
.B(n_153),
.Y(n_1209)
);

INVxp67_ASAP7_75t_SL g1210 ( 
.A(n_1120),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1126),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1175),
.B(n_154),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1154),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1160),
.B(n_390),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1154),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1151),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1154),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1121),
.B(n_157),
.Y(n_1218)
);

INVx4_ASAP7_75t_SL g1219 ( 
.A(n_1123),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1123),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1148),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1162),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1167),
.A2(n_1141),
.B1(n_1125),
.B2(n_1170),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1123),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1131),
.A2(n_158),
.B(n_159),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1130),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1129),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1130),
.Y(n_1228)
);

AOI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1174),
.A2(n_163),
.B(n_164),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1157),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1129),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1161),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1130),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1171),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1170),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1150),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1142),
.B(n_1164),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1170),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1174),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1132),
.B(n_173),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1145),
.Y(n_1241)
);

OAI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1119),
.A2(n_176),
.B1(n_178),
.B2(n_182),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1145),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1119),
.A2(n_188),
.B1(n_192),
.B2(n_194),
.Y(n_1244)
);

BUFx2_ASAP7_75t_SL g1245 ( 
.A(n_1118),
.Y(n_1245)
);

NAND2xp33_ASAP7_75t_SL g1246 ( 
.A(n_1190),
.B(n_195),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1178),
.B(n_199),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1178),
.B(n_200),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1198),
.B(n_201),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1197),
.B(n_203),
.Y(n_1250)
);

NAND2xp33_ASAP7_75t_R g1251 ( 
.A(n_1240),
.B(n_207),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1205),
.B(n_1200),
.Y(n_1252)
);

XOR2xp5_ASAP7_75t_L g1253 ( 
.A(n_1193),
.B(n_208),
.Y(n_1253)
);

XOR2xp5_ASAP7_75t_L g1254 ( 
.A(n_1245),
.B(n_209),
.Y(n_1254)
);

NAND2xp33_ASAP7_75t_R g1255 ( 
.A(n_1240),
.B(n_210),
.Y(n_1255)
);

NAND2xp33_ASAP7_75t_SL g1256 ( 
.A(n_1192),
.B(n_211),
.Y(n_1256)
);

NAND2xp33_ASAP7_75t_R g1257 ( 
.A(n_1183),
.B(n_212),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_R g1258 ( 
.A(n_1179),
.B(n_389),
.Y(n_1258)
);

BUFx5_ASAP7_75t_L g1259 ( 
.A(n_1221),
.Y(n_1259)
);

INVxp67_ASAP7_75t_L g1260 ( 
.A(n_1189),
.Y(n_1260)
);

NAND2xp33_ASAP7_75t_R g1261 ( 
.A(n_1206),
.B(n_213),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1189),
.B(n_214),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1191),
.B(n_215),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1184),
.B(n_216),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1185),
.B(n_217),
.Y(n_1265)
);

NAND2xp33_ASAP7_75t_R g1266 ( 
.A(n_1237),
.B(n_219),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1180),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1241),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1182),
.B(n_220),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1204),
.Y(n_1270)
);

NAND2xp33_ASAP7_75t_R g1271 ( 
.A(n_1179),
.B(n_221),
.Y(n_1271)
);

NAND2xp33_ASAP7_75t_R g1272 ( 
.A(n_1213),
.B(n_1215),
.Y(n_1272)
);

OR2x6_ASAP7_75t_L g1273 ( 
.A(n_1218),
.B(n_223),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1187),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1243),
.B(n_224),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1213),
.B(n_225),
.Y(n_1276)
);

XNOR2xp5_ASAP7_75t_L g1277 ( 
.A(n_1218),
.B(n_388),
.Y(n_1277)
);

NAND2xp33_ASAP7_75t_SL g1278 ( 
.A(n_1217),
.B(n_226),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1212),
.B(n_227),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1215),
.B(n_1217),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1212),
.B(n_228),
.Y(n_1281)
);

BUFx10_ASAP7_75t_L g1282 ( 
.A(n_1217),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1214),
.B(n_229),
.Y(n_1283)
);

XNOR2xp5_ASAP7_75t_L g1284 ( 
.A(n_1199),
.B(n_231),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1214),
.B(n_232),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1186),
.Y(n_1286)
);

INVxp67_ASAP7_75t_L g1287 ( 
.A(n_1217),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1221),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1196),
.Y(n_1289)
);

XNOR2xp5_ASAP7_75t_L g1290 ( 
.A(n_1223),
.B(n_235),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1196),
.B(n_240),
.Y(n_1291)
);

NAND2xp33_ASAP7_75t_R g1292 ( 
.A(n_1194),
.B(n_241),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1176),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_R g1294 ( 
.A(n_1229),
.B(n_387),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1181),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1207),
.B(n_248),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1223),
.B(n_250),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_R g1298 ( 
.A(n_1194),
.B(n_251),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_R g1299 ( 
.A(n_1201),
.B(n_386),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1207),
.B(n_253),
.Y(n_1300)
);

INVxp67_ASAP7_75t_L g1301 ( 
.A(n_1176),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1244),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1181),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1203),
.Y(n_1304)
);

BUFx8_ASAP7_75t_L g1305 ( 
.A(n_1226),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_R g1306 ( 
.A(n_1208),
.B(n_385),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1195),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_1188),
.Y(n_1308)
);

AND2x4_ASAP7_75t_SL g1309 ( 
.A(n_1288),
.B(n_1220),
.Y(n_1309)
);

AOI21xp33_ASAP7_75t_L g1310 ( 
.A1(n_1296),
.A2(n_1242),
.B(n_1244),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1307),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1274),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1293),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1260),
.B(n_1188),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1252),
.B(n_1242),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1301),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1286),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1267),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1304),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1268),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1289),
.B(n_1228),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1308),
.B(n_1220),
.Y(n_1322)
);

OAI222xp33_ASAP7_75t_L g1323 ( 
.A1(n_1302),
.A2(n_1238),
.B1(n_1235),
.B2(n_1233),
.C1(n_1224),
.C2(n_1231),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1295),
.B(n_1219),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1300),
.B(n_1236),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1297),
.B(n_1262),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1291),
.B(n_1219),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1303),
.Y(n_1328)
);

AND2x4_ASAP7_75t_SL g1329 ( 
.A(n_1288),
.B(n_1231),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1287),
.B(n_1219),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1305),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1283),
.B(n_1239),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1285),
.B(n_1177),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1259),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1280),
.B(n_1177),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1259),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1290),
.B(n_1202),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1259),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1259),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1280),
.B(n_1177),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1275),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1269),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1264),
.B(n_1177),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1270),
.B(n_1227),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1249),
.B(n_1202),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1250),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1279),
.B(n_1210),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1265),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1281),
.B(n_1210),
.Y(n_1349)
);

INVxp67_ASAP7_75t_SL g1350 ( 
.A(n_1272),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1298),
.B(n_1230),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1263),
.B(n_1230),
.Y(n_1352)
);

NOR3xp33_ASAP7_75t_L g1353 ( 
.A(n_1246),
.B(n_1216),
.C(n_1234),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1284),
.B(n_1232),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1256),
.B(n_1222),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1292),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1312),
.Y(n_1357)
);

OR2x6_ASAP7_75t_L g1358 ( 
.A(n_1356),
.B(n_1273),
.Y(n_1358)
);

OAI221xp5_ASAP7_75t_L g1359 ( 
.A1(n_1315),
.A2(n_1251),
.B1(n_1255),
.B2(n_1261),
.C(n_1257),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1316),
.B(n_1253),
.Y(n_1360)
);

OAI322xp33_ASAP7_75t_L g1361 ( 
.A1(n_1315),
.A2(n_1314),
.A3(n_1356),
.B1(n_1346),
.B2(n_1341),
.C1(n_1342),
.C2(n_1325),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1329),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1335),
.B(n_1211),
.Y(n_1363)
);

NAND3xp33_ASAP7_75t_L g1364 ( 
.A(n_1325),
.B(n_1266),
.C(n_1271),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1312),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1318),
.B(n_1320),
.Y(n_1366)
);

INVxp67_ASAP7_75t_L g1367 ( 
.A(n_1319),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1322),
.B(n_1211),
.Y(n_1368)
);

AOI221xp5_ASAP7_75t_L g1369 ( 
.A1(n_1310),
.A2(n_1277),
.B1(n_1299),
.B2(n_1306),
.C(n_1254),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1332),
.B(n_1247),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1344),
.B(n_1282),
.Y(n_1371)
);

INVxp67_ASAP7_75t_L g1372 ( 
.A(n_1319),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1350),
.B(n_1258),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1313),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1354),
.B(n_1273),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1317),
.Y(n_1376)
);

OR2x2_ASAP7_75t_SL g1377 ( 
.A(n_1331),
.B(n_1278),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1329),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1343),
.B(n_1248),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1345),
.B(n_1347),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1353),
.A2(n_1294),
.B1(n_1276),
.B2(n_1225),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1340),
.B(n_1209),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1337),
.B(n_254),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1350),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1333),
.B(n_255),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1321),
.B(n_259),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1311),
.B(n_263),
.Y(n_1387)
);

OAI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1359),
.A2(n_1355),
.B1(n_1348),
.B2(n_1349),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1384),
.B(n_1311),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1357),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1362),
.B(n_1339),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1367),
.B(n_1317),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1365),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1365),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1367),
.B(n_1328),
.Y(n_1395)
);

NAND2x1p5_ASAP7_75t_L g1396 ( 
.A(n_1362),
.B(n_1336),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1363),
.B(n_1311),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1372),
.B(n_1339),
.Y(n_1398)
);

INVx4_ASAP7_75t_L g1399 ( 
.A(n_1358),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1374),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1372),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1376),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1376),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1380),
.B(n_1334),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1363),
.B(n_1324),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1366),
.B(n_1336),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1378),
.B(n_1324),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1368),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1388),
.A2(n_1364),
.B1(n_1373),
.B2(n_1358),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1407),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1404),
.B(n_1385),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1401),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1390),
.Y(n_1413)
);

NAND2xp33_ASAP7_75t_SL g1414 ( 
.A(n_1399),
.B(n_1373),
.Y(n_1414)
);

NAND2xp33_ASAP7_75t_SL g1415 ( 
.A(n_1399),
.B(n_1375),
.Y(n_1415)
);

OAI221xp5_ASAP7_75t_L g1416 ( 
.A1(n_1404),
.A2(n_1369),
.B1(n_1358),
.B2(n_1381),
.C(n_1370),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1391),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1408),
.B(n_1406),
.Y(n_1418)
);

NAND2xp33_ASAP7_75t_R g1419 ( 
.A(n_1389),
.B(n_1360),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1396),
.Y(n_1420)
);

OAI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1396),
.A2(n_1337),
.B1(n_1386),
.B2(n_1326),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1414),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1413),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_1415),
.Y(n_1424)
);

AND2x4_ASAP7_75t_SL g1425 ( 
.A(n_1409),
.B(n_1371),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1412),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1411),
.B(n_1400),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1418),
.B(n_1416),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1420),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1410),
.B(n_1406),
.Y(n_1430)
);

OAI21xp33_ASAP7_75t_L g1431 ( 
.A1(n_1421),
.A2(n_1383),
.B(n_1381),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1417),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1419),
.B(n_1397),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1421),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1413),
.Y(n_1435)
);

INVx3_ASAP7_75t_SL g1436 ( 
.A(n_1417),
.Y(n_1436)
);

AOI221x1_ASAP7_75t_L g1437 ( 
.A1(n_1431),
.A2(n_1398),
.B1(n_1395),
.B2(n_1392),
.C(n_1353),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1433),
.B(n_1405),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1429),
.B(n_1391),
.Y(n_1439)
);

OA211x2_ASAP7_75t_L g1440 ( 
.A1(n_1431),
.A2(n_1377),
.B(n_1398),
.C(n_1395),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1423),
.Y(n_1441)
);

AOI21xp33_ASAP7_75t_L g1442 ( 
.A1(n_1422),
.A2(n_1387),
.B(n_1392),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1428),
.A2(n_1387),
.B(n_1351),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1426),
.B(n_1424),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1435),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1441),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1445),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1444),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1444),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1437),
.B(n_1422),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1439),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1440),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1446),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1447),
.Y(n_1454)
);

INVx1_ASAP7_75t_SL g1455 ( 
.A(n_1448),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1449),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1451),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_1452),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1452),
.Y(n_1459)
);

NAND4xp25_ASAP7_75t_SL g1460 ( 
.A(n_1455),
.B(n_1450),
.C(n_1434),
.D(n_1440),
.Y(n_1460)
);

NAND4xp25_ASAP7_75t_L g1461 ( 
.A(n_1456),
.B(n_1432),
.C(n_1442),
.D(n_1443),
.Y(n_1461)
);

NOR3xp33_ASAP7_75t_L g1462 ( 
.A(n_1458),
.B(n_1361),
.C(n_1427),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1457),
.B(n_1436),
.Y(n_1463)
);

AND4x1_ASAP7_75t_L g1464 ( 
.A(n_1459),
.B(n_1438),
.C(n_1425),
.D(n_1351),
.Y(n_1464)
);

NAND4xp25_ASAP7_75t_L g1465 ( 
.A(n_1453),
.B(n_1430),
.C(n_1327),
.D(n_1330),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1454),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1458),
.B(n_1402),
.Y(n_1467)
);

NOR3xp33_ASAP7_75t_L g1468 ( 
.A(n_1458),
.B(n_1336),
.C(n_1338),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1466),
.Y(n_1469)
);

AOI322xp5_ASAP7_75t_L g1470 ( 
.A1(n_1462),
.A2(n_1379),
.A3(n_1394),
.B1(n_1393),
.B2(n_1382),
.C1(n_1403),
.C2(n_1323),
.Y(n_1470)
);

AOI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1460),
.A2(n_1338),
.B1(n_1309),
.B2(n_1352),
.C(n_268),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1463),
.Y(n_1472)
);

OA22x2_ASAP7_75t_L g1473 ( 
.A1(n_1467),
.A2(n_1309),
.B1(n_1338),
.B2(n_267),
.Y(n_1473)
);

XOR2xp5_ASAP7_75t_L g1474 ( 
.A(n_1461),
.B(n_264),
.Y(n_1474)
);

AOI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1465),
.A2(n_265),
.B1(n_269),
.B2(n_271),
.C(n_272),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1464),
.Y(n_1476)
);

NOR2x1_ASAP7_75t_L g1477 ( 
.A(n_1469),
.B(n_1468),
.Y(n_1477)
);

XOR2xp5_ASAP7_75t_L g1478 ( 
.A(n_1474),
.B(n_275),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1476),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1472),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1473),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1471),
.B(n_276),
.Y(n_1482)
);

NOR2x1_ASAP7_75t_L g1483 ( 
.A(n_1475),
.B(n_278),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1470),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1479),
.B(n_279),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_SL g1486 ( 
.A(n_1477),
.B(n_1481),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1484),
.B(n_280),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1480),
.B(n_281),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1478),
.B(n_282),
.Y(n_1489)
);

NAND2xp33_ASAP7_75t_SL g1490 ( 
.A(n_1482),
.B(n_283),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_1483),
.B(n_284),
.C(n_285),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1486),
.B(n_286),
.Y(n_1492)
);

INVx1_ASAP7_75t_SL g1493 ( 
.A(n_1490),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1485),
.Y(n_1494)
);

NAND5xp2_ASAP7_75t_L g1495 ( 
.A(n_1487),
.B(n_288),
.C(n_290),
.D(n_291),
.E(n_292),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1489),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1491),
.A2(n_293),
.B1(n_295),
.B2(n_298),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1494),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1496),
.Y(n_1499)
);

NOR2x1_ASAP7_75t_L g1500 ( 
.A(n_1492),
.B(n_1488),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1493),
.Y(n_1501)
);

OAI22x1_ASAP7_75t_L g1502 ( 
.A1(n_1497),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1495),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1501),
.B(n_304),
.Y(n_1504)
);

INVx4_ASAP7_75t_L g1505 ( 
.A(n_1499),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1503),
.A2(n_305),
.B1(n_307),
.B2(n_308),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1498),
.A2(n_310),
.B1(n_311),
.B2(n_313),
.Y(n_1507)
);

AOI31xp33_ASAP7_75t_L g1508 ( 
.A1(n_1504),
.A2(n_1500),
.A3(n_1502),
.B(n_317),
.Y(n_1508)
);

AOI31xp33_ASAP7_75t_L g1509 ( 
.A1(n_1506),
.A2(n_314),
.A3(n_315),
.B(n_318),
.Y(n_1509)
);

OAI322xp33_ASAP7_75t_L g1510 ( 
.A1(n_1508),
.A2(n_1505),
.A3(n_1507),
.B1(n_331),
.B2(n_332),
.C1(n_335),
.C2(n_336),
.Y(n_1510)
);

OAI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1509),
.A2(n_319),
.B1(n_328),
.B2(n_337),
.Y(n_1511)
);

OAI221xp5_ASAP7_75t_L g1512 ( 
.A1(n_1510),
.A2(n_338),
.B1(n_343),
.B2(n_345),
.C(n_346),
.Y(n_1512)
);

AOI222xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1511),
.A2(n_347),
.B1(n_348),
.B2(n_350),
.C1(n_351),
.C2(n_353),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1512),
.Y(n_1514)
);

AOI221xp5_ASAP7_75t_L g1515 ( 
.A1(n_1514),
.A2(n_1513),
.B1(n_358),
.B2(n_359),
.C(n_361),
.Y(n_1515)
);

AOI211xp5_ASAP7_75t_L g1516 ( 
.A1(n_1515),
.A2(n_356),
.B(n_362),
.C(n_363),
.Y(n_1516)
);


endmodule