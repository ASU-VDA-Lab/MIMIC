module fake_jpeg_25630_n_322 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_59),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_30),
.B1(n_19),
.B2(n_22),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_66),
.B1(n_40),
.B2(n_39),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_30),
.B1(n_22),
.B2(n_19),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_50),
.A2(n_54),
.B1(n_20),
.B2(n_32),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_24),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_30),
.B1(n_19),
.B2(n_22),
.Y(n_54)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_58),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_25),
.B1(n_34),
.B2(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_29),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_41),
.Y(n_86)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_69),
.Y(n_93)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_39),
.C(n_41),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_77),
.C(n_60),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_95),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_75),
.B(n_79),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_41),
.C(n_37),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_18),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_94),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_18),
.B(n_28),
.C(n_31),
.Y(n_84)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_56),
.A3(n_46),
.B1(n_33),
.B2(n_24),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_28),
.B1(n_31),
.B2(n_40),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g117 ( 
.A(n_85),
.B(n_88),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_37),
.Y(n_103)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_62),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_46),
.A2(n_20),
.B1(n_21),
.B2(n_32),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_92),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_62),
.B1(n_69),
.B2(n_64),
.Y(n_96)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_29),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_29),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_96),
.A2(n_109),
.B1(n_79),
.B2(n_87),
.Y(n_125)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_100),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_24),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_99),
.B(n_119),
.Y(n_128)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_108),
.Y(n_152)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_110),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_104),
.A2(n_106),
.B(n_114),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_29),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_68),
.B1(n_61),
.B2(n_47),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_92),
.B1(n_90),
.B2(n_80),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_83),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_61),
.B1(n_47),
.B2(n_20),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_112),
.Y(n_130)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_29),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_60),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_120),
.Y(n_135)
);

BUFx10_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_27),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_106),
.B(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_82),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_115),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_124),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_97),
.B1(n_101),
.B2(n_78),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_113),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_126),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_123),
.B(n_74),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_127),
.B(n_136),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_140),
.B1(n_120),
.B2(n_112),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_138),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_137),
.B(n_114),
.Y(n_154)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_98),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_100),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_143),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_122),
.B1(n_103),
.B2(n_106),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_144),
.B1(n_109),
.B2(n_111),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_83),
.C(n_70),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_89),
.C(n_63),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_81),
.Y(n_147)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_99),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_160),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_154),
.A2(n_156),
.B(n_168),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_155),
.A2(n_161),
.B1(n_169),
.B2(n_146),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_117),
.B(n_110),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_173),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_159),
.A2(n_174),
.B1(n_182),
.B2(n_131),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_58),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_80),
.B1(n_81),
.B2(n_89),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_162),
.B(n_167),
.Y(n_189)
);

INVxp33_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_181),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_58),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_171),
.Y(n_209)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_0),
.B(n_1),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_20),
.B1(n_32),
.B2(n_21),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_23),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_134),
.B(n_129),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_125),
.A2(n_138),
.B1(n_149),
.B2(n_137),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_27),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_177),
.C(n_180),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_63),
.C(n_72),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_130),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_127),
.A2(n_118),
.B1(n_21),
.B2(n_27),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_33),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_188),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_178),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_187),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_124),
.Y(n_188)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_193),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_191),
.A2(n_195),
.B1(n_205),
.B2(n_156),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_192),
.A2(n_206),
.B1(n_210),
.B2(n_33),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_172),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_159),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_201),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_155),
.A2(n_126),
.B1(n_135),
.B2(n_133),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_147),
.Y(n_197)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_130),
.Y(n_198)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_153),
.Y(n_217)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_152),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_202),
.A2(n_186),
.B(n_208),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_140),
.Y(n_204)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_166),
.A2(n_133),
.B1(n_144),
.B2(n_146),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_139),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_166),
.B1(n_168),
.B2(n_173),
.Y(n_211)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_165),
.C(n_175),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_219),
.C(n_223),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_227),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_217),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_171),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_177),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_232),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_SL g225 ( 
.A(n_199),
.B(n_156),
.C(n_154),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_225),
.A2(n_208),
.B(n_202),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_183),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_234),
.C(n_209),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_206),
.A2(n_146),
.B1(n_158),
.B2(n_118),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_229),
.A2(n_231),
.B1(n_235),
.B2(n_190),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_195),
.A2(n_118),
.B1(n_10),
.B2(n_11),
.Y(n_230)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_230),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_191),
.A2(n_186),
.B1(n_210),
.B2(n_205),
.Y(n_231)
);

FAx1_ASAP7_75t_SL g232 ( 
.A(n_204),
.B(n_33),
.CI(n_10),
.CON(n_232),
.SN(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_33),
.C(n_9),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_216),
.B(n_197),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_247),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_213),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_251),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_238),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_184),
.Y(n_243)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_244),
.A2(n_220),
.B1(n_1),
.B2(n_2),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_200),
.C(n_202),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_250),
.C(n_219),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_246),
.A2(n_252),
.B(n_11),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_221),
.B(n_198),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_192),
.C(n_9),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_214),
.A2(n_9),
.B(n_15),
.Y(n_252)
);

BUFx24_ASAP7_75t_SL g253 ( 
.A(n_232),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_0),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_256),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_227),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_258),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_217),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_228),
.C(n_231),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_271),
.C(n_6),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_263),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_234),
.Y(n_263)
);

AO221x1_ASAP7_75t_L g265 ( 
.A1(n_255),
.A2(n_235),
.B1(n_232),
.B2(n_233),
.C(n_218),
.Y(n_265)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_266),
.A2(n_241),
.B(n_12),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_268),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_252),
.A2(n_8),
.B(n_15),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_270),
.A2(n_11),
.B(n_16),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_8),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_260),
.A2(n_244),
.B1(n_236),
.B2(n_255),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_280),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_254),
.Y(n_274)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_239),
.Y(n_276)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_278),
.B(n_279),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_272),
.B(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_283),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_242),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_285),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_286),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_259),
.C(n_257),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_290),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_261),
.C(n_258),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_297),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_263),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_285),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_275),
.A2(n_274),
.B(n_278),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_296),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_271),
.C(n_267),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_14),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_294),
.B(n_273),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_302),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_286),
.Y(n_302)
);

AOI21xp33_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_12),
.B(n_13),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_305),
.A2(n_3),
.B(n_4),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_12),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_307),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_13),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_299),
.A2(n_287),
.B1(n_293),
.B2(n_297),
.Y(n_309)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_309),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_288),
.B1(n_290),
.B2(n_295),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_310),
.B(n_312),
.Y(n_316)
);

NAND4xp25_ASAP7_75t_SL g317 ( 
.A(n_313),
.B(n_314),
.C(n_305),
.D(n_4),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_300),
.A2(n_14),
.B1(n_16),
.B2(n_3),
.Y(n_314)
);

AO21x1_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_308),
.B(n_311),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_318),
.B(n_315),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_316),
.C(n_303),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_309),
.B(n_312),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_16),
.Y(n_322)
);


endmodule