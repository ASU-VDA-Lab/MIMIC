module fake_ibex_1061_n_2077 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_403, n_423, n_357, n_88, n_412, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_421, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_407, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_199, n_410, n_308, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_385, n_414, n_118, n_378, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_408, n_119, n_361, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_393, n_297, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_2077);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_407;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_410;
input n_308;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_118;
input n_378;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_393;
input n_297;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;

output n_2077;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_766;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_1930;
wire n_452;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_1971;
wire n_879;
wire n_1957;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_641;
wire n_557;
wire n_1937;
wire n_893;
wire n_527;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_431;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_2025;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_745;
wire n_447;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_971;
wire n_702;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_1936;
wire n_1717;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_737;
wire n_606;
wire n_1571;
wire n_1980;
wire n_462;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2076;
wire n_974;
wire n_1036;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2006;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_585;
wire n_1982;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_2010;
wire n_1470;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1806;
wire n_1539;
wire n_650;
wire n_1575;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_951;
wire n_2053;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2064;
wire n_1679;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_1353;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_1830;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_1725;
wire n_1135;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_1946;
wire n_1726;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_934;
wire n_520;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_1956;
wire n_681;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_858;
wire n_1018;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_786;
wire n_505;
wire n_2043;
wire n_1621;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1433;
wire n_1314;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1893;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1961;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1542;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_753;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_1892;
wire n_1061;
wire n_682;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_886;
wire n_1010;
wire n_883;
wire n_2044;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1635;
wire n_1572;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_2013;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_1868;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_581;
wire n_1472;
wire n_1365;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_519;
wire n_1843;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_1902;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1849;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;
wire n_425;

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_22),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_262),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_57),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_192),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_27),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_416),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_167),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_120),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_214),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_93),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_91),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_366),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_383),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_254),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_409),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_399),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_327),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_349),
.Y(n_441)
);

BUFx10_ASAP7_75t_L g442 ( 
.A(n_120),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_261),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_354),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_374),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_243),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_69),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_321),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_196),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_324),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_252),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_200),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_355),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_79),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_317),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_397),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_242),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_51),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_229),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_198),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_405),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_169),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_94),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_249),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_361),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_170),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_101),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_306),
.Y(n_469)
);

INVxp33_ASAP7_75t_SL g470 ( 
.A(n_379),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_97),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_403),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_401),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_363),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_419),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_272),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_286),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_372),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_168),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_386),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_338),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_160),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_398),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_332),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_158),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_358),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_143),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_289),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_141),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_411),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_381),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_422),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_61),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_141),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_86),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_65),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_382),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_216),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_167),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_74),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_310),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_415),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_58),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_219),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_311),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_304),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_375),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_345),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_173),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_4),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_402),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_408),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_296),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_124),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_55),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_69),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_352),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_283),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_202),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_204),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_239),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_136),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_235),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_171),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_110),
.Y(n_525)
);

BUFx10_ASAP7_75t_L g526 ( 
.A(n_362),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_226),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_423),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_117),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_106),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_64),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_151),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_84),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_117),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_68),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_207),
.Y(n_536)
);

INVxp33_ASAP7_75t_L g537 ( 
.A(n_181),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_249),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_19),
.Y(n_539)
);

NOR2xp67_ASAP7_75t_L g540 ( 
.A(n_333),
.B(n_344),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_370),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_376),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_149),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_242),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_19),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_284),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_342),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_418),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_307),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_407),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_203),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_293),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_420),
.Y(n_553)
);

INVxp67_ASAP7_75t_SL g554 ( 
.A(n_292),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_334),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_168),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_309),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_357),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_79),
.B(n_54),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_119),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_339),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_111),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_22),
.Y(n_563)
);

INVxp67_ASAP7_75t_SL g564 ( 
.A(n_268),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_390),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_303),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_235),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_313),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_73),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_132),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_63),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_74),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_140),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_46),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_325),
.Y(n_575)
);

CKINVDCx14_ASAP7_75t_R g576 ( 
.A(n_412),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_368),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_56),
.Y(n_578)
);

CKINVDCx14_ASAP7_75t_R g579 ( 
.A(n_97),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_160),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_367),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_343),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_59),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_275),
.Y(n_584)
);

NOR2xp67_ASAP7_75t_L g585 ( 
.A(n_59),
.B(n_197),
.Y(n_585)
);

INVx4_ASAP7_75t_R g586 ( 
.A(n_232),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_348),
.Y(n_587)
);

CKINVDCx16_ASAP7_75t_R g588 ( 
.A(n_247),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_276),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_156),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_67),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_94),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_365),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_154),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_172),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_346),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_102),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_131),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_83),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_203),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_89),
.Y(n_601)
);

INVxp33_ASAP7_75t_SL g602 ( 
.A(n_116),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_392),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_285),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_112),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_177),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_267),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_1),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_111),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_326),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_299),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_391),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_184),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_52),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_48),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_380),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_199),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_163),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_209),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_27),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_360),
.Y(n_621)
);

NOR2xp67_ASAP7_75t_L g622 ( 
.A(n_185),
.B(n_369),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_410),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_78),
.B(n_278),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_52),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_91),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_25),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_23),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_295),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_340),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_315),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_359),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_72),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_149),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_44),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_56),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_156),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_205),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_226),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_75),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_388),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_319),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_356),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_6),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_122),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_329),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_353),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_29),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_202),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_257),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_211),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_24),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_23),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_53),
.B(n_252),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_347),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_31),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_140),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_7),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_400),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_46),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_335),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_40),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_132),
.Y(n_663)
);

NOR2xp67_ASAP7_75t_L g664 ( 
.A(n_294),
.B(n_341),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_421),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_377),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_70),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_80),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_40),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_295),
.Y(n_670)
);

CKINVDCx14_ASAP7_75t_R g671 ( 
.A(n_301),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_302),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_186),
.Y(n_673)
);

NOR2xp67_ASAP7_75t_L g674 ( 
.A(n_417),
.B(n_184),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_300),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_123),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_114),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_364),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_150),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_378),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_42),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_179),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_54),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_188),
.Y(n_684)
);

CKINVDCx14_ASAP7_75t_R g685 ( 
.A(n_115),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_41),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_128),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_250),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_218),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_238),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_323),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_304),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_190),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_387),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_128),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_0),
.Y(n_696)
);

BUFx10_ASAP7_75t_L g697 ( 
.A(n_253),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_123),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_178),
.Y(n_699)
);

INVxp67_ASAP7_75t_L g700 ( 
.A(n_351),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_50),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_300),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_328),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_393),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_157),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_113),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_179),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_16),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_389),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_223),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_350),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_503),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_579),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_503),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_671),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_443),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_685),
.A2(n_8),
.B1(n_3),
.B2(n_5),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_463),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_443),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_508),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_525),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_517),
.B(n_5),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_508),
.Y(n_723)
);

OAI22x1_ASAP7_75t_R g724 ( 
.A1(n_448),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_457),
.Y(n_725)
);

BUFx8_ASAP7_75t_SL g726 ( 
.A(n_448),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_578),
.B(n_11),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_608),
.B(n_668),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_508),
.Y(n_729)
);

INVx5_ASAP7_75t_L g730 ( 
.A(n_526),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_608),
.B(n_12),
.Y(n_731)
);

OAI22x1_ASAP7_75t_SL g732 ( 
.A1(n_467),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_442),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_466),
.Y(n_734)
);

INVx5_ASAP7_75t_L g735 ( 
.A(n_526),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_512),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_547),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_508),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_668),
.Y(n_739)
);

AND2x6_ASAP7_75t_L g740 ( 
.A(n_466),
.B(n_314),
.Y(n_740)
);

CKINVDCx11_ASAP7_75t_R g741 ( 
.A(n_467),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_584),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_688),
.B(n_14),
.Y(n_743)
);

AND2x6_ASAP7_75t_L g744 ( 
.A(n_474),
.B(n_316),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_701),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_701),
.B(n_15),
.Y(n_746)
);

BUFx8_ASAP7_75t_SL g747 ( 
.A(n_539),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_561),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_551),
.B(n_17),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_561),
.Y(n_750)
);

CKINVDCx16_ASAP7_75t_R g751 ( 
.A(n_447),
.Y(n_751)
);

OA21x2_ASAP7_75t_L g752 ( 
.A1(n_547),
.A2(n_320),
.B(n_318),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_631),
.Y(n_753)
);

BUFx12f_ASAP7_75t_L g754 ( 
.A(n_526),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_602),
.A2(n_21),
.B1(n_18),
.B2(n_20),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_593),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_553),
.Y(n_757)
);

BUFx8_ASAP7_75t_L g758 ( 
.A(n_709),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_553),
.A2(n_703),
.B(n_435),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_551),
.B(n_20),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_SL g761 ( 
.A1(n_539),
.A2(n_25),
.B1(n_21),
.B2(n_24),
.Y(n_761)
);

INVx5_ASAP7_75t_L g762 ( 
.A(n_655),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_483),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_537),
.B(n_26),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_655),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_483),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_655),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_574),
.B(n_26),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_571),
.B(n_28),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_565),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_505),
.B(n_28),
.Y(n_771)
);

OA21x2_ASAP7_75t_L g772 ( 
.A1(n_436),
.A2(n_441),
.B(n_439),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_655),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_546),
.B(n_30),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_588),
.B(n_442),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_442),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_602),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_474),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_655),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_573),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_545),
.B(n_32),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_480),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_498),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_498),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_470),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_544),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_596),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_589),
.B(n_33),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_596),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_589),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_611),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_611),
.B(n_35),
.Y(n_792)
);

AND2x6_ASAP7_75t_L g793 ( 
.A(n_445),
.B(n_322),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_446),
.B(n_36),
.Y(n_794)
);

INVx5_ASAP7_75t_L g795 ( 
.A(n_498),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_498),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_449),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_451),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_615),
.Y(n_799)
);

OA21x2_ASAP7_75t_L g800 ( 
.A1(n_462),
.A2(n_331),
.B(n_330),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_498),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_536),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_749),
.B(n_475),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_749),
.Y(n_804)
);

INVxp67_ASAP7_75t_SL g805 ( 
.A(n_780),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_731),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_718),
.B(n_706),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_749),
.B(n_478),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_730),
.B(n_444),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_760),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_759),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_783),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_783),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_730),
.B(n_700),
.Y(n_814)
);

NAND3xp33_ASAP7_75t_L g815 ( 
.A(n_764),
.B(n_601),
.C(n_562),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_783),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_775),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_720),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_784),
.Y(n_819)
);

INVxp33_ASAP7_75t_SL g820 ( 
.A(n_742),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_760),
.B(n_490),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_746),
.Y(n_822)
);

OR2x6_ASAP7_75t_L g823 ( 
.A(n_754),
.B(n_585),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_735),
.Y(n_824)
);

INVx1_ASAP7_75t_SL g825 ( 
.A(n_751),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_746),
.A2(n_769),
.B1(n_788),
.B2(n_760),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_769),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_769),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_733),
.B(n_450),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_788),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_796),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_735),
.B(n_491),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_796),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_788),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_801),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_735),
.B(n_450),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_756),
.B(n_497),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_790),
.B(n_576),
.Y(n_838)
);

INVxp67_ASAP7_75t_SL g839 ( 
.A(n_780),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_801),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_792),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_801),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_754),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_728),
.B(n_502),
.Y(n_844)
);

INVx4_ASAP7_75t_L g845 ( 
.A(n_740),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_792),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_801),
.Y(n_847)
);

BUFx10_ASAP7_75t_L g848 ( 
.A(n_728),
.Y(n_848)
);

INVx8_ASAP7_75t_L g849 ( 
.A(n_740),
.Y(n_849)
);

CKINVDCx6p67_ASAP7_75t_R g850 ( 
.A(n_741),
.Y(n_850)
);

AND3x2_ASAP7_75t_L g851 ( 
.A(n_771),
.B(n_724),
.C(n_554),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_791),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_712),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_733),
.B(n_453),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_795),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_763),
.Y(n_856)
);

BUFx16f_ASAP7_75t_R g857 ( 
.A(n_758),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_797),
.B(n_511),
.Y(n_858)
);

INVx5_ASAP7_75t_L g859 ( 
.A(n_740),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_758),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_795),
.Y(n_861)
);

INVx4_ASAP7_75t_L g862 ( 
.A(n_740),
.Y(n_862)
);

NAND3xp33_ASAP7_75t_L g863 ( 
.A(n_764),
.B(n_673),
.C(n_706),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_795),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_762),
.Y(n_865)
);

BUFx10_ASAP7_75t_L g866 ( 
.A(n_776),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_714),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_721),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_762),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_797),
.B(n_528),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_762),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_802),
.B(n_458),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_734),
.Y(n_873)
);

OAI22xp33_ASAP7_75t_L g874 ( 
.A1(n_713),
.A2(n_458),
.B1(n_460),
.B2(n_459),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_739),
.B(n_459),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_763),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_798),
.B(n_542),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_762),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_766),
.B(n_460),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_720),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_720),
.Y(n_881)
);

AOI21x1_ASAP7_75t_L g882 ( 
.A1(n_772),
.A2(n_558),
.B(n_550),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_723),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_770),
.B(n_464),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_798),
.B(n_568),
.Y(n_885)
);

AND3x2_ASAP7_75t_L g886 ( 
.A(n_722),
.B(n_564),
.C(n_424),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_723),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_772),
.A2(n_426),
.B1(n_430),
.B2(n_425),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_723),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_778),
.B(n_575),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_778),
.B(n_577),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_729),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_799),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_729),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_729),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_727),
.B(n_710),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_729),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_748),
.B(n_536),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_738),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_738),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_716),
.Y(n_901)
);

AND2x6_ASAP7_75t_L g902 ( 
.A(n_744),
.B(n_581),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_738),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_719),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_782),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_719),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_782),
.B(n_787),
.Y(n_907)
);

OAI22xp33_ASAP7_75t_L g908 ( 
.A1(n_785),
.A2(n_471),
.B1(n_476),
.B2(n_468),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_787),
.B(n_587),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_765),
.Y(n_910)
);

NAND2xp33_ASAP7_75t_SL g911 ( 
.A(n_774),
.B(n_631),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_789),
.B(n_603),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_789),
.B(n_623),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_L g914 ( 
.A(n_744),
.B(n_438),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_765),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_725),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_765),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_767),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_767),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_736),
.B(n_630),
.Y(n_920)
);

NAND3xp33_ASAP7_75t_L g921 ( 
.A(n_743),
.B(n_477),
.C(n_476),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_737),
.B(n_632),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_741),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_767),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_768),
.A2(n_614),
.B1(n_619),
.B2(n_479),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_757),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_726),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_781),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_767),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_794),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_773),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_750),
.B(n_479),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_753),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_773),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_744),
.B(n_614),
.Y(n_935)
);

NAND3xp33_ASAP7_75t_L g936 ( 
.A(n_794),
.B(n_620),
.C(n_619),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_786),
.B(n_536),
.Y(n_937)
);

NOR2x1p5_ASAP7_75t_L g938 ( 
.A(n_726),
.B(n_695),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_793),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_793),
.B(n_620),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_793),
.B(n_626),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_826),
.A2(n_777),
.B1(n_755),
.B2(n_745),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_845),
.B(n_862),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_928),
.B(n_440),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_853),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_806),
.A2(n_793),
.B1(n_432),
.B2(n_433),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_805),
.B(n_839),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_845),
.B(n_862),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_SL g949 ( 
.A(n_862),
.B(n_761),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_807),
.B(n_626),
.Y(n_950)
);

NAND3xp33_ASAP7_75t_L g951 ( 
.A(n_925),
.B(n_717),
.C(n_715),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_817),
.B(n_697),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_867),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_850),
.Y(n_954)
);

OAI22xp33_ASAP7_75t_L g955 ( 
.A1(n_852),
.A2(n_560),
.B1(n_569),
.B2(n_544),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_908),
.A2(n_635),
.B1(n_650),
.B2(n_628),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_854),
.B(n_456),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_868),
.Y(n_958)
);

NAND3xp33_ASAP7_75t_L g959 ( 
.A(n_888),
.B(n_667),
.C(n_651),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_872),
.B(n_472),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_848),
.B(n_844),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_914),
.A2(n_752),
.B(n_800),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_825),
.B(n_651),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_844),
.B(n_473),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_809),
.B(n_481),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_838),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_830),
.A2(n_654),
.B1(n_559),
.B2(n_667),
.Y(n_967)
);

OR2x6_ASAP7_75t_L g968 ( 
.A(n_860),
.B(n_938),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_836),
.B(n_822),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_896),
.B(n_484),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_930),
.B(n_484),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_856),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_863),
.B(n_486),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_829),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_856),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_856),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_875),
.B(n_555),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_876),
.Y(n_978)
);

BUFx8_ASAP7_75t_L g979 ( 
.A(n_843),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_879),
.B(n_616),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_837),
.B(n_621),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_849),
.Y(n_982)
);

AO22x1_ASAP7_75t_L g983 ( 
.A1(n_820),
.A2(n_923),
.B1(n_927),
.B2(n_933),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_837),
.B(n_621),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_841),
.B(n_803),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_921),
.B(n_793),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_808),
.B(n_821),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_874),
.A2(n_696),
.B1(n_695),
.B2(n_428),
.Y(n_988)
);

AOI221xp5_ASAP7_75t_L g989 ( 
.A1(n_820),
.A2(n_732),
.B1(n_696),
.B2(n_455),
.C(n_461),
.Y(n_989)
);

AO22x2_ASAP7_75t_L g990 ( 
.A1(n_821),
.A2(n_437),
.B1(n_465),
.B2(n_452),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_884),
.B(n_642),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_815),
.B(n_643),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_804),
.A2(n_482),
.B1(n_489),
.B2(n_487),
.Y(n_993)
);

NAND2xp33_ASAP7_75t_L g994 ( 
.A(n_849),
.B(n_646),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_810),
.B(n_691),
.Y(n_995)
);

INVx8_ASAP7_75t_L g996 ( 
.A(n_849),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_932),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_893),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_906),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_866),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_873),
.B(n_694),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_810),
.A2(n_615),
.B(n_493),
.C(n_499),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_866),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_901),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_859),
.B(n_939),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_904),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_940),
.B(n_641),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_937),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_941),
.B(n_647),
.Y(n_1009)
);

NAND3xp33_ASAP7_75t_SL g1010 ( 
.A(n_936),
.B(n_431),
.C(n_427),
.Y(n_1010)
);

NAND3xp33_ASAP7_75t_L g1011 ( 
.A(n_914),
.B(n_488),
.C(n_434),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_898),
.B(n_697),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_827),
.B(n_659),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_828),
.B(n_666),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_823),
.B(n_496),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_859),
.B(n_492),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_834),
.A2(n_510),
.B1(n_514),
.B2(n_506),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_935),
.A2(n_870),
.B(n_877),
.C(n_858),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_823),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_926),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_846),
.B(n_507),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_823),
.B(n_697),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_823),
.B(n_494),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_814),
.B(n_824),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_905),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_902),
.A2(n_524),
.B1(n_529),
.B2(n_523),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_911),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_916),
.A2(n_504),
.B1(n_513),
.B2(n_501),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_814),
.B(n_678),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_849),
.A2(n_516),
.B1(n_518),
.B2(n_515),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_907),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_811),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_902),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_858),
.B(n_870),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_911),
.A2(n_705),
.B1(n_699),
.B2(n_522),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_902),
.A2(n_909),
.B1(n_877),
.B2(n_885),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_832),
.B(n_541),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_832),
.B(n_548),
.Y(n_1038)
);

NAND3xp33_ASAP7_75t_L g1039 ( 
.A(n_886),
.B(n_531),
.C(n_521),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_890),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_890),
.B(n_582),
.Y(n_1041)
);

OR2x6_ASAP7_75t_L g1042 ( 
.A(n_857),
.B(n_485),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_891),
.B(n_429),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_850),
.Y(n_1044)
);

INVx4_ASAP7_75t_L g1045 ( 
.A(n_865),
.Y(n_1045)
);

OAI221xp5_ASAP7_75t_L g1046 ( 
.A1(n_920),
.A2(n_538),
.B1(n_629),
.B2(n_495),
.C(n_469),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_912),
.B(n_610),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_913),
.B(n_612),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_922),
.B(n_454),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_922),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_882),
.B(n_661),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_927),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_869),
.B(n_665),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_855),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_851),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_869),
.B(n_680),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_871),
.B(n_532),
.Y(n_1057)
);

AOI221xp5_ASAP7_75t_L g1058 ( 
.A1(n_855),
.A2(n_557),
.B1(n_563),
.B2(n_556),
.C(n_552),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_861),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_878),
.B(n_704),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_878),
.B(n_711),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_864),
.B(n_533),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_812),
.Y(n_1063)
);

NAND3xp33_ASAP7_75t_L g1064 ( 
.A(n_813),
.B(n_535),
.C(n_534),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_881),
.B(n_566),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_816),
.B(n_633),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_819),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_819),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_818),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_881),
.B(n_567),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_831),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_SL g1072 ( 
.A(n_831),
.B(n_560),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_SL g1073 ( 
.A(n_833),
.B(n_569),
.Y(n_1073)
);

NOR2x1p5_ASAP7_75t_L g1074 ( 
.A(n_833),
.B(n_747),
.Y(n_1074)
);

NOR3xp33_ASAP7_75t_L g1075 ( 
.A(n_835),
.B(n_648),
.C(n_636),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_840),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_842),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_842),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_847),
.Y(n_1079)
);

INVx4_ASAP7_75t_L g1080 ( 
.A(n_880),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_883),
.A2(n_752),
.B(n_800),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_887),
.B(n_570),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_880),
.B(n_500),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_889),
.B(n_572),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_892),
.A2(n_590),
.B1(n_591),
.B2(n_580),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_895),
.B(n_592),
.Y(n_1086)
);

INVxp33_ASAP7_75t_SL g1087 ( 
.A(n_897),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_897),
.A2(n_597),
.B1(n_605),
.B2(n_595),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_899),
.B(n_583),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_894),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_900),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_900),
.A2(n_752),
.B(n_800),
.Y(n_1092)
);

NOR3xp33_ASAP7_75t_L g1093 ( 
.A(n_903),
.B(n_624),
.C(n_598),
.Y(n_1093)
);

INVxp67_ASAP7_75t_L g1094 ( 
.A(n_903),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_942),
.A2(n_967),
.B(n_1002),
.C(n_947),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1031),
.B(n_600),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1032),
.Y(n_1097)
);

BUFx8_ASAP7_75t_L g1098 ( 
.A(n_1052),
.Y(n_1098)
);

CKINVDCx8_ASAP7_75t_R g1099 ( 
.A(n_954),
.Y(n_1099)
);

AND2x6_ASAP7_75t_SL g1100 ( 
.A(n_1042),
.B(n_747),
.Y(n_1100)
);

INVx11_ASAP7_75t_L g1101 ( 
.A(n_979),
.Y(n_1101)
);

CKINVDCx11_ASAP7_75t_R g1102 ( 
.A(n_1042),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_996),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_996),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_944),
.B(n_974),
.Y(n_1105)
);

OR2x2_ASAP7_75t_L g1106 ( 
.A(n_955),
.B(n_786),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_963),
.Y(n_1107)
);

NAND3xp33_ASAP7_75t_L g1108 ( 
.A(n_1075),
.B(n_613),
.C(n_604),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_997),
.B(n_594),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_945),
.B(n_657),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_1000),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_953),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_950),
.B(n_594),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1081),
.A2(n_540),
.B(n_622),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_943),
.A2(n_915),
.B(n_910),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_996),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_958),
.B(n_658),
.Y(n_1117)
);

NOR2xp67_ASAP7_75t_L g1118 ( 
.A(n_1055),
.B(n_37),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_948),
.A2(n_915),
.B(n_910),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1027),
.A2(n_607),
.B(n_609),
.C(n_606),
.Y(n_1120)
);

BUFx12f_ASAP7_75t_L g1121 ( 
.A(n_979),
.Y(n_1121)
);

OAI321xp33_ASAP7_75t_L g1122 ( 
.A1(n_1013),
.A2(n_627),
.A3(n_634),
.B1(n_640),
.B2(n_639),
.C(n_618),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1051),
.A2(n_987),
.B(n_985),
.Y(n_1123)
);

NOR3xp33_ASAP7_75t_L g1124 ( 
.A(n_955),
.B(n_989),
.C(n_951),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1092),
.A2(n_961),
.B(n_1005),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1018),
.A2(n_919),
.B(n_917),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_969),
.A2(n_919),
.B(n_917),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_1003),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_971),
.A2(n_929),
.B(n_924),
.Y(n_1129)
);

OR2x2_ASAP7_75t_L g1130 ( 
.A(n_997),
.B(n_662),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_1027),
.A2(n_1046),
.B(n_981),
.C(n_984),
.Y(n_1131)
);

AO21x1_ASAP7_75t_L g1132 ( 
.A1(n_1007),
.A2(n_645),
.B(n_644),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_982),
.B(n_672),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_957),
.B(n_676),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_1075),
.A2(n_656),
.B(n_660),
.C(n_649),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_1044),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1007),
.A2(n_674),
.B(n_664),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1009),
.A2(n_934),
.B(n_931),
.Y(n_1138)
);

NOR2x1_ASAP7_75t_R g1139 ( 
.A(n_1008),
.B(n_683),
.Y(n_1139)
);

AND2x4_ASAP7_75t_SL g1140 ( 
.A(n_968),
.B(n_617),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_957),
.B(n_684),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1012),
.B(n_617),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1019),
.B(n_637),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_960),
.B(n_669),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_960),
.B(n_675),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_998),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_990),
.A2(n_946),
.B1(n_1026),
.B2(n_993),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_977),
.B(n_679),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1021),
.A2(n_918),
.B(n_682),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_SL g1150 ( 
.A1(n_1042),
.A2(n_638),
.B1(n_652),
.B2(n_637),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1009),
.A2(n_687),
.B(n_681),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_977),
.B(n_689),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_980),
.B(n_692),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_980),
.B(n_693),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_968),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_966),
.B(n_638),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_991),
.B(n_702),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_991),
.B(n_707),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_SL g1159 ( 
.A1(n_1072),
.A2(n_652),
.B1(n_670),
.B2(n_653),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_946),
.A2(n_708),
.B(n_519),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_990),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_952),
.B(n_653),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_968),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_983),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1057),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_995),
.A2(n_527),
.B(n_509),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_990),
.A2(n_677),
.B1(n_686),
.B2(n_670),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_970),
.B(n_527),
.Y(n_1168)
);

INVx5_ASAP7_75t_L g1169 ( 
.A(n_1033),
.Y(n_1169)
);

INVx11_ASAP7_75t_L g1170 ( 
.A(n_1074),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1015),
.B(n_530),
.Y(n_1171)
);

NOR3xp33_ASAP7_75t_L g1172 ( 
.A(n_1039),
.B(n_543),
.C(n_530),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_993),
.B(n_549),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_949),
.A2(n_686),
.B1(n_690),
.B2(n_677),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1017),
.B(n_599),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_964),
.A2(n_663),
.B(n_625),
.C(n_690),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_1015),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1034),
.A2(n_663),
.B(n_625),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1017),
.B(n_520),
.Y(n_1179)
);

AO21x1_ASAP7_75t_L g1180 ( 
.A1(n_1029),
.A2(n_779),
.B(n_586),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_959),
.A2(n_698),
.B(n_336),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1013),
.A2(n_698),
.B(n_337),
.Y(n_1182)
);

CKINVDCx16_ASAP7_75t_R g1183 ( 
.A(n_1073),
.Y(n_1183)
);

AOI221xp5_ASAP7_75t_L g1184 ( 
.A1(n_1058),
.A2(n_698),
.B1(n_39),
.B2(n_37),
.C(n_38),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1023),
.B(n_43),
.Y(n_1185)
);

AND3x2_ASAP7_75t_L g1186 ( 
.A(n_1022),
.B(n_44),
.C(n_45),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1020),
.B(n_47),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1014),
.B(n_47),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_956),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_986),
.A2(n_1011),
.B(n_1029),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1004),
.B(n_1006),
.Y(n_1191)
);

CKINVDCx14_ASAP7_75t_R g1192 ( 
.A(n_988),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1045),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1035),
.B(n_49),
.Y(n_1194)
);

BUFx12f_ASAP7_75t_L g1195 ( 
.A(n_1066),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1026),
.A2(n_53),
.B1(n_49),
.B2(n_50),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_1040),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1062),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_992),
.B(n_60),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_965),
.B(n_62),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_965),
.B(n_63),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1028),
.B(n_66),
.Y(n_1202)
);

NOR3xp33_ASAP7_75t_L g1203 ( 
.A(n_1010),
.B(n_67),
.C(n_68),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1059),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1024),
.A2(n_373),
.B(n_371),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_1050),
.Y(n_1206)
);

BUFx4f_ASAP7_75t_L g1207 ( 
.A(n_1089),
.Y(n_1207)
);

INVxp67_ASAP7_75t_SL g1208 ( 
.A(n_1059),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1056),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1036),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1016),
.A2(n_1038),
.B(n_1037),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1036),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_972),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_973),
.B(n_80),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1069),
.Y(n_1215)
);

OAI321xp33_ASAP7_75t_L g1216 ( 
.A1(n_1085),
.A2(n_81),
.A3(n_82),
.B1(n_83),
.B2(n_84),
.C(n_85),
.Y(n_1216)
);

CKINVDCx10_ASAP7_75t_R g1217 ( 
.A(n_1010),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1030),
.B(n_81),
.Y(n_1218)
);

AND2x6_ASAP7_75t_SL g1219 ( 
.A(n_1043),
.B(n_82),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_975),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1065),
.A2(n_385),
.B(n_384),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1093),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_1025),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1085),
.A2(n_92),
.B1(n_88),
.B2(n_90),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1043),
.A2(n_93),
.B(n_90),
.C(n_92),
.Y(n_1225)
);

AND2x2_ASAP7_75t_SL g1226 ( 
.A(n_994),
.B(n_95),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1070),
.A2(n_396),
.B(n_395),
.Y(n_1227)
);

BUFx8_ASAP7_75t_L g1228 ( 
.A(n_976),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1049),
.B(n_95),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1070),
.A2(n_99),
.B(n_96),
.C(n_98),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_978),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1082),
.A2(n_406),
.B(n_404),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1049),
.B(n_96),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1088),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_L g1235 ( 
.A(n_1001),
.B(n_100),
.C(n_103),
.Y(n_1235)
);

BUFx12f_ASAP7_75t_L g1236 ( 
.A(n_1080),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1082),
.Y(n_1237)
);

AO21x1_ASAP7_75t_L g1238 ( 
.A1(n_1084),
.A2(n_104),
.B(n_105),
.Y(n_1238)
);

BUFx12f_ASAP7_75t_L g1239 ( 
.A(n_1080),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1041),
.A2(n_414),
.B(n_413),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1047),
.B(n_106),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1048),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1084),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1090),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1086),
.A2(n_115),
.B(n_112),
.C(n_113),
.Y(n_1245)
);

CKINVDCx10_ASAP7_75t_R g1246 ( 
.A(n_1064),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1086),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1054),
.A2(n_116),
.B(n_118),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1060),
.A2(n_118),
.B(n_121),
.Y(n_1249)
);

NOR2xp67_ASAP7_75t_L g1250 ( 
.A(n_1053),
.B(n_1061),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_999),
.A2(n_125),
.B(n_126),
.Y(n_1251)
);

AO21x1_ASAP7_75t_L g1252 ( 
.A1(n_1083),
.A2(n_125),
.B(n_126),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1087),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1078),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1094),
.A2(n_1067),
.B(n_1079),
.C(n_1076),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1091),
.A2(n_130),
.B(n_127),
.C(n_129),
.Y(n_1256)
);

AO21x1_ASAP7_75t_L g1257 ( 
.A1(n_1063),
.A2(n_129),
.B(n_130),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1068),
.A2(n_131),
.B(n_133),
.Y(n_1258)
);

CKINVDCx8_ASAP7_75t_R g1259 ( 
.A(n_1090),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1071),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1077),
.A2(n_134),
.B(n_135),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1109),
.B(n_137),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1226),
.B(n_138),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1264)
);

AO31x2_ASAP7_75t_L g1265 ( 
.A1(n_1238),
.A2(n_143),
.A3(n_139),
.B(n_142),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1106),
.B(n_1130),
.Y(n_1266)
);

AOI21xp33_ASAP7_75t_L g1267 ( 
.A1(n_1139),
.A2(n_144),
.B(n_145),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1208),
.B(n_146),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1131),
.A2(n_1190),
.B(n_1255),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1107),
.B(n_147),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1126),
.A2(n_148),
.B(n_150),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1124),
.B(n_152),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1257),
.A2(n_153),
.A3(n_154),
.B(n_155),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_SL g1274 ( 
.A1(n_1147),
.A2(n_153),
.B(n_155),
.Y(n_1274)
);

NAND2x1p5_ASAP7_75t_L g1275 ( 
.A(n_1103),
.B(n_159),
.Y(n_1275)
);

OA22x2_ASAP7_75t_L g1276 ( 
.A1(n_1167),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_1276)
);

O2A1O1Ixp5_ASAP7_75t_L g1277 ( 
.A1(n_1180),
.A2(n_164),
.B(n_165),
.C(n_166),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1146),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1244),
.Y(n_1279)
);

INVx2_ASAP7_75t_SL g1280 ( 
.A(n_1101),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1167),
.B(n_169),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1138),
.A2(n_170),
.B(n_171),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1225),
.A2(n_174),
.B(n_175),
.C(n_176),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1237),
.A2(n_175),
.B(n_176),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1149),
.A2(n_1127),
.B(n_1211),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1105),
.B(n_180),
.Y(n_1286)
);

O2A1O1Ixp5_ASAP7_75t_L g1287 ( 
.A1(n_1181),
.A2(n_181),
.B(n_182),
.C(n_183),
.Y(n_1287)
);

BUFx12f_ASAP7_75t_L g1288 ( 
.A(n_1121),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1165),
.B(n_185),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1243),
.A2(n_186),
.B(n_187),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1128),
.B(n_189),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1247),
.A2(n_189),
.B(n_190),
.Y(n_1292)
);

AND2x6_ASAP7_75t_L g1293 ( 
.A(n_1104),
.B(n_191),
.Y(n_1293)
);

OAI21xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1191),
.A2(n_192),
.B(n_193),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1207),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1195),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1132),
.A2(n_201),
.A3(n_205),
.B(n_206),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1098),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1188),
.A2(n_206),
.B(n_207),
.Y(n_1299)
);

BUFx12f_ASAP7_75t_L g1300 ( 
.A(n_1098),
.Y(n_1300)
);

AO22x2_ASAP7_75t_L g1301 ( 
.A1(n_1210),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1159),
.B(n_210),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1198),
.B(n_211),
.Y(n_1303)
);

OAI22x1_ASAP7_75t_L g1304 ( 
.A1(n_1174),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1188),
.A2(n_212),
.B(n_213),
.Y(n_1305)
);

AO31x2_ASAP7_75t_L g1306 ( 
.A1(n_1210),
.A2(n_215),
.A3(n_216),
.B(n_217),
.Y(n_1306)
);

NOR2x1_ASAP7_75t_SL g1307 ( 
.A(n_1116),
.B(n_1236),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1178),
.A2(n_219),
.B(n_220),
.C(n_221),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1212),
.A2(n_222),
.A3(n_223),
.B(n_224),
.Y(n_1309)
);

A2O1A1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1135),
.A2(n_222),
.B(n_224),
.C(n_225),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1242),
.A2(n_227),
.B(n_228),
.C(n_229),
.Y(n_1311)
);

AO31x2_ASAP7_75t_L g1312 ( 
.A1(n_1212),
.A2(n_228),
.A3(n_230),
.B(n_231),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1148),
.A2(n_1152),
.B(n_1153),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1097),
.A2(n_230),
.B(n_231),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1154),
.A2(n_232),
.B(n_233),
.Y(n_1315)
);

XNOR2xp5_ASAP7_75t_L g1316 ( 
.A(n_1140),
.B(n_233),
.Y(n_1316)
);

INVx5_ASAP7_75t_L g1317 ( 
.A(n_1116),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1194),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1166),
.A2(n_240),
.B(n_241),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1230),
.A2(n_244),
.A3(n_245),
.B(n_246),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1157),
.A2(n_244),
.B(n_245),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1151),
.B(n_246),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1228),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1245),
.A2(n_1252),
.A3(n_1256),
.B(n_1205),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1177),
.B(n_1250),
.Y(n_1325)
);

AO31x2_ASAP7_75t_L g1326 ( 
.A1(n_1196),
.A2(n_248),
.A3(n_250),
.B(n_251),
.Y(n_1326)
);

AO31x2_ASAP7_75t_L g1327 ( 
.A1(n_1196),
.A2(n_255),
.A3(n_256),
.B(n_257),
.Y(n_1327)
);

INVx4_ASAP7_75t_L g1328 ( 
.A(n_1239),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1158),
.A2(n_1145),
.B(n_1144),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1213),
.A2(n_255),
.B(n_256),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1220),
.A2(n_258),
.B(n_259),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1151),
.B(n_258),
.Y(n_1332)
);

INVx6_ASAP7_75t_SL g1333 ( 
.A(n_1171),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1231),
.A2(n_259),
.B(n_260),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1253),
.B(n_261),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1129),
.A2(n_262),
.B(n_263),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1142),
.B(n_263),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1162),
.B(n_264),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1168),
.A2(n_264),
.B(n_265),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1110),
.B(n_265),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1110),
.B(n_266),
.Y(n_1341)
);

CKINVDCx11_ASAP7_75t_R g1342 ( 
.A(n_1099),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1229),
.A2(n_269),
.B(n_270),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1233),
.A2(n_271),
.B(n_272),
.Y(n_1344)
);

INVx3_ASAP7_75t_L g1345 ( 
.A(n_1259),
.Y(n_1345)
);

AO31x2_ASAP7_75t_L g1346 ( 
.A1(n_1187),
.A2(n_273),
.A3(n_274),
.B(n_275),
.Y(n_1346)
);

NOR2xp67_ASAP7_75t_L g1347 ( 
.A(n_1155),
.B(n_276),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1254),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1224),
.A2(n_277),
.A3(n_278),
.B(n_279),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1096),
.B(n_280),
.Y(n_1350)
);

INVx4_ASAP7_75t_L g1351 ( 
.A(n_1215),
.Y(n_1351)
);

AOI221xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1176),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.C(n_283),
.Y(n_1352)
);

INVxp67_ASAP7_75t_L g1353 ( 
.A(n_1111),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1117),
.B(n_287),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1209),
.B(n_288),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1171),
.B(n_288),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1134),
.B(n_290),
.Y(n_1357)
);

AO32x2_ASAP7_75t_L g1358 ( 
.A1(n_1224),
.A2(n_290),
.A3(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_1358)
);

AOI221x1_ASAP7_75t_L g1359 ( 
.A1(n_1137),
.A2(n_1203),
.B1(n_1227),
.B2(n_1232),
.C(n_1235),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1215),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1215),
.Y(n_1361)
);

INVx4_ASAP7_75t_L g1362 ( 
.A(n_1155),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1141),
.B(n_297),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1240),
.A2(n_297),
.B(n_298),
.Y(n_1364)
);

BUFx2_ASAP7_75t_SL g1365 ( 
.A(n_1169),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1202),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1185),
.B(n_1143),
.Y(n_1367)
);

OA22x2_ASAP7_75t_L g1368 ( 
.A1(n_1150),
.A2(n_303),
.B1(n_305),
.B2(n_306),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1120),
.B(n_305),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1214),
.A2(n_307),
.B(n_308),
.Y(n_1370)
);

OAI21xp33_ASAP7_75t_L g1371 ( 
.A1(n_1156),
.A2(n_308),
.B(n_309),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1241),
.A2(n_310),
.B(n_311),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1197),
.B(n_312),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1228),
.Y(n_1374)
);

NOR2xp67_ASAP7_75t_SL g1375 ( 
.A(n_1183),
.B(n_1216),
.Y(n_1375)
);

AOI221x1_ASAP7_75t_L g1376 ( 
.A1(n_1137),
.A2(n_1261),
.B1(n_1258),
.B2(n_1251),
.C(n_1249),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1199),
.A2(n_1119),
.B(n_1115),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1200),
.A2(n_1201),
.B(n_1179),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1184),
.A2(n_1160),
.B(n_1122),
.C(n_1216),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1193),
.A2(n_1234),
.B1(n_1173),
.B2(n_1175),
.Y(n_1380)
);

INVx4_ASAP7_75t_L g1381 ( 
.A(n_1102),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1223),
.B(n_1206),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1218),
.B(n_1172),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1100),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_SL g1385 ( 
.A(n_1136),
.B(n_1163),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1189),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1108),
.A2(n_1260),
.B(n_1133),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1192),
.B(n_1164),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1118),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1186),
.B(n_1219),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1170),
.A2(n_1246),
.B(n_1217),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1392)
);

A2O1A1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1095),
.A2(n_1131),
.B(n_1225),
.C(n_1222),
.Y(n_1393)
);

A2O1A1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1095),
.A2(n_1131),
.B(n_1225),
.C(n_1222),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1105),
.B(n_1027),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1107),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1125),
.A2(n_962),
.B(n_1123),
.Y(n_1398)
);

AO32x2_ASAP7_75t_L g1399 ( 
.A1(n_1210),
.A2(n_1212),
.A3(n_1147),
.B1(n_1196),
.B2(n_1224),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1112),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1125),
.A2(n_962),
.B(n_1123),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1109),
.B(n_997),
.Y(n_1403)
);

AO31x2_ASAP7_75t_L g1404 ( 
.A1(n_1238),
.A2(n_1257),
.A3(n_1180),
.B(n_1161),
.Y(n_1404)
);

AO31x2_ASAP7_75t_L g1405 ( 
.A1(n_1238),
.A2(n_1257),
.A3(n_1180),
.B(n_1161),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1112),
.Y(n_1406)
);

OA22x2_ASAP7_75t_L g1407 ( 
.A1(n_1167),
.A2(n_1150),
.B1(n_1140),
.B2(n_1174),
.Y(n_1407)
);

AO22x2_ASAP7_75t_L g1408 ( 
.A1(n_1167),
.A2(n_1147),
.B1(n_1106),
.B2(n_1210),
.Y(n_1408)
);

A2O1A1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1095),
.A2(n_1131),
.B(n_1225),
.C(n_1222),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1121),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1128),
.B(n_1103),
.Y(n_1411)
);

OA22x2_ASAP7_75t_L g1412 ( 
.A1(n_1167),
.A2(n_1150),
.B1(n_1140),
.B2(n_1174),
.Y(n_1412)
);

OAI21xp33_ASAP7_75t_L g1413 ( 
.A1(n_1113),
.A2(n_820),
.B(n_1105),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1125),
.A2(n_962),
.B(n_1123),
.Y(n_1414)
);

AO32x2_ASAP7_75t_L g1415 ( 
.A1(n_1210),
.A2(n_1212),
.A3(n_1147),
.B1(n_1196),
.B2(n_1224),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1105),
.B(n_1027),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1109),
.B(n_997),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_SL g1418 ( 
.A1(n_1182),
.A2(n_1248),
.B(n_1147),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_SL g1419 ( 
.A(n_1226),
.B(n_1147),
.Y(n_1419)
);

AO31x2_ASAP7_75t_L g1420 ( 
.A1(n_1238),
.A2(n_1257),
.A3(n_1180),
.B(n_1161),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1121),
.Y(n_1422)
);

INVx4_ASAP7_75t_L g1423 ( 
.A(n_1101),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1244),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1125),
.A2(n_962),
.B(n_1123),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1103),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1125),
.A2(n_962),
.B(n_1123),
.Y(n_1428)
);

OAI22x1_ASAP7_75t_L g1429 ( 
.A1(n_1174),
.A2(n_748),
.B1(n_753),
.B2(n_750),
.Y(n_1429)
);

INVx2_ASAP7_75t_SL g1430 ( 
.A(n_1101),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1125),
.A2(n_962),
.B(n_1123),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1125),
.A2(n_962),
.B(n_1123),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1095),
.A2(n_1131),
.B(n_1225),
.C(n_1222),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1109),
.B(n_997),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1109),
.B(n_997),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1161),
.A2(n_1208),
.B1(n_1147),
.B2(n_826),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1439)
);

A2O1A1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1095),
.A2(n_1131),
.B(n_1225),
.C(n_1222),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1109),
.B(n_997),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1121),
.Y(n_1443)
);

AOI21xp33_ASAP7_75t_L g1444 ( 
.A1(n_1139),
.A2(n_1113),
.B(n_932),
.Y(n_1444)
);

NAND3x1_ASAP7_75t_L g1445 ( 
.A(n_1124),
.B(n_1174),
.C(n_777),
.Y(n_1445)
);

OAI22x1_ASAP7_75t_L g1446 ( 
.A1(n_1174),
.A2(n_748),
.B1(n_753),
.B2(n_750),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1109),
.B(n_997),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1448)
);

AO21x1_ASAP7_75t_L g1449 ( 
.A1(n_1182),
.A2(n_1114),
.B(n_1221),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_SL g1450 ( 
.A1(n_1182),
.A2(n_1248),
.B(n_1147),
.Y(n_1450)
);

OR2x6_ASAP7_75t_L g1451 ( 
.A(n_1121),
.B(n_1155),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1109),
.B(n_997),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_SL g1455 ( 
.A(n_1226),
.B(n_1147),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1109),
.B(n_997),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1101),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1112),
.Y(n_1459)
);

A2O1A1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1095),
.A2(n_1131),
.B(n_1225),
.C(n_1222),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1121),
.Y(n_1461)
);

NAND2x1p5_ASAP7_75t_L g1462 ( 
.A(n_1103),
.B(n_1104),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1109),
.B(n_997),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1161),
.A2(n_1208),
.B1(n_1147),
.B2(n_826),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1112),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1161),
.A2(n_1208),
.B1(n_1147),
.B2(n_826),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1125),
.A2(n_962),
.B(n_1123),
.Y(n_1468)
);

OAI21xp33_ASAP7_75t_L g1469 ( 
.A1(n_1113),
.A2(n_820),
.B(n_1105),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1095),
.B(n_1204),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1109),
.B(n_997),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1107),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1397),
.B(n_1472),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1398),
.A2(n_1414),
.B(n_1401),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1288),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1266),
.B(n_1403),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1417),
.B(n_1436),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1437),
.B(n_1441),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1398),
.A2(n_1414),
.B(n_1401),
.Y(n_1479)
);

A2O1A1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1313),
.A2(n_1329),
.B(n_1363),
.C(n_1357),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1278),
.Y(n_1481)
);

NAND3xp33_ASAP7_75t_L g1482 ( 
.A(n_1352),
.B(n_1277),
.C(n_1367),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1317),
.B(n_1307),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1400),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1379),
.A2(n_1394),
.B(n_1393),
.Y(n_1485)
);

AO31x2_ASAP7_75t_L g1486 ( 
.A1(n_1425),
.A2(n_1431),
.A3(n_1432),
.B(n_1428),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1406),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1317),
.B(n_1351),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1348),
.Y(n_1489)
);

AND2x2_ASAP7_75t_SL g1490 ( 
.A(n_1374),
.B(n_1281),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1447),
.B(n_1452),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1317),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1408),
.A2(n_1419),
.B1(n_1455),
.B2(n_1438),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1456),
.B(n_1463),
.Y(n_1494)
);

OAI21xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1263),
.A2(n_1455),
.B(n_1419),
.Y(n_1495)
);

OAI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1407),
.A2(n_1412),
.B1(n_1276),
.B2(n_1368),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1342),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1471),
.B(n_1302),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1300),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1413),
.B(n_1469),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1333),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1459),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1466),
.Y(n_1503)
);

A2O1A1Ixp33_ASAP7_75t_L g1504 ( 
.A1(n_1357),
.A2(n_1394),
.B(n_1409),
.C(n_1393),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1408),
.A2(n_1407),
.B1(n_1412),
.B2(n_1272),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1367),
.B(n_1366),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1396),
.B(n_1416),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1468),
.A2(n_1377),
.B(n_1285),
.Y(n_1508)
);

O2A1O1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1433),
.A2(n_1440),
.B(n_1460),
.C(n_1310),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1443),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_1361),
.Y(n_1511)
);

INVx8_ASAP7_75t_L g1512 ( 
.A(n_1293),
.Y(n_1512)
);

AOI21xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1316),
.A2(n_1384),
.B(n_1368),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1386),
.B(n_1296),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1262),
.B(n_1270),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1411),
.B(n_1362),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1335),
.B(n_1286),
.Y(n_1517)
);

NOR2xp67_ASAP7_75t_L g1518 ( 
.A(n_1423),
.B(n_1328),
.Y(n_1518)
);

INVx5_ASAP7_75t_L g1519 ( 
.A(n_1293),
.Y(n_1519)
);

INVx6_ASAP7_75t_L g1520 ( 
.A(n_1423),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1328),
.Y(n_1521)
);

OAI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1440),
.A2(n_1460),
.B(n_1269),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_SL g1523 ( 
.A1(n_1408),
.A2(n_1301),
.B1(n_1276),
.B2(n_1293),
.Y(n_1523)
);

OAI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1465),
.A2(n_1467),
.B1(n_1322),
.B2(n_1332),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1264),
.A2(n_1392),
.B1(n_1402),
.B2(n_1395),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1353),
.B(n_1291),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1286),
.B(n_1353),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1410),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1333),
.Y(n_1529)
);

OAI221xp5_ASAP7_75t_L g1530 ( 
.A1(n_1383),
.A2(n_1283),
.B1(n_1444),
.B2(n_1369),
.C(n_1318),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1360),
.B(n_1356),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_SL g1532 ( 
.A(n_1375),
.B(n_1293),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1289),
.B(n_1303),
.Y(n_1533)
);

OAI22x1_ASAP7_75t_L g1534 ( 
.A1(n_1291),
.A2(n_1381),
.B1(n_1323),
.B2(n_1275),
.Y(n_1534)
);

INVx6_ASAP7_75t_L g1535 ( 
.A(n_1362),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1289),
.B(n_1382),
.Y(n_1536)
);

A2O1A1Ixp33_ASAP7_75t_L g1537 ( 
.A1(n_1350),
.A2(n_1470),
.B(n_1464),
.C(n_1457),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1422),
.Y(n_1538)
);

AND2x2_ASAP7_75t_SL g1539 ( 
.A(n_1381),
.B(n_1461),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1451),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1421),
.A2(n_1426),
.B1(n_1454),
.B2(n_1453),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1303),
.B(n_1355),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_SL g1543 ( 
.A1(n_1301),
.A2(n_1290),
.B1(n_1284),
.B2(n_1292),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1434),
.A2(n_1439),
.B1(n_1448),
.B2(n_1435),
.Y(n_1544)
);

OR2x6_ASAP7_75t_L g1545 ( 
.A(n_1451),
.B(n_1280),
.Y(n_1545)
);

AO31x2_ASAP7_75t_L g1546 ( 
.A1(n_1359),
.A2(n_1376),
.A3(n_1380),
.B(n_1271),
.Y(n_1546)
);

OAI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1442),
.A2(n_1378),
.B(n_1287),
.Y(n_1547)
);

INVx5_ASAP7_75t_L g1548 ( 
.A(n_1279),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1346),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1338),
.B(n_1429),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1430),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1346),
.Y(n_1552)
);

OAI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1304),
.A2(n_1334),
.B1(n_1330),
.B2(n_1331),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1301),
.A2(n_1337),
.B1(n_1318),
.B2(n_1371),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1346),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1268),
.Y(n_1556)
);

INVx4_ASAP7_75t_SL g1557 ( 
.A(n_1306),
.Y(n_1557)
);

NOR2x1_ASAP7_75t_R g1558 ( 
.A(n_1298),
.B(n_1458),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1462),
.Y(n_1559)
);

NOR2xp67_ASAP7_75t_L g1560 ( 
.A(n_1446),
.B(n_1390),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1396),
.B(n_1416),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1462),
.Y(n_1562)
);

BUFx4f_ASAP7_75t_SL g1563 ( 
.A(n_1345),
.Y(n_1563)
);

INVx4_ASAP7_75t_L g1564 ( 
.A(n_1345),
.Y(n_1564)
);

OR2x6_ASAP7_75t_L g1565 ( 
.A(n_1365),
.B(n_1274),
.Y(n_1565)
);

OAI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1295),
.A2(n_1314),
.B1(n_1347),
.B2(n_1282),
.Y(n_1566)
);

O2A1O1Ixp33_ASAP7_75t_L g1567 ( 
.A1(n_1308),
.A2(n_1311),
.B(n_1294),
.C(n_1341),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1388),
.B(n_1340),
.Y(n_1568)
);

OAI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1336),
.A2(n_1364),
.B(n_1445),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1349),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1354),
.B(n_1373),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1349),
.Y(n_1572)
);

AOI222xp33_ASAP7_75t_L g1573 ( 
.A1(n_1385),
.A2(n_1373),
.B1(n_1391),
.B2(n_1325),
.C1(n_1319),
.C2(n_1387),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1427),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1267),
.B(n_1325),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1297),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1339),
.A2(n_1315),
.B1(n_1321),
.B2(n_1343),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1343),
.A2(n_1344),
.B1(n_1305),
.B2(n_1299),
.Y(n_1578)
);

CKINVDCx11_ASAP7_75t_R g1579 ( 
.A(n_1389),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1297),
.Y(n_1580)
);

AO31x2_ASAP7_75t_L g1581 ( 
.A1(n_1299),
.A2(n_1305),
.A3(n_1370),
.B(n_1372),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1326),
.Y(n_1582)
);

OAI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1404),
.A2(n_1405),
.B(n_1420),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1399),
.A2(n_1415),
.B1(n_1358),
.B2(n_1424),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1424),
.B(n_1399),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1415),
.A2(n_1358),
.B1(n_1327),
.B2(n_1326),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1404),
.A2(n_1420),
.B(n_1405),
.Y(n_1587)
);

AND2x2_ASAP7_75t_SL g1588 ( 
.A(n_1415),
.B(n_1358),
.Y(n_1588)
);

OAI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1404),
.A2(n_1420),
.B(n_1405),
.Y(n_1589)
);

OAI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1358),
.A2(n_1312),
.B1(n_1309),
.B2(n_1306),
.C(n_1327),
.Y(n_1590)
);

AO32x2_ASAP7_75t_L g1591 ( 
.A1(n_1306),
.A2(n_1309),
.A3(n_1312),
.B1(n_1420),
.B2(n_1405),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1404),
.A2(n_1324),
.B(n_1273),
.Y(n_1592)
);

AO32x2_ASAP7_75t_L g1593 ( 
.A1(n_1306),
.A2(n_1309),
.A3(n_1312),
.B1(n_1327),
.B2(n_1326),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1324),
.A2(n_1265),
.B(n_1320),
.Y(n_1594)
);

INVx4_ASAP7_75t_L g1595 ( 
.A(n_1327),
.Y(n_1595)
);

AO21x2_ASAP7_75t_L g1596 ( 
.A1(n_1320),
.A2(n_1309),
.B(n_1312),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_SL g1597 ( 
.A1(n_1408),
.A2(n_1167),
.B1(n_1412),
.B2(n_1407),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1288),
.Y(n_1598)
);

OAI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1281),
.A2(n_1412),
.B1(n_1407),
.B2(n_1161),
.Y(n_1599)
);

CKINVDCx20_ASAP7_75t_R g1600 ( 
.A(n_1443),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1348),
.Y(n_1601)
);

AO221x2_ASAP7_75t_L g1602 ( 
.A1(n_1304),
.A2(n_1167),
.B1(n_1150),
.B2(n_955),
.C(n_761),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1266),
.B(n_1413),
.Y(n_1603)
);

OR2x6_ASAP7_75t_L g1604 ( 
.A(n_1300),
.B(n_1121),
.Y(n_1604)
);

AOI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1407),
.A2(n_786),
.B1(n_1167),
.B2(n_1113),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1288),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1408),
.A2(n_1412),
.B1(n_1407),
.B2(n_1419),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1266),
.B(n_1413),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1397),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1398),
.A2(n_1414),
.B(n_1401),
.Y(n_1610)
);

OR2x6_ASAP7_75t_L g1611 ( 
.A(n_1300),
.B(n_1121),
.Y(n_1611)
);

AO21x2_ASAP7_75t_L g1612 ( 
.A1(n_1418),
.A2(n_1450),
.B(n_1449),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_SL g1613 ( 
.A1(n_1408),
.A2(n_1167),
.B1(n_1412),
.B2(n_1407),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_1443),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1379),
.A2(n_1329),
.B(n_1313),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1408),
.A2(n_1412),
.B1(n_1407),
.B2(n_1419),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1317),
.B(n_1307),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1379),
.A2(n_1329),
.B(n_1313),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1266),
.B(n_1413),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1408),
.A2(n_1412),
.B1(n_1407),
.B2(n_1419),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1288),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_SL g1622 ( 
.A1(n_1408),
.A2(n_1167),
.B1(n_1412),
.B2(n_1407),
.Y(n_1622)
);

O2A1O1Ixp33_ASAP7_75t_L g1623 ( 
.A1(n_1393),
.A2(n_1409),
.B(n_1433),
.C(n_1394),
.Y(n_1623)
);

BUFx3_ASAP7_75t_L g1624 ( 
.A(n_1288),
.Y(n_1624)
);

INVx6_ASAP7_75t_L g1625 ( 
.A(n_1317),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1408),
.A2(n_1167),
.B1(n_1412),
.B2(n_1407),
.Y(n_1626)
);

OAI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1605),
.A2(n_1512),
.B1(n_1476),
.B2(n_1532),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1481),
.Y(n_1628)
);

OA21x2_ASAP7_75t_L g1629 ( 
.A1(n_1508),
.A2(n_1610),
.B(n_1474),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1484),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1483),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1487),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1502),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1477),
.B(n_1494),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1522),
.B(n_1607),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1479),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_SL g1637 ( 
.A1(n_1490),
.A2(n_1602),
.B1(n_1512),
.B2(n_1532),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1597),
.A2(n_1613),
.B1(n_1626),
.B2(n_1622),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1522),
.B(n_1607),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1503),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1478),
.B(n_1491),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1483),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1507),
.B(n_1561),
.Y(n_1643)
);

NOR2x1_ASAP7_75t_SL g1644 ( 
.A(n_1519),
.B(n_1565),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_SL g1645 ( 
.A1(n_1602),
.A2(n_1519),
.B1(n_1507),
.B2(n_1603),
.Y(n_1645)
);

BUFx2_ASAP7_75t_SL g1646 ( 
.A(n_1518),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1473),
.Y(n_1647)
);

INVx5_ASAP7_75t_L g1648 ( 
.A(n_1519),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1506),
.B(n_1498),
.Y(n_1649)
);

INVx1_ASAP7_75t_SL g1650 ( 
.A(n_1600),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1609),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1548),
.B(n_1488),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1609),
.Y(n_1653)
);

AO21x2_ASAP7_75t_L g1654 ( 
.A1(n_1594),
.A2(n_1618),
.B(n_1615),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1489),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1486),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1486),
.Y(n_1657)
);

INVx4_ASAP7_75t_L g1658 ( 
.A(n_1617),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1617),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1604),
.Y(n_1660)
);

OAI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1482),
.A2(n_1480),
.B(n_1537),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1604),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1601),
.Y(n_1663)
);

AO21x2_ASAP7_75t_L g1664 ( 
.A1(n_1594),
.A2(n_1618),
.B(n_1615),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1506),
.B(n_1603),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1504),
.A2(n_1500),
.B(n_1567),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1597),
.A2(n_1613),
.B1(n_1626),
.B2(n_1622),
.Y(n_1667)
);

OAI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1500),
.A2(n_1567),
.B(n_1530),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1543),
.B(n_1566),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1616),
.B(n_1620),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1492),
.Y(n_1671)
);

INVx2_ASAP7_75t_SL g1672 ( 
.A(n_1625),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1525),
.A2(n_1544),
.B(n_1547),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1625),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1608),
.B(n_1619),
.Y(n_1675)
);

OAI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1513),
.A2(n_1599),
.B1(n_1565),
.B2(n_1545),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1548),
.B(n_1565),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1616),
.B(n_1620),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1492),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1526),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1625),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1614),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1534),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_R g1684 ( 
.A(n_1621),
.B(n_1497),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1608),
.B(n_1619),
.Y(n_1685)
);

OAI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1599),
.A2(n_1545),
.B1(n_1604),
.B2(n_1611),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1531),
.Y(n_1687)
);

BUFx12f_ASAP7_75t_L g1688 ( 
.A(n_1611),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1496),
.A2(n_1530),
.B1(n_1505),
.B2(n_1543),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1516),
.Y(n_1690)
);

OA21x2_ASAP7_75t_L g1691 ( 
.A1(n_1583),
.A2(n_1592),
.B(n_1589),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1511),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1611),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1533),
.B(n_1517),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1485),
.B(n_1505),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1549),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1527),
.B(n_1515),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1535),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1485),
.B(n_1588),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1541),
.B(n_1556),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1535),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1552),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1555),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1536),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1568),
.B(n_1571),
.Y(n_1705)
);

INVx2_ASAP7_75t_SL g1706 ( 
.A(n_1535),
.Y(n_1706)
);

OA21x2_ASAP7_75t_L g1707 ( 
.A1(n_1583),
.A2(n_1587),
.B(n_1547),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1573),
.A2(n_1496),
.B1(n_1575),
.B2(n_1544),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1528),
.Y(n_1709)
);

BUFx2_ASAP7_75t_L g1710 ( 
.A(n_1545),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_SL g1711 ( 
.A(n_1624),
.Y(n_1711)
);

NOR2x1_ASAP7_75t_SL g1712 ( 
.A(n_1559),
.B(n_1562),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1523),
.B(n_1591),
.Y(n_1713)
);

INVx4_ASAP7_75t_L g1714 ( 
.A(n_1648),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1699),
.B(n_1576),
.Y(n_1715)
);

INVx4_ASAP7_75t_L g1716 ( 
.A(n_1648),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1636),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1628),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1630),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1632),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1633),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1713),
.B(n_1580),
.Y(n_1722)
);

BUFx2_ASAP7_75t_SL g1723 ( 
.A(n_1711),
.Y(n_1723)
);

INVxp67_ASAP7_75t_L g1724 ( 
.A(n_1634),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1635),
.B(n_1639),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1640),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1692),
.Y(n_1727)
);

AND2x4_ASAP7_75t_SL g1728 ( 
.A(n_1658),
.B(n_1652),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_SL g1729 ( 
.A1(n_1638),
.A2(n_1644),
.B1(n_1658),
.B2(n_1688),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1677),
.B(n_1557),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1704),
.B(n_1573),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1677),
.B(n_1557),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1686),
.A2(n_1523),
.B1(n_1493),
.B2(n_1524),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1695),
.B(n_1595),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1677),
.B(n_1557),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1695),
.B(n_1595),
.Y(n_1736)
);

BUFx3_ASAP7_75t_L g1737 ( 
.A(n_1642),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_1648),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1643),
.B(n_1623),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1651),
.Y(n_1740)
);

NOR2x1p5_ASAP7_75t_L g1741 ( 
.A(n_1688),
.B(n_1540),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1643),
.B(n_1623),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1671),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1700),
.B(n_1570),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1700),
.B(n_1572),
.Y(n_1745)
);

INVx4_ASAP7_75t_L g1746 ( 
.A(n_1648),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1670),
.B(n_1582),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1653),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1670),
.B(n_1585),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1678),
.B(n_1591),
.Y(n_1750)
);

AND2x4_ASAP7_75t_SL g1751 ( 
.A(n_1658),
.B(n_1564),
.Y(n_1751)
);

INVxp67_ASAP7_75t_L g1752 ( 
.A(n_1634),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1654),
.B(n_1596),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1654),
.B(n_1596),
.Y(n_1754)
);

AND2x4_ASAP7_75t_SL g1755 ( 
.A(n_1652),
.B(n_1564),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1654),
.B(n_1584),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1665),
.B(n_1511),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1705),
.B(n_1509),
.Y(n_1758)
);

BUFx3_ASAP7_75t_L g1759 ( 
.A(n_1631),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1705),
.B(n_1509),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1664),
.B(n_1584),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1666),
.B(n_1612),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1668),
.B(n_1612),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1669),
.B(n_1593),
.Y(n_1764)
);

OAI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1708),
.A2(n_1660),
.B1(n_1693),
.B2(n_1662),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1669),
.B(n_1586),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1687),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1696),
.B(n_1586),
.Y(n_1768)
);

NOR2x1p5_ASAP7_75t_L g1769 ( 
.A(n_1660),
.B(n_1499),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1641),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1702),
.B(n_1546),
.Y(n_1771)
);

CKINVDCx8_ASAP7_75t_R g1772 ( 
.A(n_1646),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1703),
.B(n_1546),
.Y(n_1773)
);

OAI222xp33_ASAP7_75t_L g1774 ( 
.A1(n_1637),
.A2(n_1645),
.B1(n_1689),
.B2(n_1676),
.C1(n_1667),
.C2(n_1627),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1647),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1675),
.B(n_1685),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1661),
.B(n_1569),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1656),
.B(n_1581),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1659),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1734),
.B(n_1707),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1734),
.B(n_1707),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1771),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1771),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1736),
.B(n_1707),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_1743),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1717),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1773),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1730),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1724),
.B(n_1649),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1773),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1743),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1736),
.B(n_1657),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1722),
.B(n_1715),
.Y(n_1793)
);

CKINVDCx11_ASAP7_75t_R g1794 ( 
.A(n_1772),
.Y(n_1794)
);

INVx1_ASAP7_75t_SL g1795 ( 
.A(n_1728),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1768),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1768),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1752),
.B(n_1725),
.Y(n_1798)
);

INVxp67_ASAP7_75t_L g1799 ( 
.A(n_1740),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1748),
.Y(n_1800)
);

BUFx2_ASAP7_75t_SL g1801 ( 
.A(n_1772),
.Y(n_1801)
);

OR2x6_ASAP7_75t_L g1802 ( 
.A(n_1732),
.B(n_1673),
.Y(n_1802)
);

BUFx3_ASAP7_75t_L g1803 ( 
.A(n_1728),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1778),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1723),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1779),
.Y(n_1806)
);

INVxp67_ASAP7_75t_L g1807 ( 
.A(n_1775),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1733),
.A2(n_1667),
.B1(n_1554),
.B2(n_1694),
.Y(n_1808)
);

INVx5_ASAP7_75t_L g1809 ( 
.A(n_1738),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1750),
.B(n_1691),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1750),
.B(n_1691),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1767),
.B(n_1697),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1749),
.B(n_1629),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1755),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1727),
.Y(n_1815)
);

NOR2x1_ASAP7_75t_L g1816 ( 
.A(n_1741),
.B(n_1679),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1744),
.B(n_1691),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1770),
.B(n_1650),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1744),
.B(n_1629),
.Y(n_1819)
);

INVx4_ASAP7_75t_L g1820 ( 
.A(n_1714),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1759),
.Y(n_1821)
);

INVx2_ASAP7_75t_SL g1822 ( 
.A(n_1759),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1737),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1745),
.B(n_1763),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1780),
.B(n_1756),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1786),
.Y(n_1826)
);

AND2x4_ASAP7_75t_SL g1827 ( 
.A(n_1820),
.B(n_1735),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1785),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1804),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1813),
.B(n_1763),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1804),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1780),
.B(n_1756),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1793),
.B(n_1749),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1813),
.B(n_1766),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1781),
.B(n_1761),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1820),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1793),
.B(n_1747),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1781),
.B(n_1761),
.Y(n_1838)
);

INVx3_ASAP7_75t_L g1839 ( 
.A(n_1820),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1784),
.B(n_1753),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1791),
.Y(n_1841)
);

BUFx3_ASAP7_75t_L g1842 ( 
.A(n_1803),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_SL g1843 ( 
.A(n_1801),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1784),
.B(n_1753),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1796),
.B(n_1766),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1796),
.B(n_1797),
.Y(n_1846)
);

NOR2xp67_ASAP7_75t_L g1847 ( 
.A(n_1809),
.B(n_1714),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1824),
.B(n_1731),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1805),
.B(n_1662),
.Y(n_1849)
);

AND2x4_ASAP7_75t_L g1850 ( 
.A(n_1802),
.B(n_1754),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1810),
.B(n_1754),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1797),
.B(n_1762),
.Y(n_1852)
);

INVx4_ASAP7_75t_L g1853 ( 
.A(n_1803),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1782),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1798),
.B(n_1762),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1782),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1783),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1810),
.B(n_1764),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1787),
.Y(n_1859)
);

NAND2x1p5_ASAP7_75t_L g1860 ( 
.A(n_1816),
.B(n_1714),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1811),
.B(n_1764),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1811),
.B(n_1819),
.Y(n_1862)
);

BUFx2_ASAP7_75t_L g1863 ( 
.A(n_1785),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1854),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1848),
.B(n_1800),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1834),
.B(n_1787),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1834),
.B(n_1790),
.Y(n_1867)
);

INVx1_ASAP7_75t_SL g1868 ( 
.A(n_1843),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1854),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1845),
.B(n_1815),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1856),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1862),
.B(n_1819),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1856),
.Y(n_1873)
);

HB1xp67_ASAP7_75t_L g1874 ( 
.A(n_1841),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1862),
.B(n_1817),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1851),
.B(n_1817),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1826),
.Y(n_1877)
);

INVxp67_ASAP7_75t_L g1878 ( 
.A(n_1863),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1857),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1857),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1830),
.B(n_1851),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1859),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1859),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1863),
.Y(n_1884)
);

OR2x6_ASAP7_75t_L g1885 ( 
.A(n_1853),
.B(n_1802),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1858),
.B(n_1802),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1845),
.B(n_1806),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1829),
.Y(n_1888)
);

INVxp67_ASAP7_75t_L g1889 ( 
.A(n_1828),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1858),
.B(n_1861),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1861),
.B(n_1802),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1849),
.B(n_1807),
.Y(n_1892)
);

OR3x2_ASAP7_75t_L g1893 ( 
.A(n_1827),
.B(n_1794),
.C(n_1801),
.Y(n_1893)
);

BUFx2_ASAP7_75t_L g1894 ( 
.A(n_1853),
.Y(n_1894)
);

NAND3x1_ASAP7_75t_L g1895 ( 
.A(n_1836),
.B(n_1788),
.C(n_1818),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1830),
.B(n_1790),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1840),
.B(n_1792),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1840),
.B(n_1792),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1890),
.B(n_1872),
.Y(n_1899)
);

OAI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1894),
.A2(n_1853),
.B1(n_1836),
.B2(n_1839),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1881),
.B(n_1866),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1866),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1874),
.B(n_1799),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1890),
.B(n_1844),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_SL g1905 ( 
.A(n_1868),
.B(n_1853),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1877),
.Y(n_1906)
);

OR2x6_ASAP7_75t_L g1907 ( 
.A(n_1894),
.B(n_1836),
.Y(n_1907)
);

INVx2_ASAP7_75t_SL g1908 ( 
.A(n_1884),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1881),
.B(n_1855),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1876),
.B(n_1844),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1867),
.B(n_1855),
.Y(n_1911)
);

OAI32xp33_ASAP7_75t_L g1912 ( 
.A1(n_1889),
.A2(n_1836),
.A3(n_1839),
.B1(n_1842),
.B2(n_1860),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1867),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1877),
.Y(n_1914)
);

INVxp67_ASAP7_75t_SL g1915 ( 
.A(n_1895),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1896),
.Y(n_1916)
);

NAND3x2_ASAP7_75t_L g1917 ( 
.A(n_1886),
.B(n_1850),
.C(n_1852),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1876),
.B(n_1825),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1872),
.B(n_1825),
.Y(n_1919)
);

INVx1_ASAP7_75t_SL g1920 ( 
.A(n_1870),
.Y(n_1920)
);

OAI21xp33_ASAP7_75t_L g1921 ( 
.A1(n_1886),
.A2(n_1850),
.B(n_1846),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1896),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1875),
.B(n_1832),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1864),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1864),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1875),
.B(n_1832),
.Y(n_1926)
);

OAI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1895),
.A2(n_1847),
.B(n_1774),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1887),
.B(n_1835),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1897),
.B(n_1835),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1865),
.B(n_1837),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1869),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1869),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1871),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1878),
.B(n_1839),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1871),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1873),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1905),
.B(n_1839),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1911),
.Y(n_1938)
);

INVxp67_ASAP7_75t_L g1939 ( 
.A(n_1903),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1901),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1900),
.A2(n_1827),
.B(n_1885),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1920),
.B(n_1897),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1906),
.Y(n_1943)
);

OAI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1917),
.A2(n_1893),
.B1(n_1827),
.B2(n_1885),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1909),
.Y(n_1945)
);

OAI32xp33_ASAP7_75t_L g1946 ( 
.A1(n_1927),
.A2(n_1842),
.A3(n_1814),
.B1(n_1860),
.B2(n_1795),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1902),
.B(n_1898),
.Y(n_1947)
);

OAI21xp33_ASAP7_75t_L g1948 ( 
.A1(n_1915),
.A2(n_1891),
.B(n_1892),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1924),
.Y(n_1949)
);

OAI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1907),
.A2(n_1893),
.B1(n_1885),
.B2(n_1842),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1925),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1931),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1913),
.B(n_1898),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1906),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1907),
.A2(n_1885),
.B1(n_1891),
.B2(n_1860),
.Y(n_1955)
);

OAI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1907),
.A2(n_1885),
.B1(n_1847),
.B2(n_1833),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1916),
.B(n_1831),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1914),
.Y(n_1958)
);

INVx3_ASAP7_75t_L g1959 ( 
.A(n_1908),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1932),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1949),
.B(n_1933),
.Y(n_1961)
);

OAI221xp5_ASAP7_75t_L g1962 ( 
.A1(n_1948),
.A2(n_1915),
.B1(n_1921),
.B2(n_1934),
.C(n_1908),
.Y(n_1962)
);

AOI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1939),
.A2(n_1903),
.B1(n_1934),
.B2(n_1850),
.Y(n_1963)
);

NOR3xp33_ASAP7_75t_L g1964 ( 
.A(n_1946),
.B(n_1950),
.C(n_1944),
.Y(n_1964)
);

OAI21xp33_ASAP7_75t_SL g1965 ( 
.A1(n_1937),
.A2(n_1899),
.B(n_1926),
.Y(n_1965)
);

NOR2x1_ASAP7_75t_L g1966 ( 
.A(n_1937),
.B(n_1959),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1939),
.A2(n_1850),
.B1(n_1900),
.B2(n_1729),
.Y(n_1967)
);

INVxp33_ASAP7_75t_L g1968 ( 
.A(n_1941),
.Y(n_1968)
);

OAI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1959),
.A2(n_1956),
.B(n_1955),
.Y(n_1969)
);

NOR2xp33_ASAP7_75t_L g1970 ( 
.A(n_1945),
.B(n_1938),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1942),
.A2(n_1912),
.B(n_1693),
.Y(n_1971)
);

AOI211x1_ASAP7_75t_L g1972 ( 
.A1(n_1940),
.A2(n_1904),
.B(n_1928),
.C(n_1910),
.Y(n_1972)
);

AOI311xp33_ASAP7_75t_L g1973 ( 
.A1(n_1960),
.A2(n_1922),
.A3(n_1765),
.B(n_1789),
.C(n_1935),
.Y(n_1973)
);

INVxp67_ASAP7_75t_L g1974 ( 
.A(n_1957),
.Y(n_1974)
);

HB1xp67_ASAP7_75t_L g1975 ( 
.A(n_1951),
.Y(n_1975)
);

NOR4xp75_ASAP7_75t_SL g1976 ( 
.A(n_1947),
.B(n_1929),
.C(n_1919),
.D(n_1918),
.Y(n_1976)
);

NAND3xp33_ASAP7_75t_L g1977 ( 
.A(n_1952),
.B(n_1683),
.C(n_1709),
.Y(n_1977)
);

OAI211xp5_ASAP7_75t_L g1978 ( 
.A1(n_1953),
.A2(n_1682),
.B(n_1684),
.C(n_1808),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1943),
.B(n_1926),
.Y(n_1979)
);

OAI32xp33_ASAP7_75t_L g1980 ( 
.A1(n_1943),
.A2(n_1930),
.A3(n_1821),
.B1(n_1923),
.B2(n_1823),
.Y(n_1980)
);

AOI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1954),
.A2(n_1539),
.B(n_1751),
.Y(n_1981)
);

AOI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1954),
.A2(n_1751),
.B(n_1828),
.Y(n_1982)
);

AOI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1958),
.A2(n_1936),
.B1(n_1879),
.B2(n_1880),
.Y(n_1983)
);

NOR2x1_ASAP7_75t_L g1984 ( 
.A(n_1958),
.B(n_1769),
.Y(n_1984)
);

OAI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1937),
.A2(n_1495),
.B(n_1822),
.Y(n_1985)
);

NAND4xp25_ASAP7_75t_L g1986 ( 
.A(n_1948),
.B(n_1510),
.C(n_1560),
.D(n_1758),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1937),
.A2(n_1755),
.B(n_1822),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1974),
.B(n_1838),
.Y(n_1988)
);

O2A1O1Ixp5_ASAP7_75t_L g1989 ( 
.A1(n_1968),
.A2(n_1746),
.B(n_1716),
.C(n_1757),
.Y(n_1989)
);

NOR2xp33_ASAP7_75t_L g1990 ( 
.A(n_1965),
.B(n_1475),
.Y(n_1990)
);

AOI221x1_ASAP7_75t_L g1991 ( 
.A1(n_1964),
.A2(n_1879),
.B1(n_1882),
.B2(n_1880),
.C(n_1873),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1961),
.B(n_1846),
.Y(n_1992)
);

NAND3xp33_ASAP7_75t_L g1993 ( 
.A(n_1973),
.B(n_1579),
.C(n_1514),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1979),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1969),
.B(n_1838),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1972),
.B(n_1882),
.Y(n_1996)
);

NOR3x1_ASAP7_75t_L g1997 ( 
.A(n_1962),
.B(n_1606),
.C(n_1598),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1967),
.B(n_1914),
.Y(n_1998)
);

OAI21xp33_ASAP7_75t_L g1999 ( 
.A1(n_1966),
.A2(n_1538),
.B(n_1776),
.Y(n_1999)
);

NOR3xp33_ASAP7_75t_L g2000 ( 
.A(n_1978),
.B(n_1558),
.C(n_1521),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1963),
.B(n_1883),
.Y(n_2001)
);

NAND3xp33_ASAP7_75t_L g2002 ( 
.A(n_1985),
.B(n_1663),
.C(n_1655),
.Y(n_2002)
);

INVx1_ASAP7_75t_SL g2003 ( 
.A(n_1982),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1975),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1970),
.B(n_1883),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1986),
.B(n_1711),
.Y(n_2006)
);

NOR2x1p5_ASAP7_75t_L g2007 ( 
.A(n_2004),
.B(n_1993),
.Y(n_2007)
);

NOR2x1_ASAP7_75t_L g2008 ( 
.A(n_1990),
.B(n_1984),
.Y(n_2008)
);

NOR3xp33_ASAP7_75t_L g2009 ( 
.A(n_1989),
.B(n_1980),
.C(n_1981),
.Y(n_2009)
);

AND4x1_ASAP7_75t_L g2010 ( 
.A(n_1990),
.B(n_1971),
.C(n_1987),
.D(n_1977),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_L g2011 ( 
.A(n_2003),
.B(n_1961),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_1999),
.B(n_1983),
.Y(n_2012)
);

AND4x1_ASAP7_75t_L g2013 ( 
.A(n_2006),
.B(n_1684),
.C(n_1711),
.D(n_1976),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_L g2014 ( 
.A(n_2006),
.B(n_1551),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_2005),
.Y(n_2015)
);

NOR2x1_ASAP7_75t_L g2016 ( 
.A(n_2002),
.B(n_1716),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1992),
.Y(n_2017)
);

NAND4xp75_ASAP7_75t_L g2018 ( 
.A(n_1997),
.B(n_1706),
.C(n_1701),
.D(n_1777),
.Y(n_2018)
);

AOI31xp33_ASAP7_75t_L g2019 ( 
.A1(n_1995),
.A2(n_1550),
.A3(n_1776),
.B(n_1554),
.Y(n_2019)
);

NOR2x1_ASAP7_75t_L g2020 ( 
.A(n_1996),
.B(n_1998),
.Y(n_2020)
);

NOR3xp33_ASAP7_75t_L g2021 ( 
.A(n_1989),
.B(n_1529),
.C(n_1501),
.Y(n_2021)
);

NOR3xp33_ASAP7_75t_L g2022 ( 
.A(n_2000),
.B(n_1542),
.C(n_1710),
.Y(n_2022)
);

AND2x4_ASAP7_75t_L g2023 ( 
.A(n_2007),
.B(n_2000),
.Y(n_2023)
);

NOR2x1_ASAP7_75t_L g2024 ( 
.A(n_2018),
.B(n_1994),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_2017),
.B(n_1988),
.Y(n_2025)
);

AND2x4_ASAP7_75t_L g2026 ( 
.A(n_2021),
.B(n_2001),
.Y(n_2026)
);

NOR3xp33_ASAP7_75t_L g2027 ( 
.A(n_2011),
.B(n_1706),
.C(n_1701),
.Y(n_2027)
);

NOR3xp33_ASAP7_75t_L g2028 ( 
.A(n_2022),
.B(n_1566),
.C(n_1553),
.Y(n_2028)
);

AND2x4_ASAP7_75t_SL g2029 ( 
.A(n_2014),
.B(n_1716),
.Y(n_2029)
);

NOR2x1_ASAP7_75t_SL g2030 ( 
.A(n_2015),
.B(n_1746),
.Y(n_2030)
);

NOR2x1_ASAP7_75t_L g2031 ( 
.A(n_2008),
.B(n_1991),
.Y(n_2031)
);

NAND4xp25_ASAP7_75t_L g2032 ( 
.A(n_2022),
.B(n_1760),
.C(n_1739),
.D(n_1742),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_2013),
.B(n_1746),
.Y(n_2033)
);

NOR2x1_ASAP7_75t_L g2034 ( 
.A(n_2016),
.B(n_2012),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_2010),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2025),
.Y(n_2036)
);

XNOR2xp5_ASAP7_75t_L g2037 ( 
.A(n_2023),
.B(n_2020),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_2035),
.B(n_2009),
.Y(n_2038)
);

OR2x2_ASAP7_75t_L g2039 ( 
.A(n_2026),
.B(n_2019),
.Y(n_2039)
);

NAND3xp33_ASAP7_75t_SL g2040 ( 
.A(n_2033),
.B(n_1578),
.C(n_1577),
.Y(n_2040)
);

OAI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_2024),
.A2(n_1520),
.B1(n_1788),
.B2(n_1852),
.Y(n_2041)
);

AOI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_2034),
.A2(n_1520),
.B1(n_1563),
.B2(n_1680),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_2027),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_2030),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_L g2045 ( 
.A(n_2029),
.B(n_1520),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_2031),
.B(n_1888),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2038),
.B(n_2028),
.Y(n_2047)
);

CKINVDCx11_ASAP7_75t_R g2048 ( 
.A(n_2036),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_2043),
.B(n_2032),
.Y(n_2049)
);

XNOR2xp5_ASAP7_75t_L g2050 ( 
.A(n_2037),
.B(n_2042),
.Y(n_2050)
);

XNOR2xp5_ASAP7_75t_L g2051 ( 
.A(n_2042),
.B(n_1812),
.Y(n_2051)
);

AOI311xp33_ASAP7_75t_L g2052 ( 
.A1(n_2046),
.A2(n_1590),
.A3(n_1718),
.B(n_1720),
.C(n_1719),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_2044),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2039),
.Y(n_2054)
);

INVx1_ASAP7_75t_SL g2055 ( 
.A(n_2045),
.Y(n_2055)
);

AND3x4_ASAP7_75t_L g2056 ( 
.A(n_2040),
.B(n_1698),
.C(n_1690),
.Y(n_2056)
);

NOR4xp25_ASAP7_75t_L g2057 ( 
.A(n_2041),
.B(n_1553),
.C(n_1590),
.D(n_1721),
.Y(n_2057)
);

INVxp67_ASAP7_75t_L g2058 ( 
.A(n_2053),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_2048),
.Y(n_2059)
);

INVx2_ASAP7_75t_SL g2060 ( 
.A(n_2055),
.Y(n_2060)
);

NOR2x1_ASAP7_75t_L g2061 ( 
.A(n_2054),
.B(n_1698),
.Y(n_2061)
);

OAI221xp5_ASAP7_75t_L g2062 ( 
.A1(n_2050),
.A2(n_2057),
.B1(n_2049),
.B2(n_2047),
.C(n_2052),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2051),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_2059),
.B(n_2052),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2060),
.B(n_2056),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2058),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2061),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2063),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2062),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2066),
.Y(n_2070)
);

AOI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_2065),
.A2(n_1712),
.B(n_1674),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2069),
.B(n_1726),
.Y(n_2072)
);

OAI21xp33_ASAP7_75t_SL g2073 ( 
.A1(n_2070),
.A2(n_2064),
.B(n_2068),
.Y(n_2073)
);

OAI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_2071),
.A2(n_2067),
.B1(n_2072),
.B2(n_1563),
.Y(n_2074)
);

AOI21xp33_ASAP7_75t_L g2075 ( 
.A1(n_2073),
.A2(n_2074),
.B(n_1674),
.Y(n_2075)
);

OAI21x1_ASAP7_75t_L g2076 ( 
.A1(n_2075),
.A2(n_1681),
.B(n_1679),
.Y(n_2076)
);

AOI21xp33_ASAP7_75t_L g2077 ( 
.A1(n_2076),
.A2(n_1672),
.B(n_1574),
.Y(n_2077)
);


endmodule