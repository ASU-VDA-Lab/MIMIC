module real_aes_7646_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_449;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_729;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
INVx1_ASAP7_75t_L g516 ( .A(n_1), .Y(n_516) );
INVx1_ASAP7_75t_L g196 ( .A(n_2), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_3), .A2(n_38), .B1(n_158), .B2(n_458), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_4), .Y(n_755) );
AOI21xp33_ASAP7_75t_L g137 ( .A1(n_5), .A2(n_138), .B(n_145), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_6), .B(n_131), .Y(n_507) );
AND2x6_ASAP7_75t_L g143 ( .A(n_7), .B(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_8), .A2(n_237), .B(n_238), .Y(n_236) );
INVx1_ASAP7_75t_L g107 ( .A(n_9), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_9), .B(n_39), .Y(n_121) );
INVx1_ASAP7_75t_L g155 ( .A(n_10), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_11), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g136 ( .A(n_12), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_13), .B(n_168), .Y(n_453) );
INVx1_ASAP7_75t_L g243 ( .A(n_14), .Y(n_243) );
INVx1_ASAP7_75t_L g511 ( .A(n_15), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_16), .B(n_132), .Y(n_492) );
AO32x2_ASAP7_75t_L g473 ( .A1(n_17), .A2(n_131), .A3(n_165), .B1(n_474), .B2(n_478), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_18), .B(n_158), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_19), .B(n_184), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_20), .B(n_132), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_21), .A2(n_50), .B1(n_158), .B2(n_458), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_22), .B(n_138), .Y(n_208) );
AOI22xp33_ASAP7_75t_SL g486 ( .A1(n_23), .A2(n_77), .B1(n_158), .B2(n_168), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_24), .B(n_158), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_25), .B(n_129), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_26), .A2(n_241), .B(n_242), .C(n_244), .Y(n_240) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_27), .A2(n_74), .B1(n_727), .B2(n_728), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_27), .Y(n_728) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_28), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_29), .B(n_161), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_30), .B(n_153), .Y(n_198) );
INVx1_ASAP7_75t_L g174 ( .A(n_31), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_32), .B(n_161), .Y(n_471) );
INVx2_ASAP7_75t_L g141 ( .A(n_33), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_34), .B(n_158), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_35), .B(n_161), .Y(n_459) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_36), .A2(n_62), .B1(n_747), .B2(n_748), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_36), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_37), .A2(n_143), .B(n_148), .C(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_39), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g172 ( .A(n_40), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_41), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_42), .B(n_153), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_43), .B(n_158), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_44), .A2(n_87), .B1(n_215), .B2(n_458), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_45), .B(n_158), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_46), .B(n_158), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_47), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_48), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_49), .B(n_138), .Y(n_231) );
AOI22xp33_ASAP7_75t_SL g496 ( .A1(n_51), .A2(n_60), .B1(n_158), .B2(n_168), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_52), .A2(n_148), .B1(n_168), .B2(n_170), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_53), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_54), .B(n_158), .Y(n_452) );
CKINVDCx16_ASAP7_75t_R g193 ( .A(n_55), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_56), .B(n_158), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g151 ( .A1(n_57), .A2(n_152), .B(n_154), .C(n_157), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_58), .Y(n_261) );
INVx1_ASAP7_75t_L g146 ( .A(n_59), .Y(n_146) );
INVx1_ASAP7_75t_L g144 ( .A(n_61), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_62), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_63), .B(n_158), .Y(n_517) );
INVx1_ASAP7_75t_L g135 ( .A(n_64), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_65), .Y(n_741) );
AO32x2_ASAP7_75t_L g483 ( .A1(n_66), .A2(n_131), .A3(n_223), .B1(n_478), .B2(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g528 ( .A(n_67), .Y(n_528) );
INVx1_ASAP7_75t_L g466 ( .A(n_68), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_SL g183 ( .A1(n_69), .A2(n_157), .B(n_184), .C(n_185), .Y(n_183) );
INVxp67_ASAP7_75t_L g186 ( .A(n_70), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_71), .B(n_168), .Y(n_467) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_73), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_74), .Y(n_727) );
INVx1_ASAP7_75t_L g254 ( .A(n_75), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_76), .A2(n_102), .B1(n_113), .B2(n_758), .Y(n_101) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_78), .A2(n_143), .B(n_148), .C(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_79), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_80), .B(n_168), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_81), .B(n_197), .Y(n_211) );
INVx2_ASAP7_75t_L g133 ( .A(n_82), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_83), .B(n_184), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_84), .B(n_168), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_85), .A2(n_143), .B(n_148), .C(n_195), .Y(n_194) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_86), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g119 ( .A(n_86), .B(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g441 ( .A(n_86), .Y(n_441) );
OR2x2_ASAP7_75t_L g751 ( .A(n_86), .B(n_737), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_88), .A2(n_100), .B1(n_168), .B2(n_169), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_89), .B(n_161), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_90), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_91), .A2(n_143), .B(n_148), .C(n_226), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_92), .Y(n_233) );
INVx1_ASAP7_75t_L g182 ( .A(n_93), .Y(n_182) );
CKINVDCx16_ASAP7_75t_R g239 ( .A(n_94), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_95), .B(n_197), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_96), .B(n_168), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_97), .B(n_131), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_99), .A2(n_138), .B(n_181), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx5_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
CKINVDCx9p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_105), .Y(n_759) );
OR2x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
AND2x2_ASAP7_75t_L g120 ( .A(n_109), .B(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AO221x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_739), .B1(n_742), .B2(n_752), .C(n_754), .Y(n_113) );
OAI222xp33_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_725), .B1(n_726), .B2(n_729), .C1(n_733), .C2(n_738), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_122), .B1(n_439), .B2(n_442), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g730 ( .A(n_119), .Y(n_730) );
OR2x2_ASAP7_75t_L g440 ( .A(n_120), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g737 ( .A(n_120), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_122), .A2(n_731), .B1(n_745), .B2(n_746), .Y(n_744) );
BUFx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g731 ( .A(n_123), .Y(n_731) );
AND3x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_361), .C(n_406), .Y(n_123) );
NOR4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_284), .C(n_325), .D(n_342), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_188), .B(n_204), .C(n_246), .Y(n_125) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_162), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_127), .B(n_189), .Y(n_188) );
NOR4xp25_ASAP7_75t_L g308 ( .A(n_127), .B(n_302), .C(n_309), .D(n_315), .Y(n_308) );
AND2x2_ASAP7_75t_L g381 ( .A(n_127), .B(n_270), .Y(n_381) );
AND2x2_ASAP7_75t_L g400 ( .A(n_127), .B(n_346), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_127), .B(n_395), .Y(n_409) );
AND2x2_ASAP7_75t_L g422 ( .A(n_127), .B(n_203), .Y(n_422) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_SL g267 ( .A(n_128), .Y(n_267) );
AND2x2_ASAP7_75t_L g274 ( .A(n_128), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g324 ( .A(n_128), .B(n_163), .Y(n_324) );
AND2x2_ASAP7_75t_SL g335 ( .A(n_128), .B(n_270), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_128), .B(n_163), .Y(n_339) );
AND2x2_ASAP7_75t_L g348 ( .A(n_128), .B(n_273), .Y(n_348) );
BUFx2_ASAP7_75t_L g371 ( .A(n_128), .Y(n_371) );
AND2x2_ASAP7_75t_L g375 ( .A(n_128), .B(n_179), .Y(n_375) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_137), .B(n_160), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2xp33_ASAP7_75t_SL g217 ( .A(n_130), .B(n_218), .Y(n_217) );
NAND3xp33_ASAP7_75t_L g493 ( .A(n_130), .B(n_478), .C(n_494), .Y(n_493) );
AO21x1_ASAP7_75t_L g531 ( .A1(n_130), .A2(n_494), .B(n_532), .Y(n_531) );
INVx4_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_131), .A2(n_180), .B(n_187), .Y(n_179) );
OA21x2_ASAP7_75t_L g498 ( .A1(n_131), .A2(n_499), .B(n_507), .Y(n_498) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g165 ( .A(n_132), .Y(n_165) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_133), .B(n_134), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
BUFx2_ASAP7_75t_L g237 ( .A(n_138), .Y(n_237) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
NAND2x1p5_ASAP7_75t_L g176 ( .A(n_139), .B(n_143), .Y(n_176) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g506 ( .A(n_140), .Y(n_506) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g149 ( .A(n_141), .Y(n_149) );
INVx1_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
INVx1_ASAP7_75t_L g150 ( .A(n_142), .Y(n_150) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_142), .Y(n_153) );
INVx3_ASAP7_75t_L g156 ( .A(n_142), .Y(n_156) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_142), .Y(n_171) );
INVx1_ASAP7_75t_L g184 ( .A(n_142), .Y(n_184) );
INVx4_ASAP7_75t_SL g159 ( .A(n_143), .Y(n_159) );
OAI21xp5_ASAP7_75t_L g450 ( .A1(n_143), .A2(n_451), .B(n_455), .Y(n_450) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_143), .A2(n_465), .B(n_468), .Y(n_464) );
BUFx3_ASAP7_75t_L g478 ( .A(n_143), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_143), .A2(n_500), .B(n_503), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_143), .A2(n_510), .B(n_514), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_151), .C(n_159), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_147), .A2(n_159), .B(n_182), .C(n_183), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_147), .A2(n_159), .B(n_239), .C(n_240), .Y(n_238) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x6_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_149), .Y(n_158) );
BUFx3_ASAP7_75t_L g215 ( .A(n_149), .Y(n_215) );
INVx1_ASAP7_75t_L g458 ( .A(n_149), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_152), .A2(n_456), .B(n_457), .Y(n_455) );
O2A1O1Ixp5_ASAP7_75t_L g527 ( .A1(n_152), .A2(n_515), .B(n_528), .C(n_529), .Y(n_527) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx4_ASAP7_75t_L g229 ( .A(n_153), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_153), .A2(n_475), .B1(n_476), .B2(n_477), .Y(n_474) );
OAI22xp5_ASAP7_75t_SL g484 ( .A1(n_153), .A2(n_156), .B1(n_485), .B2(n_486), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_153), .A2(n_476), .B1(n_495), .B2(n_496), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_156), .B(n_186), .Y(n_185) );
INVx5_ASAP7_75t_L g197 ( .A(n_156), .Y(n_197) );
O2A1O1Ixp5_ASAP7_75t_SL g465 ( .A1(n_157), .A2(n_197), .B(n_466), .C(n_467), .Y(n_465) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_158), .Y(n_230) );
OAI22xp33_ASAP7_75t_L g166 ( .A1(n_159), .A2(n_167), .B1(n_175), .B2(n_176), .Y(n_166) );
INVx1_ASAP7_75t_L g202 ( .A(n_161), .Y(n_202) );
INVx2_ASAP7_75t_L g223 ( .A(n_161), .Y(n_223) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_161), .A2(n_236), .B(n_245), .Y(n_235) );
OA21x2_ASAP7_75t_L g449 ( .A1(n_161), .A2(n_450), .B(n_459), .Y(n_449) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_161), .A2(n_464), .B(n_471), .Y(n_463) );
OR2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_179), .Y(n_162) );
AND2x2_ASAP7_75t_L g203 ( .A(n_163), .B(n_179), .Y(n_203) );
BUFx2_ASAP7_75t_L g277 ( .A(n_163), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_163), .A2(n_310), .B1(n_312), .B2(n_313), .Y(n_309) );
OR2x2_ASAP7_75t_L g331 ( .A(n_163), .B(n_191), .Y(n_331) );
AND2x2_ASAP7_75t_L g395 ( .A(n_163), .B(n_273), .Y(n_395) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g263 ( .A(n_164), .B(n_191), .Y(n_263) );
AND2x2_ASAP7_75t_L g270 ( .A(n_164), .B(n_179), .Y(n_270) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_164), .Y(n_312) );
OR2x2_ASAP7_75t_L g347 ( .A(n_164), .B(n_190), .Y(n_347) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_177), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_165), .B(n_178), .Y(n_177) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_165), .A2(n_192), .B(n_200), .Y(n_191) );
INVx2_ASAP7_75t_L g216 ( .A(n_165), .Y(n_216) );
INVx2_ASAP7_75t_L g199 ( .A(n_168), .Y(n_199) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OAI22xp5_ASAP7_75t_SL g170 ( .A1(n_171), .A2(n_172), .B1(n_173), .B2(n_174), .Y(n_170) );
INVx2_ASAP7_75t_L g173 ( .A(n_171), .Y(n_173) );
INVx4_ASAP7_75t_L g241 ( .A(n_171), .Y(n_241) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_176), .A2(n_193), .B(n_194), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_176), .A2(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g266 ( .A(n_179), .Y(n_266) );
INVx3_ASAP7_75t_L g275 ( .A(n_179), .Y(n_275) );
BUFx2_ASAP7_75t_L g299 ( .A(n_179), .Y(n_299) );
AND2x2_ASAP7_75t_L g332 ( .A(n_179), .B(n_267), .Y(n_332) );
INVx1_ASAP7_75t_L g454 ( .A(n_184), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_188), .A2(n_418), .B1(n_419), .B2(n_420), .Y(n_417) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_203), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_190), .B(n_275), .Y(n_279) );
INVx1_ASAP7_75t_L g307 ( .A(n_190), .Y(n_307) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx3_ASAP7_75t_L g273 ( .A(n_191), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_198), .C(n_199), .Y(n_195) );
INVx2_ASAP7_75t_L g476 ( .A(n_197), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_197), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_197), .A2(n_525), .B(n_526), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_199), .A2(n_511), .B(n_512), .C(n_513), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_202), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_202), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g285 ( .A(n_203), .Y(n_285) );
NAND2x1_ASAP7_75t_SL g204 ( .A(n_205), .B(n_219), .Y(n_204) );
AND2x2_ASAP7_75t_L g283 ( .A(n_205), .B(n_234), .Y(n_283) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_205), .Y(n_357) );
AND2x2_ASAP7_75t_L g384 ( .A(n_205), .B(n_304), .Y(n_384) );
AND2x2_ASAP7_75t_L g392 ( .A(n_205), .B(n_354), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_205), .B(n_249), .Y(n_419) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g250 ( .A(n_206), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g268 ( .A(n_206), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g289 ( .A(n_206), .Y(n_289) );
INVx1_ASAP7_75t_L g295 ( .A(n_206), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_206), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g328 ( .A(n_206), .B(n_252), .Y(n_328) );
OR2x2_ASAP7_75t_L g366 ( .A(n_206), .B(n_321), .Y(n_366) );
AOI32xp33_ASAP7_75t_L g378 ( .A1(n_206), .A2(n_379), .A3(n_382), .B1(n_383), .B2(n_384), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_206), .B(n_354), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_206), .B(n_314), .Y(n_429) );
OR2x6_ASAP7_75t_L g206 ( .A(n_207), .B(n_217), .Y(n_206) );
AOI21xp5_ASAP7_75t_SL g207 ( .A1(n_208), .A2(n_209), .B(n_216), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_213), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_213), .A2(n_257), .B(n_258), .Y(n_256) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g244 ( .A(n_215), .Y(n_244) );
INVx1_ASAP7_75t_L g259 ( .A(n_216), .Y(n_259) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_216), .A2(n_509), .B(n_518), .Y(n_508) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_216), .A2(n_523), .B(n_530), .Y(n_522) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
OR2x2_ASAP7_75t_L g340 ( .A(n_220), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_234), .Y(n_220) );
INVx1_ASAP7_75t_L g302 ( .A(n_221), .Y(n_302) );
AND2x2_ASAP7_75t_L g304 ( .A(n_221), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_221), .B(n_251), .Y(n_321) );
AND2x2_ASAP7_75t_L g354 ( .A(n_221), .B(n_330), .Y(n_354) );
AND2x2_ASAP7_75t_L g391 ( .A(n_221), .B(n_252), .Y(n_391) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g249 ( .A(n_222), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_222), .B(n_251), .Y(n_281) );
AND2x2_ASAP7_75t_L g288 ( .A(n_222), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g329 ( .A(n_222), .B(n_330), .Y(n_329) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_232), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_231), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_230), .Y(n_226) );
INVx2_ASAP7_75t_L g305 ( .A(n_234), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_234), .B(n_251), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_234), .B(n_296), .Y(n_377) );
INVx1_ASAP7_75t_L g399 ( .A(n_234), .Y(n_399) );
INVx1_ASAP7_75t_L g416 ( .A(n_234), .Y(n_416) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g269 ( .A(n_235), .B(n_251), .Y(n_269) );
AND2x2_ASAP7_75t_L g291 ( .A(n_235), .B(n_252), .Y(n_291) );
INVx1_ASAP7_75t_L g330 ( .A(n_235), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_241), .B(n_243), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_241), .A2(n_469), .B(n_470), .Y(n_468) );
INVx1_ASAP7_75t_L g513 ( .A(n_241), .Y(n_513) );
AOI221x1_ASAP7_75t_SL g246 ( .A1(n_247), .A2(n_262), .B1(n_268), .B2(n_270), .C(n_271), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_247), .A2(n_335), .B1(n_402), .B2(n_403), .Y(n_401) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
AND2x2_ASAP7_75t_L g293 ( .A(n_248), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g388 ( .A(n_248), .B(n_268), .Y(n_388) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g344 ( .A(n_249), .B(n_269), .Y(n_344) );
INVx1_ASAP7_75t_L g356 ( .A(n_250), .Y(n_356) );
AND2x2_ASAP7_75t_L g367 ( .A(n_250), .B(n_354), .Y(n_367) );
AND2x2_ASAP7_75t_L g434 ( .A(n_250), .B(n_329), .Y(n_434) );
INVx2_ASAP7_75t_L g296 ( .A(n_251), .Y(n_296) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_259), .B(n_260), .Y(n_252) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_263), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g386 ( .A(n_263), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_264), .B(n_347), .Y(n_350) );
INVx3_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g430 ( .A1(n_265), .A2(n_386), .B(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
NOR2xp33_ASAP7_75t_SL g408 ( .A(n_268), .B(n_294), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_269), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g360 ( .A(n_269), .B(n_288), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_269), .B(n_295), .Y(n_437) );
AND2x2_ASAP7_75t_L g306 ( .A(n_270), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g373 ( .A(n_270), .Y(n_373) );
AOI21xp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_276), .B(n_280), .Y(n_271) );
NAND2x1_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_273), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g322 ( .A(n_273), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g334 ( .A(n_273), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_273), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g358 ( .A(n_274), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_274), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_274), .B(n_277), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AOI211xp5_ASAP7_75t_L g345 ( .A1(n_277), .A2(n_316), .B(n_346), .C(n_348), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_277), .A2(n_364), .B1(n_367), .B2(n_368), .C(n_372), .Y(n_363) );
AND2x2_ASAP7_75t_L g359 ( .A(n_278), .B(n_312), .Y(n_359) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g319 ( .A(n_283), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g390 ( .A(n_283), .B(n_391), .Y(n_390) );
OAI211xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_286), .B(n_292), .C(n_317), .Y(n_284) );
NAND3xp33_ASAP7_75t_SL g403 ( .A(n_285), .B(n_404), .C(n_405), .Y(n_403) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
OR2x2_ASAP7_75t_L g376 ( .A(n_287), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_297), .B1(n_300), .B2(n_306), .C(n_308), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_294), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_294), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g316 ( .A(n_299), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_299), .A2(n_356), .B1(n_357), .B2(n_358), .Y(n_355) );
OR2x2_ASAP7_75t_L g436 ( .A(n_299), .B(n_347), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVxp67_ASAP7_75t_L g410 ( .A(n_302), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_304), .B(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g311 ( .A(n_305), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_307), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_307), .B(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_307), .B(n_374), .Y(n_413) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_311), .Y(n_337) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g427 ( .A(n_316), .B(n_347), .Y(n_427) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_322), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g405 ( .A(n_322), .Y(n_405) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI322xp33_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_331), .A3(n_332), .B1(n_333), .B2(n_336), .C1(n_338), .C2(n_340), .Y(n_325) );
OAI322xp33_ASAP7_75t_L g407 ( .A1(n_326), .A2(n_408), .A3(n_409), .B1(n_410), .B2(n_411), .C1(n_412), .C2(n_414), .Y(n_407) );
CKINVDCx16_ASAP7_75t_R g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx4_ASAP7_75t_L g341 ( .A(n_328), .Y(n_341) );
AND2x2_ASAP7_75t_L g402 ( .A(n_328), .B(n_354), .Y(n_402) );
AND2x2_ASAP7_75t_L g415 ( .A(n_328), .B(n_416), .Y(n_415) );
CKINVDCx16_ASAP7_75t_R g426 ( .A(n_331), .Y(n_426) );
INVx1_ASAP7_75t_L g404 ( .A(n_332), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
OR2x2_ASAP7_75t_L g338 ( .A(n_334), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g421 ( .A(n_334), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_334), .B(n_375), .Y(n_432) );
OR2x2_ASAP7_75t_L g365 ( .A(n_337), .B(n_366), .Y(n_365) );
INVxp33_ASAP7_75t_L g382 ( .A(n_337), .Y(n_382) );
OAI221xp5_ASAP7_75t_SL g342 ( .A1(n_341), .A2(n_343), .B1(n_345), .B2(n_349), .C(n_351), .Y(n_342) );
NOR2xp67_ASAP7_75t_L g398 ( .A(n_341), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g425 ( .A(n_341), .Y(n_425) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx3_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AOI322xp5_ASAP7_75t_L g389 ( .A1(n_348), .A2(n_373), .A3(n_390), .B1(n_392), .B2(n_393), .C1(n_396), .C2(n_400), .Y(n_389) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_355), .B1(n_359), .B2(n_360), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_385), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_363), .B(n_378), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_366), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
NAND2xp33_ASAP7_75t_SL g383 ( .A(n_369), .B(n_380), .Y(n_383) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
OAI322xp33_ASAP7_75t_L g423 ( .A1(n_371), .A2(n_424), .A3(n_426), .B1(n_427), .B2(n_428), .C1(n_430), .C2(n_433), .Y(n_423) );
AOI21xp33_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_374), .B(n_376), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_381), .B(n_429), .Y(n_438) );
OAI211xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_387), .B(n_389), .C(n_401), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NOR4xp25_ASAP7_75t_L g406 ( .A(n_407), .B(n_417), .C(n_423), .D(n_435), .Y(n_406) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
CKINVDCx14_ASAP7_75t_R g433 ( .A(n_434), .Y(n_433) );
OAI21xp5_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_437), .B(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx6_ASAP7_75t_L g732 ( .A(n_440), .Y(n_732) );
NOR2x2_ASAP7_75t_L g736 ( .A(n_441), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_443), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_729) );
OR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_647), .Y(n_443) );
NAND5xp2_ASAP7_75t_L g444 ( .A(n_445), .B(n_566), .C(n_581), .D(n_607), .E(n_629), .Y(n_444) );
NOR2xp33_ASAP7_75t_SL g445 ( .A(n_446), .B(n_546), .Y(n_445) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_487), .B1(n_519), .B2(n_535), .C(n_536), .Y(n_446) );
NOR2xp33_ASAP7_75t_SL g447 ( .A(n_448), .B(n_479), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_448), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_SL g723 ( .A(n_448), .Y(n_723) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_460), .Y(n_448) );
INVx1_ASAP7_75t_L g563 ( .A(n_449), .Y(n_563) );
AND2x2_ASAP7_75t_L g565 ( .A(n_449), .B(n_473), .Y(n_565) );
AND2x2_ASAP7_75t_L g575 ( .A(n_449), .B(n_472), .Y(n_575) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_449), .Y(n_593) );
INVx1_ASAP7_75t_L g603 ( .A(n_449), .Y(n_603) );
OR2x2_ASAP7_75t_L g641 ( .A(n_449), .B(n_540), .Y(n_641) );
INVx2_ASAP7_75t_L g691 ( .A(n_449), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_449), .B(n_539), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B(n_454), .Y(n_451) );
NOR2xp67_ASAP7_75t_L g460 ( .A(n_461), .B(n_472), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_462), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_462), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_SL g623 ( .A(n_462), .B(n_563), .Y(n_623) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_463), .Y(n_481) );
INVx2_ASAP7_75t_L g540 ( .A(n_463), .Y(n_540) );
OR2x2_ASAP7_75t_L g602 ( .A(n_463), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g541 ( .A(n_472), .B(n_483), .Y(n_541) );
AND2x2_ASAP7_75t_L g558 ( .A(n_472), .B(n_538), .Y(n_558) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g482 ( .A(n_473), .B(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_L g561 ( .A(n_473), .Y(n_561) );
AND2x2_ASAP7_75t_L g690 ( .A(n_473), .B(n_691), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_476), .A2(n_504), .B(n_505), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_476), .A2(n_515), .B(n_516), .C(n_517), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_478), .A2(n_524), .B(n_527), .Y(n_523) );
INVx1_ASAP7_75t_L g535 ( .A(n_479), .Y(n_535) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
AND2x2_ASAP7_75t_L g653 ( .A(n_480), .B(n_541), .Y(n_653) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g654 ( .A(n_481), .B(n_565), .Y(n_654) );
O2A1O1Ixp33_ASAP7_75t_L g621 ( .A1(n_482), .A2(n_622), .B(n_624), .C(n_626), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_482), .B(n_622), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_482), .A2(n_552), .B1(n_695), .B2(n_696), .C(n_698), .Y(n_694) );
INVx1_ASAP7_75t_L g538 ( .A(n_483), .Y(n_538) );
INVx1_ASAP7_75t_L g574 ( .A(n_483), .Y(n_574) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_483), .Y(n_583) );
INVx1_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_497), .Y(n_488) );
AND2x2_ASAP7_75t_L g600 ( .A(n_489), .B(n_545), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_489), .B(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_490), .B(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g692 ( .A(n_490), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g724 ( .A(n_490), .Y(n_724) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g554 ( .A(n_491), .Y(n_554) );
AND2x2_ASAP7_75t_L g580 ( .A(n_491), .B(n_534), .Y(n_580) );
NOR2x1_ASAP7_75t_L g589 ( .A(n_491), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g596 ( .A(n_491), .B(n_597), .Y(n_596) );
AND2x4_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g532 ( .A(n_492), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_497), .B(n_636), .Y(n_671) );
INVx1_ASAP7_75t_SL g675 ( .A(n_497), .Y(n_675) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_508), .Y(n_497) );
INVx3_ASAP7_75t_L g534 ( .A(n_498), .Y(n_534) );
AND2x2_ASAP7_75t_L g545 ( .A(n_498), .B(n_522), .Y(n_545) );
AND2x2_ASAP7_75t_L g567 ( .A(n_498), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g612 ( .A(n_498), .B(n_606), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_498), .B(n_544), .Y(n_693) );
INVx2_ASAP7_75t_L g515 ( .A(n_506), .Y(n_515) );
AND2x2_ASAP7_75t_L g533 ( .A(n_508), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g544 ( .A(n_508), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_508), .B(n_522), .Y(n_569) );
AND2x2_ASAP7_75t_L g605 ( .A(n_508), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_533), .Y(n_520) );
INVx1_ASAP7_75t_L g585 ( .A(n_521), .Y(n_585) );
AND2x2_ASAP7_75t_L g627 ( .A(n_521), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_521), .B(n_548), .Y(n_633) );
AOI21xp5_ASAP7_75t_SL g707 ( .A1(n_521), .A2(n_539), .B(n_562), .Y(n_707) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_531), .Y(n_521) );
OR2x2_ASAP7_75t_L g550 ( .A(n_522), .B(n_531), .Y(n_550) );
AND2x2_ASAP7_75t_L g597 ( .A(n_522), .B(n_534), .Y(n_597) );
INVx2_ASAP7_75t_L g606 ( .A(n_522), .Y(n_606) );
INVx1_ASAP7_75t_L g712 ( .A(n_522), .Y(n_712) );
AND2x2_ASAP7_75t_L g636 ( .A(n_531), .B(n_606), .Y(n_636) );
INVx1_ASAP7_75t_L g661 ( .A(n_531), .Y(n_661) );
AND2x2_ASAP7_75t_L g570 ( .A(n_533), .B(n_554), .Y(n_570) );
AND2x2_ASAP7_75t_L g582 ( .A(n_533), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_SL g700 ( .A(n_533), .Y(n_700) );
INVx2_ASAP7_75t_L g590 ( .A(n_534), .Y(n_590) );
AND2x2_ASAP7_75t_L g628 ( .A(n_534), .B(n_544), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_534), .B(n_712), .Y(n_711) );
OAI21xp33_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_541), .B(n_542), .Y(n_536) );
AND2x2_ASAP7_75t_L g643 ( .A(n_537), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g697 ( .A(n_537), .Y(n_697) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g617 ( .A(n_538), .Y(n_617) );
BUFx2_ASAP7_75t_L g716 ( .A(n_538), .Y(n_716) );
BUFx2_ASAP7_75t_L g587 ( .A(n_539), .Y(n_587) );
AND2x2_ASAP7_75t_L g689 ( .A(n_539), .B(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g672 ( .A(n_540), .Y(n_672) );
AND2x4_ASAP7_75t_L g599 ( .A(n_541), .B(n_562), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_541), .B(n_623), .Y(n_635) );
AOI32xp33_ASAP7_75t_L g559 ( .A1(n_542), .A2(n_560), .A3(n_562), .B1(n_564), .B2(n_565), .Y(n_559) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
INVx3_ASAP7_75t_L g548 ( .A(n_543), .Y(n_548) );
OR2x2_ASAP7_75t_L g684 ( .A(n_543), .B(n_640), .Y(n_684) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g553 ( .A(n_544), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g660 ( .A(n_544), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g552 ( .A(n_545), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g564 ( .A(n_545), .B(n_554), .Y(n_564) );
INVx1_ASAP7_75t_L g685 ( .A(n_545), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_545), .B(n_660), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_551), .B(n_555), .C(n_559), .Y(n_546) );
OAI322xp33_ASAP7_75t_L g655 ( .A1(n_547), .A2(n_592), .A3(n_656), .B1(n_658), .B2(n_662), .C1(n_663), .C2(n_667), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
INVxp67_ASAP7_75t_L g620 ( .A(n_548), .Y(n_620) );
INVx1_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g674 ( .A(n_550), .B(n_675), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_550), .B(n_590), .Y(n_721) );
INVxp67_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g613 ( .A(n_553), .Y(n_613) );
OR2x2_ASAP7_75t_L g699 ( .A(n_554), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_557), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g608 ( .A(n_558), .B(n_587), .Y(n_608) );
AND2x2_ASAP7_75t_L g679 ( .A(n_558), .B(n_592), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_558), .B(n_666), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g566 ( .A1(n_560), .A2(n_567), .B1(n_570), .B2(n_571), .C(n_576), .Y(n_566) );
OR2x2_ASAP7_75t_L g577 ( .A(n_560), .B(n_573), .Y(n_577) );
AND2x2_ASAP7_75t_L g665 ( .A(n_560), .B(n_666), .Y(n_665) );
AOI32xp33_ASAP7_75t_L g704 ( .A1(n_560), .A2(n_590), .A3(n_705), .B1(n_706), .B2(n_709), .Y(n_704) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_561), .B(n_597), .C(n_620), .Y(n_638) );
AND2x2_ASAP7_75t_L g664 ( .A(n_561), .B(n_657), .Y(n_664) );
INVxp67_ASAP7_75t_L g644 ( .A(n_562), .Y(n_644) );
BUFx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_565), .B(n_617), .Y(n_673) );
INVx2_ASAP7_75t_L g683 ( .A(n_565), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_565), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g652 ( .A(n_568), .Y(n_652) );
OR2x2_ASAP7_75t_L g578 ( .A(n_569), .B(n_579), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_571), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_574), .Y(n_657) );
AND2x2_ASAP7_75t_L g616 ( .A(n_575), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g662 ( .A(n_575), .Y(n_662) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_575), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
AOI21xp33_ASAP7_75t_SL g601 ( .A1(n_577), .A2(n_602), .B(n_604), .Y(n_601) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g695 ( .A(n_580), .B(n_605), .Y(n_695) );
AOI211xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_584), .B(n_594), .C(n_601), .Y(n_581) );
AND2x2_ASAP7_75t_L g625 ( .A(n_583), .B(n_593), .Y(n_625) );
INVx2_ASAP7_75t_L g640 ( .A(n_583), .Y(n_640) );
OR2x2_ASAP7_75t_L g678 ( .A(n_583), .B(n_641), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_583), .B(n_721), .Y(n_720) );
AOI211xp5_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_586), .B(n_588), .C(n_591), .Y(n_584) );
INVxp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_587), .B(n_625), .Y(n_624) );
OAI211xp5_ASAP7_75t_L g706 ( .A1(n_588), .A2(n_683), .B(n_707), .C(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2x1p5_ASAP7_75t_L g604 ( .A(n_589), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g646 ( .A(n_590), .B(n_636), .Y(n_646) );
INVx1_ASAP7_75t_L g651 ( .A(n_590), .Y(n_651) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_595), .B(n_598), .Y(n_594) );
INVxp33_ASAP7_75t_L g702 ( .A(n_596), .Y(n_702) );
AND2x2_ASAP7_75t_L g681 ( .A(n_597), .B(n_660), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_602), .A2(n_664), .B(n_665), .Y(n_663) );
OAI322xp33_ASAP7_75t_L g682 ( .A1(n_604), .A2(n_683), .A3(n_684), .B1(n_685), .B2(n_686), .C1(n_688), .C2(n_692), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B1(n_614), .B2(n_618), .C(n_621), .Y(n_607) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g659 ( .A(n_612), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g703 ( .A(n_616), .Y(n_703) );
INVxp67_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_619), .B(n_639), .Y(n_705) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g668 ( .A(n_628), .B(n_636), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .B1(n_634), .B2(n_636), .C(n_637), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_632), .A2(n_649), .B1(n_653), .B2(n_654), .C(n_655), .Y(n_648) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVxp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_636), .B(n_651), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B1(n_642), .B2(n_645), .Y(n_637) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx2_ASAP7_75t_SL g666 ( .A(n_641), .Y(n_666) );
INVxp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND5xp2_ASAP7_75t_L g647 ( .A(n_648), .B(n_669), .C(n_694), .D(n_704), .E(n_714), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_650), .B(n_652), .Y(n_649) );
NOR4xp25_ASAP7_75t_L g722 ( .A(n_651), .B(n_657), .C(n_723), .D(n_724), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_654), .A2(n_715), .B1(n_717), .B2(n_719), .C(n_722), .Y(n_714) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g713 ( .A(n_660), .Y(n_713) );
OAI322xp33_ASAP7_75t_L g670 ( .A1(n_664), .A2(n_671), .A3(n_672), .B1(n_673), .B2(n_674), .C1(n_676), .C2(n_680), .Y(n_670) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_682), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g715 ( .A(n_690), .B(n_716), .Y(n_715) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_698) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
OR2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_713), .Y(n_710) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
BUFx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_SL g753 ( .A(n_740), .Y(n_753) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_744), .B(n_749), .Y(n_743) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_SL g757 ( .A(n_751), .Y(n_757) );
BUFx3_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
endmodule