module real_jpeg_10717_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_311, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_311;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_52),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_3),
.A2(n_52),
.B1(n_59),
.B2(n_60),
.Y(n_120)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_5),
.A2(n_32),
.B(n_43),
.C(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_5),
.B(n_32),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_8),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_8),
.A2(n_59),
.B1(n_60),
.B2(n_153),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_153),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_8),
.A2(n_27),
.B1(n_35),
.B2(n_153),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_9),
.A2(n_27),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_9),
.A2(n_38),
.B1(n_45),
.B2(n_46),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_9),
.A2(n_38),
.B1(n_59),
.B2(n_60),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_10),
.A2(n_59),
.B1(n_60),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_10),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_144),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_144),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_10),
.A2(n_27),
.B1(n_35),
.B2(n_144),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_11),
.A2(n_27),
.B1(n_35),
.B2(n_50),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_11),
.A2(n_50),
.B1(n_59),
.B2(n_60),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_12),
.A2(n_45),
.B(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_12),
.B(n_45),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_12),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_12),
.A2(n_82),
.B1(n_85),
.B2(n_162),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_12),
.A2(n_32),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_12),
.B(n_32),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_12),
.B(n_209),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g228 ( 
.A1(n_12),
.A2(n_29),
.B(n_33),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_12),
.A2(n_27),
.B1(n_35),
.B2(n_164),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_14),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_63),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_15),
.A2(n_27),
.B1(n_35),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_15),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_15),
.A2(n_59),
.B1(n_60),
.B2(n_92),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_15),
.A2(n_45),
.B1(n_46),
.B2(n_92),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_92),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_16),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_16),
.A2(n_36),
.B1(n_59),
.B2(n_60),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_16),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_17),
.A2(n_27),
.B1(n_35),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_17),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_17),
.A2(n_59),
.B1(n_60),
.B2(n_126),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_17),
.A2(n_45),
.B1(n_46),
.B2(n_126),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_126),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_107),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_93),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_22),
.B(n_93),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_65),
.C(n_78),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_23),
.A2(n_65),
.B1(n_66),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_23),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_24),
.A2(n_25),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_25),
.B(n_53),
.C(n_64),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_26),
.A2(n_31),
.B1(n_34),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_26),
.A2(n_31),
.B1(n_37),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_26),
.A2(n_31),
.B1(n_91),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_26),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_26),
.A2(n_31),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_26),
.A2(n_31),
.B1(n_125),
.B2(n_260),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_28),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_27),
.A2(n_28),
.B(n_164),
.C(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_31),
.Y(n_209)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_53),
.B1(n_54),
.B2(n_64),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_48),
.B2(n_51),
.Y(n_41)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_42),
.A2(n_44),
.B1(n_51),
.B2(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_42),
.A2(n_44),
.B1(n_70),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_42),
.A2(n_44),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_42),
.A2(n_44),
.B1(n_189),
.B2(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_42),
.A2(n_44),
.B1(n_205),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_42),
.A2(n_44),
.B1(n_244),
.B2(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_42),
.A2(n_44),
.B1(n_129),
.B2(n_256),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_43),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_44),
.B(n_164),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_56),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_45),
.B(n_47),
.Y(n_193)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_46),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_53),
.A2(n_54),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_58),
.B(n_62),
.Y(n_54)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_58),
.B1(n_74),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_55),
.A2(n_58),
.B1(n_88),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_55),
.A2(n_58),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_55),
.A2(n_58),
.B1(n_152),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_55),
.A2(n_58),
.B1(n_177),
.B2(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_55),
.A2(n_58),
.B1(n_185),
.B2(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_55),
.A2(n_58),
.B1(n_122),
.B2(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_56),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_56),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_57),
.Y(n_157)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_58),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_59),
.B(n_61),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_59),
.B(n_168),
.Y(n_167)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_60),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_66),
.A2(n_67),
.B(n_72),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_72),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_75),
.A2(n_77),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_89),
.B(n_90),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_80),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_81),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_89),
.B1(n_90),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_81),
.A2(n_87),
.B1(n_89),
.B2(n_291),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B(n_86),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_82),
.A2(n_85),
.B1(n_143),
.B2(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_82),
.A2(n_85),
.B1(n_146),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_82),
.A2(n_85),
.B1(n_179),
.B2(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_82),
.A2(n_85),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_82),
.A2(n_85),
.B1(n_120),
.B2(n_232),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_83),
.A2(n_84),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_83),
.A2(n_84),
.B1(n_197),
.B2(n_211),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_84),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_85),
.B(n_164),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_87),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_105),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B1(n_100),
.B2(n_104),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_101),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_133),
.B(n_309),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_130),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_109),
.B(n_130),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_116),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_110),
.A2(n_114),
.B1(n_115),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_110),
.Y(n_296)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_116),
.A2(n_117),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_123),
.C(n_127),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_118),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_119),
.B(n_121),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

AOI321xp33_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_285),
.A3(n_297),
.B1(n_303),
.B2(n_308),
.C(n_311),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_250),
.C(n_281),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_221),
.B(n_249),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_199),
.B(n_220),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_181),
.B(n_198),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_171),
.B(n_180),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_159),
.B(n_170),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_147),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_141),
.B(n_147),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_154),
.B2(n_158),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_148),
.B(n_158),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_151),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_154),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_165),
.B(n_169),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_163),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_172),
.B(n_173),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_176),
.C(n_178),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_182),
.B(n_183),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_183),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_186),
.CI(n_190),
.CON(n_183),
.SN(n_183)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_188),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_195),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_200),
.B(n_201),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_213),
.B2(n_214),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_216),
.C(n_218),
.Y(n_222)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_206),
.B1(n_207),
.B2(n_212),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_204),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_210),
.C(n_212),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_209),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_211),
.Y(n_231)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_215),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_216),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_217),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_223),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_236),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_225),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_225),
.B(n_235),
.C(n_236),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_229),
.B2(n_230),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_230),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_245),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_242),
.B2(n_243),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_242),
.C(n_245),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_241),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_248),
.Y(n_259)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

AOI21xp33_ASAP7_75t_L g304 ( 
.A1(n_251),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_268),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_252),
.B(n_268),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_263),
.C(n_267),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_262),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_257),
.B1(n_258),
.B2(n_261),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_255),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_SL g279 ( 
.A(n_257),
.B(n_261),
.C(n_262),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_267),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_265),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_279),
.B2(n_280),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_272),
.C(n_280),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_276),
.C(n_278),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_275),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_279),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_283),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_293),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_286),
.B(n_293),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_290),
.C(n_292),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_290),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_304),
.B(n_307),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_299),
.B(n_300),
.Y(n_307)
);


endmodule