module real_jpeg_6730_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_1),
.A2(n_25),
.B1(n_103),
.B2(n_106),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_1),
.A2(n_25),
.B1(n_165),
.B2(n_168),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_1),
.A2(n_25),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_1),
.B(n_31),
.Y(n_274)
);

O2A1O1Ixp33_ASAP7_75t_L g331 ( 
.A1(n_1),
.A2(n_263),
.B(n_332),
.C(n_333),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_1),
.B(n_356),
.C(n_357),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_1),
.B(n_138),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_1),
.B(n_193),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_1),
.B(n_94),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_2),
.A2(n_44),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_2),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_2),
.A2(n_212),
.B1(n_247),
.B2(n_250),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_2),
.A2(n_212),
.B1(n_345),
.B2(n_347),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_2),
.A2(n_212),
.B1(n_366),
.B2(n_368),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_3),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_3),
.Y(n_167)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_3),
.Y(n_200)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_4),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_5),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_5),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_5),
.Y(n_193)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_5),
.Y(n_278)
);

INVx8_ASAP7_75t_L g384 ( 
.A(n_5),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_6),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_6),
.A2(n_45),
.B1(n_133),
.B2(n_136),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_6),
.A2(n_45),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_6),
.A2(n_45),
.B1(n_198),
.B2(n_201),
.Y(n_197)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_10),
.Y(n_216)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_11),
.Y(n_85)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_11),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_11),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g356 ( 
.A(n_11),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_12),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_12),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_12),
.A2(n_127),
.B1(n_173),
.B2(n_177),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_12),
.A2(n_127),
.B1(n_214),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_12),
.A2(n_127),
.B1(n_267),
.B2(n_269),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_13),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_440),
.Y(n_19)
);

OAI221xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_59),
.B1(n_63),
.B2(n_435),
.C(n_438),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_21),
.B(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_21),
.B(n_59),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_22),
.B(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_23),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_31),
.Y(n_23)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_24),
.B(n_48),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_28),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_25),
.B(n_29),
.Y(n_28)
);

OAI21xp33_ASAP7_75t_L g333 ( 
.A1(n_25),
.A2(n_334),
.B(n_337),
.Y(n_333)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVxp33_ASAP7_75t_L g260 ( 
.A(n_28),
.Y(n_260)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_31),
.B(n_41),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_31),
.B(n_211),
.Y(n_241)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_31)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_32),
.Y(n_259)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_34),
.Y(n_126)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_36),
.Y(n_117)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_36),
.Y(n_135)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_36),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_36),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_36),
.Y(n_263)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_38),
.Y(n_206)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_38),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_40),
.A2(n_61),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_40),
.B(n_241),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_48),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_48),
.B(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_54),
.B2(n_57),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_53),
.Y(n_264)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_58),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_59),
.A2(n_154),
.B(n_179),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_59),
.A2(n_156),
.B1(n_179),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_59),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B(n_62),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_60),
.A2(n_72),
.B(n_223),
.Y(n_431)
);

A2O1A1O1Ixp25_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_234),
.B(n_424),
.C(n_427),
.D(n_434),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_217),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_180),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_66),
.B(n_180),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_153),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_139),
.B2(n_140),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_69),
.B(n_139),
.C(n_153),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_70),
.A2(n_71),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_71),
.B(n_76),
.C(n_109),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_71),
.B(n_220),
.C(n_232),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_72),
.B(n_210),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_73),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_108),
.B2(n_109),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_76),
.A2(n_77),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_76),
.A2(n_77),
.B1(n_243),
.B2(n_253),
.Y(n_242)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_77),
.B(n_240),
.C(n_243),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_77),
.B(n_228),
.C(n_231),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_100),
.B(n_101),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_78),
.A2(n_172),
.B(n_178),
.Y(n_171)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_79),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_79),
.B(n_102),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_79),
.B(n_344),
.Y(n_343)
);

NOR2x1_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_94),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B1(n_86),
.B2(n_90),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_83),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AO22x1_ASAP7_75t_SL g94 ( 
.A1(n_88),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_94)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_113),
.B1(n_121),
.B2(n_123),
.Y(n_120)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_91),
.Y(n_346)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_93),
.Y(n_177)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_94),
.B(n_145),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_94),
.B(n_344),
.Y(n_360)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_97),
.Y(n_201)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_97),
.Y(n_268)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_100),
.B(n_101),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_100),
.A2(n_144),
.B(n_172),
.Y(n_202)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_107),
.B(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_125),
.B(n_130),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_110),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_110),
.B(n_246),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_110),
.A2(n_138),
.B(n_205),
.Y(n_301)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_111),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_120),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_114),
.Y(n_336)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_115),
.Y(n_332)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_117),
.Y(n_208)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_120),
.B(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_138),
.B(n_151),
.Y(n_150)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_131),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_131),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_138),
.Y(n_131)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_138),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_140),
.A2(n_141),
.B(n_150),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_150),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_142),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_144),
.B(n_360),
.Y(n_404)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_149),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_151),
.B(n_229),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_151),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_155),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_171),
.Y(n_155)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_156),
.A2(n_171),
.B1(n_179),
.B2(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_156),
.B(n_331),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_156),
.A2(n_179),
.B1(n_331),
.B2(n_407),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_162),
.B(n_164),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_157),
.B(n_164),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_157),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_157),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_167),
.Y(n_358)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_171),
.Y(n_313)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g285 ( 
.A(n_178),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_178),
.B(n_343),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.C(n_187),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_181),
.A2(n_185),
.B1(n_186),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_181),
.Y(n_317)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_187),
.B(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_203),
.C(n_209),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_188),
.A2(n_189),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_202),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_190),
.B(n_202),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_191),
.B(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_192),
.A2(n_196),
.B(n_266),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_195),
.B(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_197),
.B(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_198),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_199),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_200),
.Y(n_367)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_201),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_203),
.B(n_209),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_204),
.B(n_245),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g230 ( 
.A(n_205),
.Y(n_230)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI32xp33_ASAP7_75t_L g256 ( 
.A1(n_214),
.A2(n_257),
.A3(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_256)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_217),
.A2(n_425),
.B(n_426),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_233),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_218),
.B(n_233),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_232),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_225),
.B1(n_226),
.B2(n_231),
.Y(n_221)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_222),
.Y(n_231)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_229),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_416),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_306),
.C(n_321),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_293),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_279),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_238),
.B(n_279),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_254),
.C(n_270),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_239),
.B(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_243),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_254),
.A2(n_255),
.B1(n_270),
.B2(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_265),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_256),
.B(n_265),
.Y(n_288)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp33_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

INVx6_ASAP7_75t_SL g262 ( 
.A(n_263),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_277),
.B(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_270),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.C(n_275),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_271),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_275),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_276),
.B(n_380),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_277),
.B(n_364),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_287),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_282),
.C(n_287),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_285),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_286),
.B(n_360),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_290),
.C(n_291),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_293),
.A2(n_419),
.B(n_420),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_305),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_294),
.B(n_305),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_297),
.C(n_298),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_302),
.C(n_303),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_301),
.A2(n_303),
.B1(n_430),
.B2(n_431),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_301),
.B(n_431),
.C(n_432),
.Y(n_437)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_302),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_318),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_307),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_315),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_308),
.B(n_315),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_312),
.C(n_314),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g319 ( 
.A(n_309),
.B(n_312),
.CI(n_314),
.CON(n_319),
.SN(n_319)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_318),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_319),
.B(n_320),
.Y(n_421)
);

BUFx24_ASAP7_75t_SL g441 ( 
.A(n_319),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_348),
.B(n_415),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_326),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_323),
.B(n_326),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_330),
.C(n_340),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_327),
.B(n_411),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_330),
.A2(n_340),
.B1(n_341),
.B2(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_331),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_339),
.Y(n_347)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_409),
.B(n_414),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_350),
.A2(n_399),
.B(n_408),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_374),
.B(n_398),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_361),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_352),
.B(n_361),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_359),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_353),
.A2(n_354),
.B1(n_359),
.B2(n_377),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_359),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_369),
.Y(n_361)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_362),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_381),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_370),
.A2(n_371),
.B1(n_372),
.B2(n_373),
.Y(n_369)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_370),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_371),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_372),
.C(n_401),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_375),
.A2(n_385),
.B(n_397),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_378),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_378),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx8_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_393),
.B(n_396),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_392),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_391),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx6_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_394),
.B(n_395),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_402),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_402),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_406),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_404),
.B(n_405),
.C(n_406),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_413),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_410),
.B(n_413),
.Y(n_414)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g416 ( 
.A1(n_417),
.A2(n_418),
.B(n_421),
.C(n_422),
.D(n_423),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_433),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_428),
.B(n_433),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_432),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_437),
.Y(n_439)
);


endmodule