module real_aes_16284_n_376 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1888;
wire n_1217;
wire n_1423;
wire n_571;
wire n_1034;
wire n_1328;
wire n_549;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_1382;
wire n_951;
wire n_875;
wire n_1199;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1893;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1914;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1760;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_733;
wire n_602;
wire n_402;
wire n_1404;
wire n_676;
wire n_658;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1855;
wire n_1605;
wire n_1592;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_1838;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1790;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1457;
wire n_465;
wire n_719;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_1777;
wire n_458;
wire n_444;
wire n_1200;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_517;
wire n_1851;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1891;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1925;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1868;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1280;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g1125 ( .A(n_0), .Y(n_1125) );
AOI22xp33_ASAP7_75t_SL g1460 ( .A1(n_1), .A2(n_331), .B1(n_725), .B2(n_1169), .Y(n_1460) );
INVxp67_ASAP7_75t_SL g1480 ( .A(n_1), .Y(n_1480) );
INVx1_ASAP7_75t_L g898 ( .A(n_2), .Y(n_898) );
AO22x1_ASAP7_75t_L g923 ( .A1(n_2), .A2(n_251), .B1(n_526), .B2(n_609), .Y(n_923) );
INVx1_ASAP7_75t_L g389 ( .A(n_3), .Y(n_389) );
AND2x2_ASAP7_75t_L g460 ( .A(n_3), .B(n_272), .Y(n_460) );
AND2x2_ASAP7_75t_L g477 ( .A(n_3), .B(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_3), .B(n_399), .Y(n_696) );
INVx1_ASAP7_75t_L g907 ( .A(n_4), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_4), .A2(n_136), .B1(n_479), .B2(n_493), .Y(n_922) );
AOI22xp33_ASAP7_75t_SL g1212 ( .A1(n_5), .A2(n_334), .B1(n_467), .B2(n_1169), .Y(n_1212) );
AOI221xp5_ASAP7_75t_L g1226 ( .A1(n_5), .A2(n_7), .B1(n_498), .B2(n_1227), .C(n_1229), .Y(n_1226) );
AOI22xp33_ASAP7_75t_SL g1493 ( .A1(n_6), .A2(n_52), .B1(n_724), .B2(n_725), .Y(n_1493) );
INVxp67_ASAP7_75t_SL g1515 ( .A(n_6), .Y(n_1515) );
AOI22xp33_ASAP7_75t_SL g1217 ( .A1(n_7), .A2(n_13), .B1(n_642), .B2(n_1026), .Y(n_1217) );
AOI22xp33_ASAP7_75t_SL g1168 ( .A1(n_8), .A2(n_330), .B1(n_1014), .B2(n_1169), .Y(n_1168) );
AOI221xp5_ASAP7_75t_L g1185 ( .A1(n_8), .A2(n_280), .B1(n_833), .B2(n_1141), .C(n_1186), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_9), .A2(n_217), .B1(n_647), .B2(n_1133), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_9), .A2(n_197), .B1(n_611), .B2(n_1044), .Y(n_1143) );
AOI22xp5_ASAP7_75t_L g1536 ( .A1(n_10), .A2(n_64), .B1(n_1537), .B2(n_1539), .Y(n_1536) );
INVx1_ASAP7_75t_L g1306 ( .A(n_11), .Y(n_1306) );
OAI22xp5_ASAP7_75t_L g1324 ( .A1(n_11), .A2(n_364), .B1(n_534), .B2(n_594), .Y(n_1324) );
CKINVDCx5p33_ASAP7_75t_R g1344 ( .A(n_12), .Y(n_1344) );
A2O1A1Ixp33_ASAP7_75t_L g1240 ( .A1(n_13), .A2(n_1062), .B(n_1241), .C(n_1247), .Y(n_1240) );
AOI22xp33_ASAP7_75t_SL g1022 ( .A1(n_14), .A2(n_244), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
INVxp67_ASAP7_75t_SL g1060 ( .A(n_14), .Y(n_1060) );
INVxp67_ASAP7_75t_SL g588 ( .A(n_15), .Y(n_588) );
AND4x1_ASAP7_75t_L g658 ( .A(n_15), .B(n_590), .C(n_595), .D(n_628), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_16), .A2(n_303), .B1(n_579), .B2(n_1266), .Y(n_1265) );
AOI221xp5_ASAP7_75t_L g1270 ( .A1(n_16), .A2(n_96), .B1(n_493), .B2(n_517), .C(n_607), .Y(n_1270) );
INVx2_ASAP7_75t_L g420 ( .A(n_17), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_18), .A2(n_132), .B1(n_1081), .B2(n_1354), .Y(n_1353) );
AOI22xp33_ASAP7_75t_L g1367 ( .A1(n_18), .A2(n_183), .B1(n_705), .B2(n_1193), .Y(n_1367) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_19), .A2(n_248), .B1(n_733), .B2(n_1263), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g1271 ( .A1(n_19), .A2(n_151), .B1(n_1272), .B2(n_1274), .Y(n_1271) );
XNOR2xp5_ASAP7_75t_L g1861 ( .A(n_20), .B(n_1862), .Y(n_1861) );
INVx1_ASAP7_75t_L g993 ( .A(n_21), .Y(n_993) );
OAI22xp33_ASAP7_75t_L g1464 ( .A1(n_22), .A2(n_279), .B1(n_581), .B2(n_631), .Y(n_1464) );
INVx1_ASAP7_75t_L g1477 ( .A(n_22), .Y(n_1477) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_23), .A2(n_178), .B1(n_534), .B2(n_594), .Y(n_593) );
OAI211xp5_ASAP7_75t_L g596 ( .A1(n_23), .A2(n_524), .B(n_597), .C(n_600), .Y(n_596) );
INVx1_ASAP7_75t_L g1382 ( .A(n_24), .Y(n_1382) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_25), .A2(n_139), .B1(n_647), .B2(n_1081), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_25), .A2(n_306), .B1(n_1045), .B2(n_1106), .Y(n_1105) );
OAI22xp33_ASAP7_75t_L g1362 ( .A1(n_26), .A2(n_232), .B1(n_581), .B2(n_1087), .Y(n_1362) );
INVx1_ASAP7_75t_L g1369 ( .A(n_26), .Y(n_1369) );
AOI22xp33_ASAP7_75t_SL g1358 ( .A1(n_27), .A2(n_101), .B1(n_1026), .B2(n_1266), .Y(n_1358) );
AOI22xp33_ASAP7_75t_SL g1375 ( .A1(n_27), .A2(n_259), .B1(n_1273), .B2(n_1274), .Y(n_1375) );
AOI22xp5_ASAP7_75t_L g1561 ( .A1(n_28), .A2(n_241), .B1(n_1529), .B2(n_1534), .Y(n_1561) );
OAI22xp5_ASAP7_75t_L g1435 ( .A1(n_29), .A2(n_324), .B1(n_534), .B2(n_594), .Y(n_1435) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_30), .A2(n_103), .B1(n_609), .B2(n_611), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_30), .A2(n_42), .B1(n_645), .B2(n_647), .Y(n_649) );
CKINVDCx5p33_ASAP7_75t_R g1293 ( .A(n_31), .Y(n_1293) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_32), .Y(n_384) );
AND2x2_ASAP7_75t_L g1530 ( .A(n_32), .B(n_382), .Y(n_1530) );
AOI22xp5_ASAP7_75t_L g1528 ( .A1(n_33), .A2(n_212), .B1(n_1529), .B2(n_1534), .Y(n_1528) );
OA22x2_ASAP7_75t_L g1743 ( .A1(n_33), .A2(n_1744), .B1(n_1851), .B2(n_1852), .Y(n_1743) );
INVxp67_ASAP7_75t_L g1852 ( .A(n_33), .Y(n_1852) );
AOI22xp33_ASAP7_75t_L g1856 ( .A1(n_33), .A2(n_1857), .B1(n_1860), .B2(n_1921), .Y(n_1856) );
OAI22xp5_ASAP7_75t_SL g960 ( .A1(n_34), .A2(n_307), .B1(n_961), .B2(n_962), .Y(n_960) );
INVxp67_ASAP7_75t_SL g996 ( .A(n_34), .Y(n_996) );
CKINVDCx5p33_ASAP7_75t_R g1001 ( .A(n_35), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1429 ( .A1(n_36), .A2(n_243), .B1(n_733), .B2(n_1428), .Y(n_1429) );
AOI221xp5_ASAP7_75t_L g1448 ( .A1(n_36), .A2(n_338), .B1(n_604), .B2(n_627), .C(n_1318), .Y(n_1448) );
INVx1_ASAP7_75t_L g423 ( .A(n_37), .Y(n_423) );
OAI211xp5_ASAP7_75t_L g472 ( .A1(n_37), .A2(n_473), .B(n_481), .C(n_500), .Y(n_472) );
INVxp67_ASAP7_75t_L g1162 ( .A(n_38), .Y(n_1162) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_39), .Y(n_592) );
INVx1_ASAP7_75t_L g1785 ( .A(n_40), .Y(n_1785) );
AOI22xp5_ASAP7_75t_L g1545 ( .A1(n_41), .A2(n_290), .B1(n_1529), .B2(n_1534), .Y(n_1545) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_42), .A2(n_355), .B1(n_493), .B2(n_626), .C(n_627), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_43), .A2(n_58), .B1(n_648), .B2(n_652), .Y(n_793) );
INVx1_ASAP7_75t_L g806 ( .A(n_43), .Y(n_806) );
INVx1_ASAP7_75t_L g1424 ( .A(n_44), .Y(n_1424) );
OAI221xp5_ASAP7_75t_L g1444 ( .A1(n_44), .A2(n_264), .B1(n_507), .B2(n_614), .C(n_1445), .Y(n_1444) );
INVx1_ASAP7_75t_L g706 ( .A(n_45), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_46), .A2(n_56), .B1(n_669), .B2(n_670), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_46), .A2(n_176), .B1(n_651), .B2(n_733), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g1213 ( .A1(n_47), .A2(n_108), .B1(n_1131), .B2(n_1133), .Y(n_1213) );
AOI221xp5_ASAP7_75t_L g1242 ( .A1(n_47), .A2(n_221), .B1(n_1186), .B2(n_1243), .C(n_1244), .Y(n_1242) );
AOI221xp5_ASAP7_75t_L g516 ( .A1(n_48), .A2(n_326), .B1(n_493), .B2(n_517), .C(n_518), .Y(n_516) );
INVxp67_ASAP7_75t_SL g546 ( .A(n_48), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g1557 ( .A1(n_49), .A2(n_129), .B1(n_1529), .B2(n_1534), .Y(n_1557) );
INVx1_ASAP7_75t_L g465 ( .A(n_50), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_50), .A2(n_234), .B1(n_521), .B2(n_524), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g783 ( .A1(n_51), .A2(n_366), .B1(n_434), .B2(n_784), .C(n_785), .Y(n_783) );
AOI221xp5_ASAP7_75t_L g804 ( .A1(n_51), .A2(n_130), .B1(n_797), .B2(n_798), .C(n_805), .Y(n_804) );
AOI221xp5_ASAP7_75t_L g1506 ( .A1(n_52), .A2(n_111), .B1(n_1227), .B2(n_1507), .C(n_1508), .Y(n_1506) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_53), .A2(n_296), .B1(n_856), .B2(n_1020), .Y(n_1019) );
INVx1_ASAP7_75t_L g1051 ( .A(n_53), .Y(n_1051) );
NAND5xp2_ASAP7_75t_L g821 ( .A(n_54), .B(n_822), .C(n_851), .D(n_867), .E(n_874), .Y(n_821) );
INVx1_ASAP7_75t_L g883 ( .A(n_54), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g1555 ( .A1(n_54), .A2(n_189), .B1(n_1537), .B2(n_1556), .Y(n_1555) );
OAI22xp5_ASAP7_75t_L g1467 ( .A1(n_55), .A2(n_161), .B1(n_534), .B2(n_594), .Y(n_1467) );
OAI211xp5_ASAP7_75t_SL g1469 ( .A1(n_55), .A2(n_524), .B(n_1470), .C(n_1475), .Y(n_1469) );
AOI22xp33_ASAP7_75t_SL g719 ( .A1(n_56), .A2(n_191), .B1(n_720), .B2(n_722), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g1311 ( .A1(n_57), .A2(n_202), .B1(n_1189), .B2(n_1193), .Y(n_1311) );
AOI22xp33_ASAP7_75t_SL g1331 ( .A1(n_57), .A2(n_340), .B1(n_643), .B2(n_725), .Y(n_1331) );
INVx1_ASAP7_75t_L g800 ( .A(n_58), .Y(n_800) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_59), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_59), .A2(n_148), .B1(n_578), .B2(n_579), .Y(n_577) );
INVxp67_ASAP7_75t_L g1342 ( .A(n_60), .Y(n_1342) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_61), .Y(n_396) );
INVx1_ASAP7_75t_L g598 ( .A(n_62), .Y(n_598) );
OAI22xp33_ASAP7_75t_L g630 ( .A1(n_62), .A2(n_112), .B1(n_631), .B2(n_636), .Y(n_630) );
AOI22xp33_ASAP7_75t_SL g1128 ( .A1(n_63), .A2(n_65), .B1(n_725), .B2(n_1024), .Y(n_1128) );
INVx1_ASAP7_75t_L g1147 ( .A(n_63), .Y(n_1147) );
AOI221xp5_ASAP7_75t_L g1140 ( .A1(n_65), .A2(n_149), .B1(n_602), .B2(n_607), .C(n_1141), .Y(n_1140) );
XOR2x2_ASAP7_75t_L g1298 ( .A(n_66), .B(n_1299), .Y(n_1298) );
XOR2xp5_ASAP7_75t_L g1452 ( .A(n_67), .B(n_1453), .Y(n_1452) );
INVx1_ASAP7_75t_L g1009 ( .A(n_68), .Y(n_1009) );
INVx1_ASAP7_75t_L g1256 ( .A(n_69), .Y(n_1256) );
OAI222xp33_ASAP7_75t_L g1280 ( .A1(n_69), .A2(n_371), .B1(n_615), .B2(n_1094), .C1(n_1281), .C2(n_1286), .Y(n_1280) );
AOI22xp33_ASAP7_75t_SL g1461 ( .A1(n_70), .A2(n_302), .B1(n_1020), .B2(n_1081), .Y(n_1461) );
AOI221xp5_ASAP7_75t_L g1483 ( .A1(n_70), .A2(n_273), .B1(n_1038), .B2(n_1041), .C(n_1244), .Y(n_1483) );
AOI22xp33_ASAP7_75t_L g1494 ( .A1(n_71), .A2(n_281), .B1(n_647), .B2(n_1495), .Y(n_1494) );
AOI22xp33_ASAP7_75t_L g1509 ( .A1(n_71), .A2(n_153), .B1(n_1188), .B2(n_1234), .Y(n_1509) );
AOI22xp33_ASAP7_75t_L g1615 ( .A1(n_72), .A2(n_262), .B1(n_1537), .B2(n_1539), .Y(n_1615) );
CKINVDCx5p33_ASAP7_75t_R g1279 ( .A(n_73), .Y(n_1279) );
AOI221xp5_ASAP7_75t_L g830 ( .A1(n_74), .A2(n_187), .B1(n_479), .B2(n_493), .C(n_518), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_74), .A2(n_255), .B1(n_733), .B2(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g1396 ( .A(n_75), .Y(n_1396) );
CKINVDCx5p33_ASAP7_75t_R g1221 ( .A(n_76), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_77), .A2(n_255), .B1(n_609), .B2(n_829), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_77), .A2(n_187), .B1(n_733), .B2(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g1874 ( .A(n_78), .Y(n_1874) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_79), .A2(n_171), .B1(n_1020), .B2(n_1130), .Y(n_1172) );
AOI21xp33_ASAP7_75t_L g1195 ( .A1(n_79), .A2(n_602), .B(n_627), .Y(n_1195) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_80), .A2(n_354), .B1(n_602), .B2(n_604), .C(n_607), .Y(n_601) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_80), .A2(n_315), .B1(n_651), .B2(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g1209 ( .A(n_81), .Y(n_1209) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_82), .A2(n_351), .B1(n_672), .B2(n_675), .C(n_679), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_82), .A2(n_311), .B1(n_728), .B2(n_729), .C(n_731), .Y(n_727) );
AOI22xp33_ASAP7_75t_SL g1013 ( .A1(n_83), .A2(n_193), .B1(n_728), .B2(n_1014), .Y(n_1013) );
INVxp67_ASAP7_75t_SL g1057 ( .A(n_83), .Y(n_1057) );
AOI22xp33_ASAP7_75t_SL g1386 ( .A1(n_84), .A2(n_301), .B1(n_725), .B2(n_1026), .Y(n_1386) );
AOI22xp33_ASAP7_75t_L g1408 ( .A1(n_84), .A2(n_322), .B1(n_1188), .B2(n_1234), .Y(n_1408) );
OAI211xp5_ASAP7_75t_SL g774 ( .A1(n_85), .A2(n_742), .B(n_749), .C(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g811 ( .A(n_85), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g1895 ( .A1(n_86), .A2(n_271), .B1(n_1896), .B2(n_1898), .Y(n_1895) );
OAI22xp5_ASAP7_75t_L g1912 ( .A1(n_86), .A2(n_271), .B1(n_1913), .B2(n_1914), .Y(n_1912) );
CKINVDCx5p33_ASAP7_75t_R g1175 ( .A(n_87), .Y(n_1175) );
CKINVDCx5p33_ASAP7_75t_R g842 ( .A(n_88), .Y(n_842) );
OAI21xp5_ASAP7_75t_SL g1200 ( .A1(n_89), .A2(n_534), .B(n_1201), .Y(n_1200) );
INVxp67_ASAP7_75t_SL g712 ( .A(n_90), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_90), .A2(n_361), .B1(n_735), .B2(n_738), .Y(n_734) );
AOI22xp33_ASAP7_75t_SL g1430 ( .A1(n_91), .A2(n_367), .B1(n_725), .B2(n_1431), .Y(n_1430) );
AOI221xp5_ASAP7_75t_L g1440 ( .A1(n_91), .A2(n_156), .B1(n_497), .B2(n_833), .C(n_1099), .Y(n_1440) );
AOI22xp33_ASAP7_75t_SL g1171 ( .A1(n_92), .A2(n_280), .B1(n_642), .B2(n_1024), .Y(n_1171) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_92), .A2(n_330), .B1(n_611), .B2(n_1193), .Y(n_1192) );
AOI22xp33_ASAP7_75t_L g1498 ( .A1(n_93), .A2(n_111), .B1(n_724), .B2(n_1078), .Y(n_1498) );
INVxp67_ASAP7_75t_SL g1516 ( .A(n_93), .Y(n_1516) );
OR2x2_ASAP7_75t_L g449 ( .A(n_94), .B(n_450), .Y(n_449) );
OAI221xp5_ASAP7_75t_L g502 ( .A1(n_95), .A2(n_231), .B1(n_503), .B2(n_507), .C(n_512), .Y(n_502) );
OAI322xp33_ASAP7_75t_L g544 ( .A1(n_95), .A2(n_545), .A3(n_553), .B1(n_556), .B2(n_564), .C1(n_570), .C2(n_581), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_96), .A2(n_142), .B1(n_579), .B2(n_1263), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g1572 ( .A1(n_97), .A2(n_190), .B1(n_1529), .B2(n_1537), .Y(n_1572) );
OAI21xp5_ASAP7_75t_L g1412 ( .A1(n_98), .A2(n_534), .B(n_1413), .Y(n_1412) );
AOI22xp33_ASAP7_75t_SL g965 ( .A1(n_99), .A2(n_174), .B1(n_526), .B2(n_966), .Y(n_965) );
INVxp67_ASAP7_75t_SL g989 ( .A(n_99), .Y(n_989) );
OAI22xp33_ASAP7_75t_L g1774 ( .A1(n_100), .A2(n_209), .B1(n_1775), .B2(n_1777), .Y(n_1774) );
OAI22xp5_ASAP7_75t_L g1837 ( .A1(n_100), .A2(n_209), .B1(n_1838), .B2(n_1842), .Y(n_1837) );
AOI221xp5_ASAP7_75t_L g1366 ( .A1(n_101), .A2(n_336), .B1(n_493), .B2(n_498), .C(n_1318), .Y(n_1366) );
INVx1_ASAP7_75t_L g1065 ( .A(n_102), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_103), .A2(n_355), .B1(n_645), .B2(n_647), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g1571 ( .A1(n_104), .A2(n_317), .B1(n_1534), .B2(n_1539), .Y(n_1571) );
AOI22xp5_ASAP7_75t_L g1547 ( .A1(n_105), .A2(n_168), .B1(n_1537), .B2(n_1548), .Y(n_1547) );
OAI21xp33_ASAP7_75t_L g1289 ( .A1(n_106), .A2(n_1290), .B(n_1291), .Y(n_1289) );
INVx1_ASAP7_75t_L g1804 ( .A(n_107), .Y(n_1804) );
AOI22xp33_ASAP7_75t_SL g1232 ( .A1(n_108), .A2(n_145), .B1(n_1233), .B2(n_1234), .Y(n_1232) );
INVx1_ASAP7_75t_L g1873 ( .A(n_109), .Y(n_1873) );
CKINVDCx5p33_ASAP7_75t_R g1183 ( .A(n_110), .Y(n_1183) );
INVx1_ASAP7_75t_L g599 ( .A(n_112), .Y(n_599) );
OAI211xp5_ASAP7_75t_L g835 ( .A1(n_113), .A2(n_836), .B(n_838), .C(n_840), .Y(n_835) );
INVx1_ASAP7_75t_L g879 ( .A(n_113), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g1387 ( .A1(n_114), .A2(n_332), .B1(n_1354), .B2(n_1388), .Y(n_1387) );
AOI221xp5_ASAP7_75t_L g1409 ( .A1(n_114), .A2(n_358), .B1(n_1108), .B2(n_1229), .C(n_1410), .Y(n_1409) );
INVx1_ASAP7_75t_L g1123 ( .A(n_115), .Y(n_1123) );
OAI221xp5_ASAP7_75t_L g1145 ( .A1(n_115), .A2(n_150), .B1(n_507), .B2(n_614), .C(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_L g513 ( .A(n_116), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g1616 ( .A1(n_117), .A2(n_348), .B1(n_1529), .B2(n_1534), .Y(n_1616) );
CKINVDCx5p33_ASAP7_75t_R g1178 ( .A(n_118), .Y(n_1178) );
OAI22xp5_ASAP7_75t_L g1196 ( .A1(n_118), .A2(n_133), .B1(n_1197), .B2(n_1198), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_119), .A2(n_254), .B1(n_526), .B2(n_828), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_119), .A2(n_274), .B1(n_642), .B2(n_724), .Y(n_985) );
INVx1_ASAP7_75t_L g1882 ( .A(n_120), .Y(n_1882) );
INVx1_ASAP7_75t_L g1807 ( .A(n_121), .Y(n_1807) );
AOI22xp33_ASAP7_75t_L g1393 ( .A1(n_122), .A2(n_322), .B1(n_724), .B2(n_725), .Y(n_1393) );
AOI221xp5_ASAP7_75t_L g1404 ( .A1(n_122), .A2(n_301), .B1(n_497), .B2(n_498), .C(n_1405), .Y(n_1404) );
INVx1_ASAP7_75t_L g951 ( .A(n_123), .Y(n_951) );
INVx1_ASAP7_75t_L g1126 ( .A(n_124), .Y(n_1126) );
OAI221xp5_ASAP7_75t_L g613 ( .A1(n_125), .A2(n_287), .B1(n_614), .B2(n_615), .C(n_617), .Y(n_613) );
INVx1_ASAP7_75t_L g657 ( .A(n_125), .Y(n_657) );
INVx1_ASAP7_75t_L g382 ( .A(n_126), .Y(n_382) );
AOI22xp33_ASAP7_75t_SL g1463 ( .A1(n_127), .A2(n_300), .B1(n_725), .B2(n_1026), .Y(n_1463) );
INVxp67_ASAP7_75t_SL g1482 ( .A(n_127), .Y(n_1482) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_128), .A2(n_200), .B1(n_856), .B2(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g1055 ( .A(n_128), .Y(n_1055) );
INVx1_ASAP7_75t_L g790 ( .A(n_130), .Y(n_790) );
OAI222xp33_ASAP7_75t_L g913 ( .A1(n_131), .A2(n_350), .B1(n_745), .B2(n_747), .C1(n_914), .C2(n_916), .Y(n_913) );
INVx1_ASAP7_75t_L g926 ( .A(n_131), .Y(n_926) );
AOI21xp33_ASAP7_75t_L g1374 ( .A1(n_132), .A2(n_518), .B(n_606), .Y(n_1374) );
CKINVDCx5p33_ASAP7_75t_R g1177 ( .A(n_133), .Y(n_1177) );
INVx1_ASAP7_75t_L g1491 ( .A(n_134), .Y(n_1491) );
OAI221xp5_ASAP7_75t_L g1513 ( .A1(n_134), .A2(n_135), .B1(n_507), .B2(n_614), .C(n_1514), .Y(n_1513) );
INVx1_ASAP7_75t_L g1490 ( .A(n_135), .Y(n_1490) );
INVx1_ASAP7_75t_L g903 ( .A(n_136), .Y(n_903) );
OAI211xp5_ASAP7_75t_L g954 ( .A1(n_137), .A2(n_955), .B(n_956), .C(n_957), .Y(n_954) );
INVxp33_ASAP7_75t_SL g977 ( .A(n_137), .Y(n_977) );
OAI22xp33_ASAP7_75t_L g752 ( .A1(n_138), .A2(n_184), .B1(n_753), .B2(n_756), .Y(n_752) );
INVxp67_ASAP7_75t_SL g761 ( .A(n_138), .Y(n_761) );
AOI221xp5_ASAP7_75t_L g1098 ( .A1(n_139), .A2(n_258), .B1(n_517), .B2(n_627), .C(n_1099), .Y(n_1098) );
INVxp67_ASAP7_75t_SL g1314 ( .A(n_140), .Y(n_1314) );
AOI22xp33_ASAP7_75t_L g1332 ( .A1(n_140), .A2(n_276), .B1(n_1333), .B2(n_1334), .Y(n_1332) );
AOI22xp33_ASAP7_75t_SL g1544 ( .A1(n_141), .A2(n_235), .B1(n_1537), .B2(n_1539), .Y(n_1544) );
INVx1_ASAP7_75t_L g1284 ( .A(n_142), .Y(n_1284) );
INVx1_ASAP7_75t_L g1005 ( .A(n_143), .Y(n_1005) );
OAI222xp33_ASAP7_75t_L g1049 ( .A1(n_143), .A2(n_228), .B1(n_473), .B2(n_615), .C1(n_1050), .C2(n_1056), .Y(n_1049) );
INVx1_ASAP7_75t_L g1305 ( .A(n_144), .Y(n_1305) );
OAI22xp33_ASAP7_75t_L g1339 ( .A1(n_144), .A2(n_195), .B1(n_636), .B2(n_1087), .Y(n_1339) );
AOI22xp33_ASAP7_75t_L g1214 ( .A1(n_145), .A2(n_221), .B1(n_1131), .B2(n_1215), .Y(n_1214) );
XOR2x2_ASAP7_75t_L g1069 ( .A(n_146), .B(n_1070), .Y(n_1069) );
INVxp67_ASAP7_75t_SL g1309 ( .A(n_147), .Y(n_1309) );
AOI22xp33_ASAP7_75t_SL g1335 ( .A1(n_147), .A2(n_220), .B1(n_647), .B2(n_1336), .Y(n_1335) );
AOI221xp5_ASAP7_75t_L g492 ( .A1(n_148), .A2(n_242), .B1(n_493), .B2(n_497), .C(n_498), .Y(n_492) );
AOI22xp33_ASAP7_75t_SL g1135 ( .A1(n_149), .A2(n_154), .B1(n_1026), .B2(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1122 ( .A(n_150), .Y(n_1122) );
AOI22xp33_ASAP7_75t_SL g1261 ( .A1(n_151), .A2(n_250), .B1(n_733), .B2(n_1023), .Y(n_1261) );
OAI22xp33_ASAP7_75t_L g773 ( .A1(n_152), .A2(n_370), .B1(n_753), .B2(n_756), .Y(n_773) );
INVxp33_ASAP7_75t_SL g815 ( .A(n_152), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g1497 ( .A1(n_153), .A2(n_192), .B1(n_647), .B2(n_1495), .Y(n_1497) );
INVxp67_ASAP7_75t_SL g1148 ( .A(n_154), .Y(n_1148) );
CKINVDCx5p33_ASAP7_75t_R g776 ( .A(n_155), .Y(n_776) );
AOI22xp33_ASAP7_75t_SL g1426 ( .A1(n_156), .A2(n_206), .B1(n_724), .B2(n_725), .Y(n_1426) );
INVx1_ASAP7_75t_L g780 ( .A(n_157), .Y(n_780) );
AOI221xp5_ASAP7_75t_L g796 ( .A1(n_157), .A2(n_266), .B1(n_797), .B2(n_798), .C(n_799), .Y(n_796) );
AOI22xp33_ASAP7_75t_SL g1077 ( .A1(n_158), .A2(n_185), .B1(n_1026), .B2(n_1078), .Y(n_1077) );
AOI221xp5_ASAP7_75t_L g1107 ( .A1(n_158), .A2(n_207), .B1(n_498), .B2(n_1041), .C(n_1108), .Y(n_1107) );
OAI22xp33_ASAP7_75t_L g1086 ( .A1(n_159), .A2(n_316), .B1(n_581), .B2(n_1087), .Y(n_1086) );
INVx1_ASAP7_75t_L g1112 ( .A(n_159), .Y(n_1112) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_160), .A2(n_176), .B1(n_670), .B2(n_691), .C(n_692), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_160), .A2(n_351), .B1(n_724), .B2(n_725), .C(n_726), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g1427 ( .A1(n_162), .A2(n_338), .B1(n_1334), .B2(n_1428), .Y(n_1427) );
AOI22xp33_ASAP7_75t_L g1439 ( .A1(n_162), .A2(n_243), .B1(n_1044), .B2(n_1189), .Y(n_1439) );
OAI22xp33_ASAP7_75t_L g1499 ( .A1(n_163), .A2(n_295), .B1(n_581), .B2(n_631), .Y(n_1499) );
INVx1_ASAP7_75t_L g1512 ( .A(n_163), .Y(n_1512) );
INVx1_ASAP7_75t_L g1030 ( .A(n_164), .Y(n_1030) );
INVx1_ASAP7_75t_L g1347 ( .A(n_165), .Y(n_1347) );
OAI221xp5_ASAP7_75t_SL g1371 ( .A1(n_165), .A2(n_277), .B1(n_614), .B2(n_615), .C(n_1372), .Y(n_1371) );
CKINVDCx5p33_ASAP7_75t_R g1434 ( .A(n_166), .Y(n_1434) );
OAI22xp33_ASAP7_75t_L g1903 ( .A1(n_167), .A2(n_177), .B1(n_1904), .B2(n_1906), .Y(n_1903) );
OAI22xp33_ASAP7_75t_L g1909 ( .A1(n_167), .A2(n_177), .B1(n_1910), .B2(n_1911), .Y(n_1909) );
INVx1_ASAP7_75t_L g1294 ( .A(n_168), .Y(n_1294) );
AO22x1_ASAP7_75t_L g1166 ( .A1(n_169), .A2(n_219), .B1(n_1130), .B2(n_1131), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_169), .B(n_1099), .Y(n_1191) );
INVx1_ASAP7_75t_L g873 ( .A(n_170), .Y(n_873) );
AOI22xp33_ASAP7_75t_SL g1187 ( .A1(n_171), .A2(n_219), .B1(n_1188), .B2(n_1189), .Y(n_1187) );
CKINVDCx5p33_ASAP7_75t_R g1090 ( .A(n_172), .Y(n_1090) );
INVx1_ASAP7_75t_L g1901 ( .A(n_173), .Y(n_1901) );
INVx1_ASAP7_75t_L g984 ( .A(n_174), .Y(n_984) );
CKINVDCx5p33_ASAP7_75t_R g1466 ( .A(n_175), .Y(n_1466) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_179), .A2(n_359), .B1(n_534), .B2(n_594), .Y(n_1091) );
INVx1_ASAP7_75t_L g1879 ( .A(n_180), .Y(n_1879) );
OAI22xp5_ASAP7_75t_L g1119 ( .A1(n_181), .A2(n_305), .B1(n_534), .B2(n_594), .Y(n_1119) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_182), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g1355 ( .A1(n_183), .A2(n_328), .B1(n_1354), .B2(n_1356), .Y(n_1355) );
INVxp67_ASAP7_75t_SL g701 ( .A(n_184), .Y(n_701) );
INVxp67_ASAP7_75t_SL g1096 ( .A(n_185), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g1502 ( .A1(n_186), .A2(n_205), .B1(n_534), .B2(n_594), .Y(n_1502) );
OAI211xp5_ASAP7_75t_L g1504 ( .A1(n_186), .A2(n_1103), .B(n_1505), .C(n_1510), .Y(n_1504) );
INVx1_ASAP7_75t_L g900 ( .A(n_188), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_188), .A2(n_282), .B1(n_609), .B2(n_829), .Y(n_934) );
INVx1_ASAP7_75t_L g1415 ( .A(n_190), .Y(n_1415) );
INVx1_ASAP7_75t_L g693 ( .A(n_191), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g1517 ( .A1(n_192), .A2(n_281), .B1(n_517), .B2(n_627), .C(n_1518), .Y(n_1517) );
AOI221xp5_ASAP7_75t_L g1037 ( .A1(n_193), .A2(n_244), .B1(n_607), .B2(n_1038), .C(n_1041), .Y(n_1037) );
CKINVDCx5p33_ASAP7_75t_R g958 ( .A(n_194), .Y(n_958) );
INVx1_ASAP7_75t_L g1303 ( .A(n_195), .Y(n_1303) );
INVx1_ASAP7_75t_L g969 ( .A(n_196), .Y(n_969) );
AOI22xp33_ASAP7_75t_SL g1129 ( .A1(n_197), .A2(n_288), .B1(n_1130), .B2(n_1131), .Y(n_1129) );
OAI211xp5_ASAP7_75t_L g823 ( .A1(n_198), .A2(n_824), .B(n_826), .C(n_834), .Y(n_823) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_198), .B(n_438), .Y(n_850) );
XNOR2x2_ASAP7_75t_L g1418 ( .A(n_199), .B(n_1419), .Y(n_1418) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_200), .A2(n_296), .B1(n_1044), .B2(n_1045), .Y(n_1043) );
INVx1_ASAP7_75t_L g1075 ( .A(n_201), .Y(n_1075) );
OAI221xp5_ASAP7_75t_L g1093 ( .A1(n_201), .A2(n_333), .B1(n_507), .B2(n_1094), .C(n_1095), .Y(n_1093) );
AOI22xp33_ASAP7_75t_SL g1338 ( .A1(n_202), .A2(n_368), .B1(n_653), .B2(n_725), .Y(n_1338) );
INVx2_ASAP7_75t_L g1532 ( .A(n_203), .Y(n_1532) );
AND2x2_ASAP7_75t_L g1535 ( .A(n_203), .B(n_1533), .Y(n_1535) );
AND2x2_ASAP7_75t_L g1540 ( .A(n_203), .B(n_314), .Y(n_1540) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_204), .Y(n_543) );
INVxp67_ASAP7_75t_SL g1446 ( .A(n_206), .Y(n_1446) );
AOI22xp33_ASAP7_75t_SL g1085 ( .A1(n_207), .A2(n_309), .B1(n_642), .B2(n_724), .Y(n_1085) );
INVx1_ASAP7_75t_L g1402 ( .A(n_208), .Y(n_1402) );
OAI22xp5_ASAP7_75t_L g1222 ( .A1(n_210), .A2(n_297), .B1(n_438), .B2(n_534), .Y(n_1222) );
OAI211xp5_ASAP7_75t_L g1224 ( .A1(n_210), .A2(n_524), .B(n_1225), .C(n_1235), .Y(n_1224) );
AOI22xp5_ASAP7_75t_L g1563 ( .A1(n_211), .A2(n_269), .B1(n_1534), .B2(n_1537), .Y(n_1563) );
CKINVDCx5p33_ASAP7_75t_R g1182 ( .A(n_213), .Y(n_1182) );
XOR2x2_ASAP7_75t_L g1485 ( .A(n_214), .B(n_1486), .Y(n_1485) );
OAI22xp33_ASAP7_75t_L g1432 ( .A1(n_215), .A2(n_283), .B1(n_581), .B2(n_1087), .Y(n_1432) );
INVx1_ASAP7_75t_L g1442 ( .A(n_215), .Y(n_1442) );
AOI22xp33_ASAP7_75t_L g1390 ( .A1(n_216), .A2(n_358), .B1(n_647), .B2(n_1388), .Y(n_1390) );
AOI22xp33_ASAP7_75t_L g1406 ( .A1(n_216), .A2(n_332), .B1(n_1233), .B2(n_1234), .Y(n_1406) );
AOI221xp5_ASAP7_75t_L g1149 ( .A1(n_217), .A2(n_288), .B1(n_493), .B2(n_518), .C(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g1361 ( .A(n_218), .Y(n_1361) );
INVxp67_ASAP7_75t_SL g1316 ( .A(n_220), .Y(n_1316) );
INVx1_ASAP7_75t_L g941 ( .A(n_222), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g1564 ( .A1(n_223), .A2(n_227), .B1(n_1529), .B2(n_1548), .Y(n_1564) );
NOR2xp33_ASAP7_75t_L g1319 ( .A(n_224), .B(n_1094), .Y(n_1319) );
INVx1_ASAP7_75t_L g1329 ( .A(n_224), .Y(n_1329) );
INVx1_ASAP7_75t_L g1029 ( .A(n_225), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_226), .A2(n_293), .B1(n_828), .B2(n_829), .Y(n_827) );
AOI22xp33_ASAP7_75t_SL g859 ( .A1(n_226), .A2(n_313), .B1(n_725), .B2(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g1006 ( .A(n_228), .Y(n_1006) );
INVx1_ASAP7_75t_L g1259 ( .A(n_229), .Y(n_1259) );
OAI211xp5_ASAP7_75t_L g1268 ( .A1(n_229), .A2(n_1103), .B(n_1269), .C(n_1276), .Y(n_1268) );
OAI211xp5_ASAP7_75t_L g1899 ( .A1(n_230), .A2(n_1762), .B(n_1891), .C(n_1900), .Y(n_1899) );
INVx1_ASAP7_75t_L g1920 ( .A(n_230), .Y(n_1920) );
INVx1_ASAP7_75t_L g409 ( .A(n_231), .Y(n_409) );
INVx1_ASAP7_75t_L g1370 ( .A(n_232), .Y(n_1370) );
CKINVDCx5p33_ASAP7_75t_R g902 ( .A(n_233), .Y(n_902) );
INVx1_ASAP7_75t_L g436 ( .A(n_234), .Y(n_436) );
INVx1_ASAP7_75t_L g584 ( .A(n_235), .Y(n_584) );
CKINVDCx5p33_ASAP7_75t_R g845 ( .A(n_236), .Y(n_845) );
INVx2_ASAP7_75t_L g422 ( .A(n_237), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_237), .B(n_420), .Y(n_457) );
INVx1_ASAP7_75t_L g569 ( .A(n_237), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g1277 ( .A(n_238), .Y(n_1277) );
AOI22xp5_ASAP7_75t_L g1549 ( .A1(n_239), .A2(n_362), .B1(n_1529), .B2(n_1534), .Y(n_1549) );
INVx1_ASAP7_75t_L g911 ( .A(n_240), .Y(n_911) );
NAND2xp33_ASAP7_75t_SL g935 ( .A(n_240), .B(n_479), .Y(n_935) );
INVx1_ASAP7_75t_L g561 ( .A(n_242), .Y(n_561) );
INVx1_ASAP7_75t_L g1881 ( .A(n_245), .Y(n_1881) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_246), .A2(n_321), .B1(n_836), .B2(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g877 ( .A(n_246), .Y(n_877) );
INVx1_ASAP7_75t_L g491 ( .A(n_247), .Y(n_491) );
INVx1_ASAP7_75t_L g1283 ( .A(n_248), .Y(n_1283) );
INVx1_ASAP7_75t_L g1794 ( .A(n_249), .Y(n_1794) );
INVx1_ASAP7_75t_L g1287 ( .A(n_250), .Y(n_1287) );
AOI21xp5_ASAP7_75t_L g912 ( .A1(n_251), .A2(n_652), .B(n_726), .Y(n_912) );
INVx1_ASAP7_75t_L g937 ( .A(n_252), .Y(n_937) );
BUFx3_ASAP7_75t_L g414 ( .A(n_253), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_254), .A2(n_289), .B1(n_724), .B2(n_991), .Y(n_990) );
CKINVDCx20_ASAP7_75t_R g1395 ( .A(n_256), .Y(n_1395) );
CKINVDCx5p33_ASAP7_75t_R g777 ( .A(n_257), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_258), .A2(n_306), .B1(n_573), .B2(n_647), .Y(n_1083) );
AOI22xp33_ASAP7_75t_SL g1352 ( .A1(n_259), .A2(n_336), .B1(n_1024), .B2(n_1266), .Y(n_1352) );
INVx1_ASAP7_75t_L g893 ( .A(n_260), .Y(n_893) );
NOR2xp33_ASAP7_75t_L g895 ( .A(n_260), .B(n_753), .Y(n_895) );
OAI211xp5_ASAP7_75t_SL g1759 ( .A1(n_261), .A2(n_1760), .B(n_1762), .C(n_1764), .Y(n_1759) );
INVx1_ASAP7_75t_L g1833 ( .A(n_261), .Y(n_1833) );
AOI21xp33_ASAP7_75t_L g972 ( .A1(n_263), .A2(n_518), .B(n_798), .Y(n_972) );
INVx1_ASAP7_75t_L g983 ( .A(n_263), .Y(n_983) );
INVx1_ASAP7_75t_L g1423 ( .A(n_264), .Y(n_1423) );
INVx1_ASAP7_75t_L g1400 ( .A(n_265), .Y(n_1400) );
AOI21xp33_ASAP7_75t_L g792 ( .A1(n_266), .A2(n_573), .B(n_731), .Y(n_792) );
XOR2x2_ASAP7_75t_L g946 ( .A(n_267), .B(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g1773 ( .A(n_268), .Y(n_1773) );
OAI211xp5_ASAP7_75t_SL g1823 ( .A1(n_268), .A2(n_1824), .B(n_1826), .C(n_1829), .Y(n_1823) );
OAI22xp33_ASAP7_75t_L g1218 ( .A1(n_270), .A2(n_285), .B1(n_581), .B2(n_631), .Y(n_1218) );
INVx1_ASAP7_75t_L g1236 ( .A(n_270), .Y(n_1236) );
BUFx3_ASAP7_75t_L g399 ( .A(n_272), .Y(n_399) );
INVx1_ASAP7_75t_L g478 ( .A(n_272), .Y(n_478) );
AOI22xp33_ASAP7_75t_SL g1462 ( .A1(n_273), .A2(n_325), .B1(n_1020), .B2(n_1081), .Y(n_1462) );
NAND2xp5_ASAP7_75t_SL g964 ( .A(n_274), .B(n_798), .Y(n_964) );
INVxp67_ASAP7_75t_SL g1350 ( .A(n_275), .Y(n_1350) );
OAI211xp5_ASAP7_75t_SL g1364 ( .A1(n_275), .A2(n_524), .B(n_1365), .C(n_1368), .Y(n_1364) );
AOI21xp5_ASAP7_75t_L g1312 ( .A1(n_276), .A2(n_518), .B(n_1141), .Y(n_1312) );
INVx1_ASAP7_75t_L g1348 ( .A(n_277), .Y(n_1348) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_278), .Y(n_782) );
INVx1_ASAP7_75t_L g1476 ( .A(n_279), .Y(n_1476) );
INVx1_ASAP7_75t_L g909 ( .A(n_282), .Y(n_909) );
INVx1_ASAP7_75t_L g1443 ( .A(n_283), .Y(n_1443) );
INVx1_ASAP7_75t_L g1210 ( .A(n_284), .Y(n_1210) );
INVx1_ASAP7_75t_L g1237 ( .A(n_285), .Y(n_1237) );
INVx1_ASAP7_75t_L g484 ( .A(n_286), .Y(n_484) );
INVx1_ASAP7_75t_L g655 ( .A(n_287), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g967 ( .A(n_289), .B(n_497), .Y(n_967) );
INVx1_ASAP7_75t_L g764 ( .A(n_291), .Y(n_764) );
XNOR2x2_ASAP7_75t_L g1204 ( .A(n_292), .B(n_1205), .Y(n_1204) );
AOI22xp33_ASAP7_75t_SL g853 ( .A1(n_293), .A2(n_372), .B1(n_725), .B2(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g430 ( .A(n_294), .Y(n_430) );
INVx1_ASAP7_75t_L g444 ( .A(n_294), .Y(n_444) );
INVx1_ASAP7_75t_L g1511 ( .A(n_295), .Y(n_1511) );
CKINVDCx5p33_ASAP7_75t_R g1118 ( .A(n_298), .Y(n_1118) );
INVx1_ASAP7_75t_L g1797 ( .A(n_299), .Y(n_1797) );
AOI221xp5_ASAP7_75t_L g1471 ( .A1(n_300), .A2(n_331), .B1(n_607), .B2(n_1405), .C(n_1472), .Y(n_1471) );
AOI22xp33_ASAP7_75t_L g1474 ( .A1(n_302), .A2(n_325), .B1(n_1233), .B2(n_1234), .Y(n_1474) );
INVx1_ASAP7_75t_L g1288 ( .A(n_303), .Y(n_1288) );
INVx1_ASAP7_75t_L g1798 ( .A(n_304), .Y(n_1798) );
OAI211xp5_ASAP7_75t_L g1138 ( .A1(n_305), .A2(n_1103), .B(n_1139), .C(n_1144), .Y(n_1138) );
OAI21xp33_ASAP7_75t_L g975 ( .A1(n_307), .A2(n_869), .B(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g1790 ( .A(n_308), .Y(n_1790) );
INVxp67_ASAP7_75t_SL g1097 ( .A(n_309), .Y(n_1097) );
AOI22xp5_ASAP7_75t_SL g1560 ( .A1(n_310), .A2(n_369), .B1(n_1537), .B2(n_1548), .Y(n_1560) );
INVx1_ASAP7_75t_L g694 ( .A(n_311), .Y(n_694) );
CKINVDCx5p33_ASAP7_75t_R g892 ( .A(n_312), .Y(n_892) );
AOI221xp5_ASAP7_75t_SL g832 ( .A1(n_313), .A2(n_372), .B1(n_479), .B2(n_606), .C(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g1533 ( .A(n_314), .Y(n_1533) );
AND2x2_ASAP7_75t_L g1538 ( .A(n_314), .B(n_1532), .Y(n_1538) );
INVxp67_ASAP7_75t_SL g624 ( .A(n_315), .Y(n_624) );
INVx1_ASAP7_75t_L g1113 ( .A(n_316), .Y(n_1113) );
INVx1_ASAP7_75t_L g1902 ( .A(n_318), .Y(n_1902) );
OAI211xp5_ASAP7_75t_L g1918 ( .A1(n_318), .A2(n_1795), .B(n_1826), .C(n_1919), .Y(n_1918) );
OAI211xp5_ASAP7_75t_SL g1307 ( .A1(n_319), .A2(n_507), .B(n_1308), .C(n_1313), .Y(n_1307) );
INVx1_ASAP7_75t_L g1328 ( .A(n_319), .Y(n_1328) );
OAI22xp33_ASAP7_75t_L g1752 ( .A1(n_320), .A2(n_375), .B1(n_1753), .B2(n_1756), .Y(n_1752) );
OAI22xp33_ASAP7_75t_L g1845 ( .A1(n_320), .A2(n_375), .B1(n_391), .B2(n_1846), .Y(n_1845) );
INVx1_ASAP7_75t_L g866 ( .A(n_321), .Y(n_866) );
XNOR2xp5_ASAP7_75t_L g765 ( .A(n_323), .B(n_766), .Y(n_765) );
OAI211xp5_ASAP7_75t_L g1437 ( .A1(n_324), .A2(n_524), .B(n_1438), .C(n_1441), .Y(n_1437) );
INVxp67_ASAP7_75t_SL g574 ( .A(n_326), .Y(n_574) );
INVx1_ASAP7_75t_L g1868 ( .A(n_327), .Y(n_1868) );
INVx1_ASAP7_75t_L g1373 ( .A(n_328), .Y(n_1373) );
CKINVDCx16_ASAP7_75t_R g915 ( .A(n_329), .Y(n_915) );
INVx1_ASAP7_75t_L g1074 ( .A(n_333), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_334), .B(n_1246), .Y(n_1245) );
OAI21xp33_ASAP7_75t_L g1027 ( .A1(n_335), .A2(n_534), .B(n_1028), .Y(n_1027) );
INVx1_ASAP7_75t_L g768 ( .A(n_337), .Y(n_768) );
INVx1_ASAP7_75t_L g788 ( .A(n_339), .Y(n_788) );
AOI221xp5_ASAP7_75t_L g1317 ( .A1(n_340), .A2(n_368), .B1(n_498), .B2(n_604), .C(n_1318), .Y(n_1317) );
INVx1_ASAP7_75t_L g1878 ( .A(n_341), .Y(n_1878) );
INVx1_ASAP7_75t_L g1869 ( .A(n_342), .Y(n_1869) );
INVx1_ASAP7_75t_L g1769 ( .A(n_343), .Y(n_1769) );
CKINVDCx5p33_ASAP7_75t_R g1203 ( .A(n_344), .Y(n_1203) );
CKINVDCx5p33_ASAP7_75t_R g1383 ( .A(n_345), .Y(n_1383) );
INVxp67_ASAP7_75t_SL g620 ( .A(n_346), .Y(n_620) );
AOI22xp33_ASAP7_75t_SL g641 ( .A1(n_346), .A2(n_354), .B1(n_642), .B2(n_643), .Y(n_641) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_347), .Y(n_395) );
INVx1_ASAP7_75t_L g1323 ( .A(n_349), .Y(n_1323) );
NOR2xp33_ASAP7_75t_R g928 ( .A(n_350), .B(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g888 ( .A(n_352), .Y(n_888) );
INVx1_ASAP7_75t_L g1457 ( .A(n_353), .Y(n_1457) );
OAI221xp5_ASAP7_75t_SL g1478 ( .A1(n_353), .A2(n_374), .B1(n_614), .B2(n_615), .C(n_1479), .Y(n_1478) );
INVxp67_ASAP7_75t_SL g710 ( .A(n_356), .Y(n_710) );
OAI221xp5_ASAP7_75t_L g744 ( .A1(n_356), .A2(n_357), .B1(n_745), .B2(n_747), .C(n_749), .Y(n_744) );
OAI221xp5_ASAP7_75t_L g681 ( .A1(n_357), .A2(n_361), .B1(n_682), .B2(n_687), .C(n_688), .Y(n_681) );
OAI211xp5_ASAP7_75t_L g1102 ( .A1(n_359), .A2(n_1103), .B(n_1104), .C(n_1111), .Y(n_1102) );
XOR2x2_ASAP7_75t_L g1115 ( .A(n_360), .B(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g417 ( .A(n_363), .Y(n_417) );
INVx1_ASAP7_75t_L g448 ( .A(n_363), .Y(n_448) );
INVx2_ASAP7_75t_L g531 ( .A(n_363), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g1501 ( .A(n_365), .Y(n_1501) );
INVx1_ASAP7_75t_L g801 ( .A(n_366), .Y(n_801) );
INVxp67_ASAP7_75t_SL g1447 ( .A(n_367), .Y(n_1447) );
INVxp67_ASAP7_75t_SL g771 ( .A(n_370), .Y(n_771) );
INVx1_ASAP7_75t_L g1255 ( .A(n_371), .Y(n_1255) );
INVx1_ASAP7_75t_L g1792 ( .A(n_373), .Y(n_1792) );
INVx1_ASAP7_75t_L g1458 ( .A(n_374), .Y(n_1458) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_400), .B(n_1521), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_385), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g1855 ( .A(n_379), .B(n_388), .Y(n_1855) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g1859 ( .A(n_381), .B(n_384), .Y(n_1859) );
INVx1_ASAP7_75t_L g1924 ( .A(n_381), .Y(n_1924) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g1926 ( .A(n_384), .B(n_1924), .Y(n_1926) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g1849 ( .A(n_388), .B(n_1850), .Y(n_1849) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g499 ( .A(n_389), .B(n_399), .Y(n_499) );
AND2x4_ASAP7_75t_L g519 ( .A(n_389), .B(n_398), .Y(n_519) );
AND2x4_ASAP7_75t_SL g1854 ( .A(n_390), .B(n_1855), .Y(n_1854) );
INVx1_ASAP7_75t_L g1910 ( .A(n_390), .Y(n_1910) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x6_ASAP7_75t_L g391 ( .A(n_392), .B(n_397), .Y(n_391) );
INVxp67_ASAP7_75t_L g1246 ( .A(n_392), .Y(n_1246) );
INVx1_ASAP7_75t_L g1789 ( .A(n_392), .Y(n_1789) );
OR2x6_ASAP7_75t_L g1840 ( .A(n_392), .B(n_1841), .Y(n_1840) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g483 ( .A(n_393), .Y(n_483) );
BUFx4f_ASAP7_75t_L g837 ( .A(n_393), .Y(n_837) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx2_ASAP7_75t_L g462 ( .A(n_395), .Y(n_462) );
AND2x2_ASAP7_75t_L g480 ( .A(n_395), .B(n_396), .Y(n_480) );
INVx2_ASAP7_75t_L g490 ( .A(n_395), .Y(n_490) );
AND2x2_ASAP7_75t_L g495 ( .A(n_395), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g538 ( .A(n_395), .Y(n_538) );
NAND2x1_ASAP7_75t_L g678 ( .A(n_395), .B(n_396), .Y(n_678) );
INVx1_ASAP7_75t_L g463 ( .A(n_396), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_396), .B(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g496 ( .A(n_396), .Y(n_496) );
BUFx2_ASAP7_75t_L g510 ( .A(n_396), .Y(n_510) );
AND2x2_ASAP7_75t_L g527 ( .A(n_396), .B(n_490), .Y(n_527) );
OR2x2_ASAP7_75t_L g674 ( .A(n_396), .B(n_462), .Y(n_674) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g1828 ( .A(n_398), .Y(n_1828) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_L g1832 ( .A(n_399), .Y(n_1832) );
AND2x4_ASAP7_75t_L g1836 ( .A(n_399), .B(n_537), .Y(n_1836) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_1154), .B2(n_1155), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
XNOR2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_659), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_585), .B2(n_586), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
XNOR2x1_ASAP7_75t_L g405 ( .A(n_406), .B(n_584), .Y(n_405) );
NOR2x1_ASAP7_75t_L g406 ( .A(n_407), .B(n_470), .Y(n_406) );
NAND5xp2_ASAP7_75t_L g407 ( .A(n_408), .B(n_431), .C(n_435), .D(n_449), .E(n_464), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_423), .B2(n_424), .Y(n_408) );
AO22x1_ASAP7_75t_L g1004 ( .A1(n_410), .A2(n_424), .B1(n_1005), .B2(n_1006), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1176 ( .A1(n_410), .A2(n_424), .B1(n_1177), .B2(n_1178), .Y(n_1176) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_410), .A2(n_424), .B1(n_1209), .B2(n_1210), .Y(n_1208) );
AOI22xp33_ASAP7_75t_L g1456 ( .A1(n_410), .A2(n_424), .B1(n_1457), .B2(n_1458), .Y(n_1456) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_415), .Y(n_410) );
AND2x2_ASAP7_75t_L g656 ( .A(n_411), .B(n_415), .Y(n_656) );
AND2x6_ASAP7_75t_L g746 ( .A(n_411), .B(n_418), .Y(n_746) );
AND2x4_ASAP7_75t_SL g864 ( .A(n_411), .B(n_415), .Y(n_864) );
NAND2x1_ASAP7_75t_L g980 ( .A(n_411), .B(n_415), .Y(n_980) );
INVx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2x1p5_ASAP7_75t_L g541 ( .A(n_413), .B(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g648 ( .A(n_413), .B(n_428), .Y(n_648) );
BUFx2_ASAP7_75t_L g1768 ( .A(n_413), .Y(n_1768) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g434 ( .A(n_414), .B(n_429), .Y(n_434) );
INVx2_ASAP7_75t_L g441 ( .A(n_414), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_414), .B(n_430), .Y(n_454) );
OR2x2_ASAP7_75t_L g560 ( .A(n_414), .B(n_443), .Y(n_560) );
AND2x4_ASAP7_75t_L g424 ( .A(n_415), .B(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_L g432 ( .A(n_415), .B(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_SL g865 ( .A(n_415), .B(n_425), .Y(n_865) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
OR2x2_ASAP7_75t_L g458 ( .A(n_416), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g699 ( .A(n_416), .Y(n_699) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g568 ( .A(n_417), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_417), .B(n_477), .Y(n_704) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_418), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g748 ( .A(n_418), .B(n_427), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_418), .Y(n_751) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
NAND3x1_ASAP7_75t_L g567 ( .A(n_419), .B(n_568), .C(n_569), .Y(n_567) );
NAND2x1p5_ASAP7_75t_L g726 ( .A(n_419), .B(n_569), .Y(n_726) );
OR2x4_ASAP7_75t_L g1755 ( .A(n_419), .B(n_560), .Y(n_1755) );
INVx1_ASAP7_75t_L g1758 ( .A(n_419), .Y(n_1758) );
AND2x4_ASAP7_75t_L g1763 ( .A(n_419), .B(n_434), .Y(n_1763) );
OR2x6_ASAP7_75t_L g1779 ( .A(n_419), .B(n_576), .Y(n_1779) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND2xp33_ASAP7_75t_SL g555 ( .A(n_420), .B(n_422), .Y(n_555) );
BUFx3_ASAP7_75t_L g639 ( .A(n_420), .Y(n_639) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND3x4_ASAP7_75t_L g638 ( .A(n_422), .B(n_639), .C(n_640), .Y(n_638) );
AND2x2_ASAP7_75t_L g904 ( .A(n_422), .B(n_639), .Y(n_904) );
HB1xp67_ASAP7_75t_L g1748 ( .A(n_422), .Y(n_1748) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_424), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_654) );
AOI221x1_ASAP7_75t_L g978 ( .A1(n_424), .A2(n_951), .B1(n_958), .B2(n_979), .C(n_981), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_424), .A2(n_979), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_424), .A2(n_979), .B1(n_1122), .B2(n_1123), .Y(n_1121) );
HB1xp67_ASAP7_75t_L g1257 ( .A(n_424), .Y(n_1257) );
AOI22xp33_ASAP7_75t_L g1327 ( .A1(n_424), .A2(n_656), .B1(n_1328), .B2(n_1329), .Y(n_1327) );
AOI22xp5_ASAP7_75t_L g1346 ( .A1(n_424), .A2(n_656), .B1(n_1347), .B2(n_1348), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1394 ( .A1(n_424), .A2(n_979), .B1(n_1395), .B2(n_1396), .Y(n_1394) );
AOI22xp33_ASAP7_75t_L g1422 ( .A1(n_424), .A2(n_979), .B1(n_1423), .B2(n_1424), .Y(n_1422) );
AOI22xp33_ASAP7_75t_L g1489 ( .A1(n_424), .A2(n_979), .B1(n_1490), .B2(n_1491), .Y(n_1489) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g542 ( .A(n_430), .Y(n_542) );
AND4x1_ASAP7_75t_L g628 ( .A(n_431), .B(n_629), .C(n_637), .D(n_654), .Y(n_628) );
AND5x1_ASAP7_75t_L g947 ( .A(n_431), .B(n_948), .C(n_978), .D(n_992), .E(n_995), .Y(n_947) );
INVx2_ASAP7_75t_SL g1088 ( .A(n_431), .Y(n_1088) );
NAND4xp75_ASAP7_75t_L g1116 ( .A(n_431), .B(n_1117), .C(n_1120), .D(n_1137), .Y(n_1116) );
AND4x1_ASAP7_75t_L g1253 ( .A(n_431), .B(n_1254), .C(n_1258), .D(n_1260), .Y(n_1253) );
NAND3xp33_ASAP7_75t_SL g1384 ( .A(n_431), .B(n_1385), .C(n_1394), .Y(n_1384) );
INVx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g863 ( .A1(n_432), .A2(n_842), .B1(n_864), .B2(n_865), .C(n_866), .Y(n_863) );
INVx3_ASAP7_75t_L g1010 ( .A(n_432), .Y(n_1010) );
HB1xp67_ASAP7_75t_L g1219 ( .A(n_432), .Y(n_1219) );
BUFx2_ASAP7_75t_L g1169 ( .A(n_433), .Y(n_1169) );
BUFx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g580 ( .A(n_434), .Y(n_580) );
BUFx2_ASAP7_75t_L g643 ( .A(n_434), .Y(n_643) );
BUFx3_ASAP7_75t_L g724 ( .A(n_434), .Y(n_724) );
AND2x2_ASAP7_75t_L g739 ( .A(n_434), .B(n_737), .Y(n_739) );
BUFx2_ASAP7_75t_L g854 ( .A(n_434), .Y(n_854) );
BUFx2_ASAP7_75t_L g1026 ( .A(n_434), .Y(n_1026) );
BUFx2_ASAP7_75t_L g1431 ( .A(n_434), .Y(n_1431) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g1174 ( .A(n_437), .B(n_1175), .Y(n_1174) );
AOI221xp5_ASAP7_75t_L g1381 ( .A1(n_437), .A2(n_591), .B1(n_1382), .B2(n_1383), .C(n_1384), .Y(n_1381) );
INVx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx5_ASAP7_75t_L g997 ( .A(n_438), .Y(n_997) );
OR2x6_ASAP7_75t_L g438 ( .A(n_439), .B(n_445), .Y(n_438) );
OR2x2_ASAP7_75t_L g594 ( .A(n_439), .B(n_445), .Y(n_594) );
INVx2_ASAP7_75t_L g743 ( .A(n_439), .Y(n_743) );
INVx8_ASAP7_75t_L g468 ( .A(n_440), .Y(n_468) );
BUFx3_ASAP7_75t_L g642 ( .A(n_440), .Y(n_642) );
BUFx3_ASAP7_75t_L g652 ( .A(n_440), .Y(n_652) );
AND2x2_ASAP7_75t_L g736 ( .A(n_440), .B(n_737), .Y(n_736) );
HB1xp67_ASAP7_75t_L g991 ( .A(n_440), .Y(n_991) );
AND2x4_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
AND2x4_ASAP7_75t_L g549 ( .A(n_441), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVxp67_ASAP7_75t_L g550 ( .A(n_444), .Y(n_550) );
INVxp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g535 ( .A(n_446), .B(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g687 ( .A(n_446), .B(n_536), .Y(n_687) );
INVx1_ASAP7_75t_L g716 ( .A(n_446), .Y(n_716) );
INVx1_ASAP7_75t_L g1850 ( .A(n_446), .Y(n_1850) );
BUFx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g456 ( .A(n_447), .Y(n_456) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx8_ASAP7_75t_L g591 ( .A(n_450), .Y(n_591) );
AND2x4_ASAP7_75t_L g450 ( .A(n_451), .B(n_458), .Y(n_450) );
INVx1_ASAP7_75t_L g878 ( .A(n_451), .Y(n_878) );
OR2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_455), .Y(n_451) );
BUFx3_ASAP7_75t_L g781 ( .A(n_452), .Y(n_781) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_453), .Y(n_552) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g576 ( .A(n_454), .Y(n_576) );
INVx1_ASAP7_75t_L g469 ( .A(n_455), .Y(n_469) );
OR2x2_ASAP7_75t_L g539 ( .A(n_455), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g635 ( .A(n_455), .Y(n_635) );
OR2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
OR2x2_ASAP7_75t_L g554 ( .A(n_456), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_SL g680 ( .A(n_456), .B(n_499), .Y(n_680) );
INVx1_ASAP7_75t_L g809 ( .A(n_456), .Y(n_809) );
HB1xp67_ASAP7_75t_L g1750 ( .A(n_456), .Y(n_1750) );
INVx1_ASAP7_75t_L g737 ( .A(n_457), .Y(n_737) );
INVx1_ASAP7_75t_L g755 ( .A(n_457), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_458), .B(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g700 ( .A(n_459), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
AND2x6_ASAP7_75t_L g501 ( .A(n_460), .B(n_479), .Y(n_501) );
INVx1_ASAP7_75t_L g511 ( .A(n_460), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_460), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_460), .B(n_531), .Y(n_684) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_460), .B(n_841), .Y(n_1199) );
AND2x2_ASAP7_75t_L g523 ( .A(n_461), .B(n_477), .Y(n_523) );
INVx3_ASAP7_75t_L g610 ( .A(n_461), .Y(n_610) );
BUFx6f_ASAP7_75t_L g828 ( .A(n_461), .Y(n_828) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_462), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_466), .A2(n_582), .B1(n_1029), .B2(n_1030), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_466), .A2(n_582), .B1(n_1182), .B2(n_1183), .Y(n_1201) );
AOI22xp33_ASAP7_75t_L g1291 ( .A1(n_466), .A2(n_582), .B1(n_1277), .B2(n_1279), .Y(n_1291) );
AOI22xp33_ASAP7_75t_L g1413 ( .A1(n_466), .A2(n_582), .B1(n_1400), .B2(n_1402), .Y(n_1413) );
AND2x4_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
AND2x4_ASAP7_75t_L g876 ( .A(n_467), .B(n_469), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_467), .A2(n_860), .B1(n_892), .B2(n_915), .Y(n_914) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g578 ( .A(n_468), .Y(n_578) );
INVx8_ASAP7_75t_L g725 ( .A(n_468), .Y(n_725) );
CKINVDCx5p33_ASAP7_75t_R g784 ( .A(n_468), .Y(n_784) );
INVx3_ASAP7_75t_L g1023 ( .A(n_468), .Y(n_1023) );
AND2x4_ASAP7_75t_L g582 ( .A(n_469), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_532), .Y(n_470) );
OAI31xp33_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_502), .A3(n_520), .B(n_528), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g614 ( .A(n_474), .Y(n_614) );
INVx2_ASAP7_75t_L g1094 ( .A(n_474), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g1247 ( .A1(n_474), .A2(n_508), .B1(n_1209), .B2(n_1210), .Y(n_1247) );
INVx4_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx3_ASAP7_75t_L g952 ( .A(n_476), .Y(n_952) );
AND2x4_ASAP7_75t_SL g476 ( .A(n_477), .B(n_479), .Y(n_476) );
AND2x4_ASAP7_75t_L g505 ( .A(n_477), .B(n_506), .Y(n_505) );
AND2x4_ASAP7_75t_L g525 ( .A(n_477), .B(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g763 ( .A(n_477), .B(n_506), .Y(n_763) );
AND2x2_ASAP7_75t_L g825 ( .A(n_477), .B(n_705), .Y(n_825) );
BUFx2_ASAP7_75t_L g847 ( .A(n_477), .Y(n_847) );
HB1xp67_ASAP7_75t_L g1841 ( .A(n_478), .Y(n_1841) );
BUFx3_ASAP7_75t_L g497 ( .A(n_479), .Y(n_497) );
BUFx3_ASAP7_75t_L g517 ( .A(n_479), .Y(n_517) );
INVx1_ASAP7_75t_L g603 ( .A(n_479), .Y(n_603) );
BUFx3_ASAP7_75t_L g797 ( .A(n_479), .Y(n_797) );
BUFx6f_ASAP7_75t_L g1228 ( .A(n_479), .Y(n_1228) );
BUFx3_ASAP7_75t_L g1318 ( .A(n_479), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1827 ( .A(n_479), .B(n_1828), .Y(n_1827) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g1040 ( .A(n_480), .Y(n_1040) );
OAI221xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_484), .B1(n_485), .B2(n_491), .C(n_492), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g512 ( .A1(n_482), .A2(n_513), .B1(n_514), .B2(n_515), .C(n_516), .Y(n_512) );
INVx1_ASAP7_75t_L g670 ( .A(n_482), .Y(n_670) );
OAI221xp5_ASAP7_75t_L g1146 ( .A1(n_482), .A2(n_622), .B1(n_1147), .B2(n_1148), .C(n_1149), .Y(n_1146) );
OAI22xp5_ASAP7_75t_L g1286 ( .A1(n_482), .A2(n_621), .B1(n_1287), .B2(n_1288), .Y(n_1286) );
OAI221xp5_ASAP7_75t_L g1313 ( .A1(n_482), .A2(n_1314), .B1(n_1315), .B2(n_1316), .C(n_1317), .Y(n_1313) );
OAI221xp5_ASAP7_75t_L g1445 ( .A1(n_482), .A2(n_1315), .B1(n_1446), .B2(n_1447), .C(n_1448), .Y(n_1445) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_SL g619 ( .A(n_483), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_483), .A2(n_800), .B1(n_801), .B2(n_802), .Y(n_799) );
OAI22x1_ASAP7_75t_SL g805 ( .A1(n_483), .A2(n_782), .B1(n_802), .B2(n_806), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_484), .A2(n_546), .B1(n_547), .B2(n_551), .Y(n_545) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
HB1xp67_ASAP7_75t_L g1315 ( .A(n_486), .Y(n_1315) );
INVx2_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g623 ( .A(n_487), .Y(n_623) );
INVx2_ASAP7_75t_L g802 ( .A(n_487), .Y(n_802) );
INVx4_ASAP7_75t_L g962 ( .A(n_487), .Y(n_962) );
BUFx6f_ASAP7_75t_L g1062 ( .A(n_487), .Y(n_1062) );
INVx1_ASAP7_75t_L g1481 ( .A(n_487), .Y(n_1481) );
INVx1_ASAP7_75t_L g1806 ( .A(n_487), .Y(n_1806) );
INVx8_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g514 ( .A(n_488), .Y(n_514) );
OR2x2_ASAP7_75t_L g1844 ( .A(n_488), .B(n_1832), .Y(n_1844) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OAI221xp5_ASAP7_75t_L g570 ( .A1(n_491), .A2(n_571), .B1(n_574), .B2(n_575), .C(n_577), .Y(n_570) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g606 ( .A(n_494), .Y(n_606) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_495), .Y(n_506) );
BUFx3_ASAP7_75t_L g798 ( .A(n_495), .Y(n_798) );
AND2x4_ASAP7_75t_L g1847 ( .A(n_495), .B(n_1841), .Y(n_1847) );
HB1xp67_ASAP7_75t_SL g1508 ( .A(n_498), .Y(n_1508) );
INVx4_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_SL g607 ( .A(n_499), .Y(n_607) );
AND2x4_ASAP7_75t_L g807 ( .A(n_499), .B(n_808), .Y(n_807) );
INVx4_ASAP7_75t_L g833 ( .A(n_499), .Y(n_833) );
NAND4xp25_ASAP7_75t_L g963 ( .A(n_499), .B(n_964), .C(n_965), .D(n_967), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g1801 ( .A(n_499), .B(n_808), .Y(n_1801) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_501), .A2(n_601), .B(n_608), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g1036 ( .A1(n_501), .A2(n_1037), .B(n_1043), .Y(n_1036) );
AOI21xp5_ASAP7_75t_L g1104 ( .A1(n_501), .A2(n_1105), .B(n_1107), .Y(n_1104) );
AOI21xp5_ASAP7_75t_SL g1139 ( .A1(n_501), .A2(n_1140), .B(n_1143), .Y(n_1139) );
AOI221xp5_ASAP7_75t_SL g1184 ( .A1(n_501), .A2(n_525), .B1(n_1175), .B2(n_1185), .C(n_1187), .Y(n_1184) );
AOI21xp5_ASAP7_75t_L g1225 ( .A1(n_501), .A2(n_1226), .B(n_1232), .Y(n_1225) );
AOI21xp5_ASAP7_75t_L g1269 ( .A1(n_501), .A2(n_1270), .B(n_1271), .Y(n_1269) );
AOI21xp5_ASAP7_75t_L g1302 ( .A1(n_501), .A2(n_504), .B(n_1303), .Y(n_1302) );
AOI21xp5_ASAP7_75t_L g1365 ( .A1(n_501), .A2(n_1366), .B(n_1367), .Y(n_1365) );
AOI221xp5_ASAP7_75t_L g1403 ( .A1(n_501), .A2(n_525), .B1(n_1382), .B2(n_1404), .C(n_1406), .Y(n_1403) );
AOI21xp5_ASAP7_75t_L g1438 ( .A1(n_501), .A2(n_1439), .B(n_1440), .Y(n_1438) );
AOI21xp5_ASAP7_75t_L g1470 ( .A1(n_501), .A2(n_1471), .B(n_1474), .Y(n_1470) );
AOI21xp5_ASAP7_75t_SL g1505 ( .A1(n_501), .A2(n_1506), .B(n_1509), .Y(n_1505) );
INVxp67_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_504), .A2(n_522), .B1(n_598), .B2(n_599), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_504), .A2(n_1034), .B1(n_1112), .B2(n_1113), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1368 ( .A1(n_504), .A2(n_522), .B1(n_1369), .B2(n_1370), .Y(n_1368) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_504), .A2(n_1400), .B1(n_1401), .B2(n_1402), .Y(n_1399) );
AOI22xp5_ASAP7_75t_L g1441 ( .A1(n_504), .A2(n_1034), .B1(n_1442), .B2(n_1443), .Y(n_1441) );
AOI22xp33_ASAP7_75t_L g1510 ( .A1(n_504), .A2(n_1034), .B1(n_1511), .B2(n_1512), .Y(n_1510) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_505), .A2(n_1029), .B1(n_1030), .B2(n_1034), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1144 ( .A1(n_505), .A2(n_522), .B1(n_1125), .B2(n_1126), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_505), .A2(n_522), .B1(n_1182), .B2(n_1183), .Y(n_1181) );
INVx1_ASAP7_75t_L g1239 ( .A(n_505), .Y(n_1239) );
HB1xp67_ASAP7_75t_L g1278 ( .A(n_505), .Y(n_1278) );
BUFx6f_ASAP7_75t_L g1042 ( .A(n_506), .Y(n_1042) );
INVx2_ASAP7_75t_L g1101 ( .A(n_506), .Y(n_1101) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g616 ( .A(n_508), .Y(n_616) );
NOR2x1_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g686 ( .A(n_510), .Y(n_686) );
BUFx2_ASAP7_75t_L g841 ( .A(n_510), .Y(n_841) );
AND2x4_ASAP7_75t_L g1831 ( .A(n_510), .B(n_1832), .Y(n_1831) );
INVx1_ASAP7_75t_L g846 ( .A(n_511), .Y(n_846) );
OAI22xp33_ASAP7_75t_L g556 ( .A1(n_513), .A2(n_557), .B1(n_561), .B2(n_562), .Y(n_556) );
INVx1_ASAP7_75t_L g691 ( .A(n_514), .Y(n_691) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g627 ( .A(n_519), .Y(n_627) );
OAI221xp5_ASAP7_75t_L g1050 ( .A1(n_519), .A2(n_676), .B1(n_1051), .B2(n_1052), .C(n_1055), .Y(n_1050) );
INVx2_ASAP7_75t_L g1244 ( .A(n_519), .Y(n_1244) );
INVx1_ASAP7_75t_L g1410 ( .A(n_519), .Y(n_1410) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_522), .A2(n_525), .B1(n_1305), .B2(n_1306), .Y(n_1304) );
HB1xp67_ASAP7_75t_L g1401 ( .A(n_522), .Y(n_1401) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x4_ASAP7_75t_L g715 ( .A(n_523), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g1035 ( .A(n_523), .Y(n_1035) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_R g1048 ( .A(n_525), .B(n_1009), .Y(n_1048) );
INVx2_ASAP7_75t_SL g1103 ( .A(n_525), .Y(n_1103) );
BUFx2_ASAP7_75t_L g1189 ( .A(n_526), .Y(n_1189) );
INVx1_ASAP7_75t_L g1275 ( .A(n_526), .Y(n_1275) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g612 ( .A(n_527), .Y(n_612) );
BUFx3_ASAP7_75t_L g829 ( .A(n_527), .Y(n_829) );
BUFx3_ASAP7_75t_L g1047 ( .A(n_527), .Y(n_1047) );
OAI21xp5_ASAP7_75t_L g595 ( .A1(n_528), .A2(n_596), .B(n_613), .Y(n_595) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_529), .B(n_757), .Y(n_943) );
BUFx2_ASAP7_75t_L g1064 ( .A(n_529), .Y(n_1064) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g695 ( .A(n_530), .B(n_696), .Y(n_695) );
OR2x6_ASAP7_75t_L g862 ( .A(n_530), .B(n_726), .Y(n_862) );
BUFx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g640 ( .A(n_531), .Y(n_640) );
AOI21xp5_ASAP7_75t_SL g532 ( .A1(n_533), .A2(n_543), .B(n_544), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g1360 ( .A1(n_533), .A2(n_1361), .B(n_1362), .Y(n_1360) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
HB1xp67_ASAP7_75t_L g1290 ( .A(n_534), .Y(n_1290) );
AND2x4_ASAP7_75t_L g534 ( .A(n_535), .B(n_539), .Y(n_534) );
INVx2_ASAP7_75t_SL g813 ( .A(n_535), .Y(n_813) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g875 ( .A(n_539), .Y(n_875) );
INVx3_ASAP7_75t_L g563 ( .A(n_540), .Y(n_563) );
BUFx6f_ASAP7_75t_L g1816 ( .A(n_540), .Y(n_1816) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
BUFx2_ASAP7_75t_L g750 ( .A(n_541), .Y(n_750) );
BUFx3_ASAP7_75t_L g1892 ( .A(n_541), .Y(n_1892) );
BUFx2_ASAP7_75t_L g1772 ( .A(n_542), .Y(n_1772) );
INVx1_ASAP7_75t_L g1428 ( .A(n_547), .Y(n_1428) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g646 ( .A(n_548), .Y(n_646) );
BUFx6f_ASAP7_75t_L g856 ( .A(n_548), .Y(n_856) );
BUFx6f_ASAP7_75t_L g858 ( .A(n_548), .Y(n_858) );
AND2x4_ASAP7_75t_L g1757 ( .A(n_548), .B(n_1758), .Y(n_1757) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_549), .Y(n_573) );
BUFx8_ASAP7_75t_L g583 ( .A(n_549), .Y(n_583) );
INVx2_ASAP7_75t_L g721 ( .A(n_549), .Y(n_721) );
OAI221xp5_ASAP7_75t_L g982 ( .A1(n_551), .A2(n_906), .B1(n_983), .B2(n_984), .C(n_985), .Y(n_982) );
OAI22xp5_ASAP7_75t_L g1893 ( .A1(n_551), .A2(n_557), .B1(n_1874), .B2(n_1882), .Y(n_1893) );
INVx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx3_ASAP7_75t_L g899 ( .A(n_552), .Y(n_899) );
INVx3_ASAP7_75t_L g908 ( .A(n_552), .Y(n_908) );
OAI22xp5_ASAP7_75t_SL g981 ( .A1(n_553), .A2(n_982), .B1(n_986), .B2(n_988), .Y(n_981) );
BUFx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx4f_ASAP7_75t_L g1810 ( .A(n_554), .Y(n_1810) );
BUFx2_ASAP7_75t_L g731 ( .A(n_555), .Y(n_731) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_559), .A2(n_898), .B1(n_899), .B2(n_900), .Y(n_897) );
HB1xp67_ASAP7_75t_L g1885 ( .A(n_559), .Y(n_1885) );
BUFx4f_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g633 ( .A(n_560), .Y(n_633) );
OR2x4_ASAP7_75t_L g1776 ( .A(n_560), .B(n_1758), .Y(n_1776) );
BUFx3_ASAP7_75t_L g1814 ( .A(n_560), .Y(n_1814) );
OAI22xp5_ASAP7_75t_L g1821 ( .A1(n_562), .A2(n_632), .B1(n_1790), .B2(n_1798), .Y(n_1821) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx3_ASAP7_75t_L g791 ( .A(n_563), .Y(n_791) );
OAI33xp33_ASAP7_75t_L g1883 ( .A1(n_564), .A2(n_1809), .A3(n_1884), .B1(n_1888), .B2(n_1889), .B3(n_1893), .Y(n_1883) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AOI33xp33_ASAP7_75t_L g637 ( .A1(n_565), .A2(n_638), .A3(n_641), .B1(n_644), .B2(n_649), .B3(n_650), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g1170 ( .A(n_565), .B(n_1171), .C(n_1172), .Y(n_1170) );
BUFx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
BUFx2_ASAP7_75t_L g1021 ( .A(n_566), .Y(n_1021) );
BUFx2_ASAP7_75t_L g1084 ( .A(n_566), .Y(n_1084) );
BUFx2_ASAP7_75t_L g1216 ( .A(n_566), .Y(n_1216) );
INVx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx3_ASAP7_75t_L g987 ( .A(n_567), .Y(n_987) );
INVx1_ASAP7_75t_L g1263 ( .A(n_571), .Y(n_1263) );
BUFx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OAI221xp5_ASAP7_75t_L g988 ( .A1(n_572), .A2(n_781), .B1(n_969), .B2(n_989), .C(n_990), .Y(n_988) );
INVx8_ASAP7_75t_L g1215 ( .A(n_572), .Y(n_1215) );
INVx5_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx3_ASAP7_75t_L g730 ( .A(n_573), .Y(n_730) );
INVx2_ASAP7_75t_SL g906 ( .A(n_573), .Y(n_906) );
HB1xp67_ASAP7_75t_L g1333 ( .A(n_573), .Y(n_1333) );
INVx2_ASAP7_75t_SL g1337 ( .A(n_573), .Y(n_1337) );
OAI22xp5_ASAP7_75t_L g1818 ( .A1(n_575), .A2(n_1794), .B1(n_1807), .B2(n_1819), .Y(n_1818) );
BUFx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g653 ( .A(n_580), .Y(n_653) );
INVx2_ASAP7_75t_L g728 ( .A(n_580), .Y(n_728) );
INVx2_ASAP7_75t_L g860 ( .A(n_580), .Y(n_860) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g636 ( .A(n_582), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_582), .A2(n_876), .B1(n_1125), .B2(n_1126), .Y(n_1124) );
HB1xp67_ASAP7_75t_L g1130 ( .A(n_583), .Y(n_1130) );
INVx3_ASAP7_75t_L g1357 ( .A(n_583), .Y(n_1357) );
INVx2_ASAP7_75t_SL g1389 ( .A(n_583), .Y(n_1389) );
INVx3_ASAP7_75t_L g1496 ( .A(n_583), .Y(n_1496) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AO21x2_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B(n_658), .Y(n_587) );
NAND3xp33_ASAP7_75t_SL g589 ( .A(n_590), .B(n_595), .C(n_628), .Y(n_589) );
AOI21xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B(n_593), .Y(n_590) );
AOI211x1_ASAP7_75t_L g1000 ( .A1(n_591), .A2(n_1001), .B(n_1002), .C(n_1027), .Y(n_1000) );
AOI21xp33_ASAP7_75t_SL g1089 ( .A1(n_591), .A2(n_1090), .B(n_1091), .Y(n_1089) );
AOI21xp5_ASAP7_75t_L g1117 ( .A1(n_591), .A2(n_1118), .B(n_1119), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_591), .B(n_1203), .Y(n_1202) );
AOI21xp5_ASAP7_75t_L g1220 ( .A1(n_591), .A2(n_1221), .B(n_1222), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_591), .B(n_1293), .Y(n_1292) );
AOI21xp33_ASAP7_75t_SL g1322 ( .A1(n_591), .A2(n_1323), .B(n_1324), .Y(n_1322) );
AOI211x1_ASAP7_75t_L g1343 ( .A1(n_591), .A2(n_1344), .B(n_1345), .C(n_1359), .Y(n_1343) );
AOI21xp33_ASAP7_75t_SL g1433 ( .A1(n_591), .A2(n_1434), .B(n_1435), .Y(n_1433) );
AOI21xp5_ASAP7_75t_L g1465 ( .A1(n_591), .A2(n_1466), .B(n_1467), .Y(n_1465) );
AOI21xp33_ASAP7_75t_SL g1500 ( .A1(n_591), .A2(n_1501), .B(n_1502), .Y(n_1500) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_594), .B(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g626 ( .A(n_603), .Y(n_626) );
INVx1_ASAP7_75t_L g1150 ( .A(n_603), .Y(n_1150) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g1142 ( .A(n_606), .Y(n_1142) );
HB1xp67_ASAP7_75t_L g1243 ( .A(n_606), .Y(n_1243) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g966 ( .A(n_610), .Y(n_966) );
INVx2_ASAP7_75t_L g1044 ( .A(n_610), .Y(n_1044) );
INVx1_ASAP7_75t_L g1106 ( .A(n_610), .Y(n_1106) );
INVx2_ASAP7_75t_SL g1188 ( .A(n_610), .Y(n_1188) );
INVx2_ASAP7_75t_L g1233 ( .A(n_610), .Y(n_1233) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx3_ASAP7_75t_L g705 ( .A(n_612), .Y(n_705) );
BUFx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OAI221xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_620), .B1(n_621), .B2(n_624), .C(n_625), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g1872 ( .A1(n_618), .A2(n_1873), .B1(n_1874), .B2(n_1875), .Y(n_1872) );
OAI22xp33_ASAP7_75t_L g1877 ( .A1(n_618), .A2(n_1795), .B1(n_1878), .B2(n_1879), .Y(n_1877) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
BUFx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g669 ( .A(n_622), .Y(n_669) );
OAI221xp5_ASAP7_75t_L g1514 ( .A1(n_622), .A2(n_1058), .B1(n_1515), .B2(n_1516), .C(n_1517), .Y(n_1514) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g1285 ( .A(n_627), .Y(n_1285) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_631), .B(n_714), .Y(n_994) );
OR2x6_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
OR2x2_ASAP7_75t_L g1087 ( .A(n_632), .B(n_634), .Y(n_1087) );
INVx2_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
INVxp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g870 ( .A(n_635), .B(n_871), .Y(n_870) );
AOI33xp33_ASAP7_75t_L g852 ( .A1(n_638), .A2(n_853), .A3(n_855), .B1(n_857), .B2(n_859), .B3(n_861), .Y(n_852) );
BUFx3_ASAP7_75t_L g1012 ( .A(n_638), .Y(n_1012) );
AOI33xp33_ASAP7_75t_L g1076 ( .A1(n_638), .A2(n_1077), .A3(n_1080), .B1(n_1083), .B2(n_1084), .B3(n_1085), .Y(n_1076) );
AOI33xp33_ASAP7_75t_L g1330 ( .A1(n_638), .A2(n_1216), .A3(n_1331), .B1(n_1332), .B2(n_1335), .B3(n_1338), .Y(n_1330) );
AOI33xp33_ASAP7_75t_L g1425 ( .A1(n_638), .A2(n_1216), .A3(n_1426), .B1(n_1427), .B2(n_1429), .B3(n_1430), .Y(n_1425) );
AOI33xp33_ASAP7_75t_L g1492 ( .A1(n_638), .A2(n_1216), .A3(n_1493), .B1(n_1494), .B2(n_1497), .B3(n_1498), .Y(n_1492) );
INVx3_ASAP7_75t_L g1767 ( .A(n_639), .Y(n_1767) );
INVx1_ASAP7_75t_L g759 ( .A(n_640), .Y(n_759) );
OAI31xp33_ASAP7_75t_SL g772 ( .A1(n_640), .A2(n_773), .A3(n_774), .B(n_778), .Y(n_772) );
OAI31xp33_ASAP7_75t_L g894 ( .A1(n_640), .A2(n_895), .A3(n_896), .B(n_913), .Y(n_894) );
INVx2_ASAP7_75t_SL g1114 ( .A(n_640), .Y(n_1114) );
INVx2_ASAP7_75t_SL g1015 ( .A(n_642), .Y(n_1015) );
INVx1_ASAP7_75t_L g1079 ( .A(n_642), .Y(n_1079) );
BUFx3_ASAP7_75t_L g1136 ( .A(n_642), .Y(n_1136) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g1888 ( .A1(n_646), .A2(n_908), .B1(n_1868), .B2(n_1878), .Y(n_1888) );
BUFx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
BUFx2_ASAP7_75t_L g722 ( .A(n_648), .Y(n_722) );
BUFx12f_ASAP7_75t_L g733 ( .A(n_648), .Y(n_733) );
AND2x4_ASAP7_75t_L g757 ( .A(n_648), .B(n_755), .Y(n_757) );
INVx5_ASAP7_75t_L g1018 ( .A(n_648), .Y(n_1018) );
BUFx3_ASAP7_75t_L g1131 ( .A(n_648), .Y(n_1131) );
BUFx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AO22x2_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_1068), .B1(n_1152), .B2(n_1153), .Y(n_659) );
XOR2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_817), .Y(n_660) );
XNOR2x1_ASAP7_75t_L g1153 ( .A(n_661), .B(n_817), .Y(n_1153) );
BUFx2_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
INVxp67_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
XNOR2x1_ASAP7_75t_L g663 ( .A(n_664), .B(n_765), .Y(n_663) );
XNOR2x1_ASAP7_75t_L g664 ( .A(n_665), .B(n_764), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_717), .Y(n_665) );
NAND3xp33_ASAP7_75t_SL g666 ( .A(n_667), .B(n_697), .C(n_711), .Y(n_666) );
AOI211xp5_ASAP7_75t_SL g667 ( .A1(n_668), .A2(n_671), .B(n_681), .C(n_690), .Y(n_667) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g692 ( .A1(n_673), .A2(n_676), .B1(n_693), .B2(n_694), .C(n_695), .Y(n_692) );
BUFx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g933 ( .A(n_674), .Y(n_933) );
BUFx2_ASAP7_75t_L g961 ( .A(n_674), .Y(n_961) );
BUFx2_ASAP7_75t_L g1054 ( .A(n_674), .Y(n_1054) );
INVxp67_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
BUFx4f_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OR2x6_ASAP7_75t_L g688 ( .A(n_677), .B(n_689), .Y(n_688) );
INVx4_ASAP7_75t_L g839 ( .A(n_677), .Y(n_839) );
BUFx4f_ASAP7_75t_L g849 ( .A(n_677), .Y(n_849) );
BUFx4f_ASAP7_75t_L g1310 ( .A(n_677), .Y(n_1310) );
BUFx6f_ASAP7_75t_L g1795 ( .A(n_677), .Y(n_1795) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
BUFx3_ASAP7_75t_L g709 ( .A(n_678), .Y(n_709) );
OAI21xp5_ASAP7_75t_L g930 ( .A1(n_679), .A2(n_688), .B(n_931), .Y(n_930) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g812 ( .A(n_682), .Y(n_812) );
INVx2_ASAP7_75t_SL g927 ( .A(n_682), .Y(n_927) );
NAND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_685), .Y(n_682) );
INVx1_ASAP7_75t_L g689 ( .A(n_683), .Y(n_689) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_SL g925 ( .A(n_687), .Y(n_925) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_688), .Y(n_816) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_695), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_695), .B(n_922), .Y(n_921) );
INVx2_ASAP7_75t_L g1783 ( .A(n_695), .Y(n_1783) );
INVx2_ASAP7_75t_L g1871 ( .A(n_695), .Y(n_1871) );
AOI222xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_701), .B1(n_702), .B2(n_706), .C1(n_707), .C2(n_710), .Y(n_697) );
AOI21xp33_ASAP7_75t_SL g814 ( .A1(n_698), .A2(n_815), .B(n_816), .Y(n_814) );
AND2x4_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
AOI222xp33_ASAP7_75t_L g810 ( .A1(n_702), .A2(n_776), .B1(n_788), .B2(n_811), .C1(n_812), .C2(n_813), .Y(n_810) );
INVx1_ASAP7_75t_L g939 ( .A(n_702), .Y(n_939) );
AND2x4_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g708 ( .A(n_704), .B(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g929 ( .A(n_704), .B(n_709), .Y(n_929) );
AOI211xp5_ASAP7_75t_L g740 ( .A1(n_706), .A2(n_741), .B(n_744), .C(n_752), .Y(n_740) );
AOI222xp33_ASAP7_75t_L g795 ( .A1(n_707), .A2(n_777), .B1(n_796), .B2(n_803), .C1(n_804), .C2(n_807), .Y(n_795) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_SL g971 ( .A(n_709), .Y(n_971) );
BUFx2_ASAP7_75t_SL g1282 ( .A(n_709), .Y(n_1282) );
BUFx3_ASAP7_75t_L g1825 ( .A(n_709), .Y(n_1825) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx3_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_715), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_715), .A2(n_762), .B1(n_892), .B2(n_893), .Y(n_891) );
AND2x4_ASAP7_75t_L g762 ( .A(n_716), .B(n_763), .Y(n_762) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_740), .B(n_758), .C(n_760), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_723), .B1(n_727), .B2(n_732), .C(n_734), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
OR2x6_ASAP7_75t_SL g753 ( .A(n_721), .B(n_754), .Y(n_753) );
INVx3_ASAP7_75t_L g871 ( .A(n_721), .Y(n_871) );
BUFx2_ASAP7_75t_L g1082 ( .A(n_721), .Y(n_1082) );
BUFx2_ASAP7_75t_L g1134 ( .A(n_721), .Y(n_1134) );
BUFx2_ASAP7_75t_L g1266 ( .A(n_725), .Y(n_1266) );
INVx3_ASAP7_75t_L g786 ( .A(n_726), .Y(n_786) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI221xp5_ASAP7_75t_L g779 ( .A1(n_730), .A2(n_780), .B1(n_781), .B2(n_782), .C(n_783), .Y(n_779) );
OAI221xp5_ASAP7_75t_L g901 ( .A1(n_730), .A2(n_750), .B1(n_902), .B2(n_903), .C(n_904), .Y(n_901) );
BUFx2_ASAP7_75t_L g1020 ( .A(n_733), .Y(n_1020) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_736), .A2(n_739), .B1(n_768), .B2(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx4_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_746), .A2(n_748), .B1(n_776), .B2(n_777), .Y(n_775) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI221xp5_ASAP7_75t_L g896 ( .A1(n_749), .A2(n_897), .B1(n_901), .B2(n_905), .C(n_910), .Y(n_896) );
OR2x6_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g1761 ( .A(n_750), .Y(n_1761) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
HB1xp67_ASAP7_75t_L g917 ( .A(n_755), .Y(n_917) );
INVx3_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
HB1xp67_ASAP7_75t_L g974 ( .A(n_758), .Y(n_974) );
INVx1_ASAP7_75t_L g1249 ( .A(n_758), .Y(n_1249) );
INVx1_ASAP7_75t_L g1321 ( .A(n_758), .Y(n_1321) );
BUFx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AOI21x1_ASAP7_75t_L g822 ( .A1(n_759), .A2(n_823), .B(n_850), .Y(n_822) );
HB1xp67_ASAP7_75t_L g1151 ( .A(n_759), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_762), .B(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g872 ( .A(n_762), .Y(n_872) );
AOI211x1_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_768), .B(n_769), .C(n_794), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
NAND3xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_787), .C(n_789), .Y(n_778) );
INVx3_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
OAI211xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_791), .B(n_792), .C(n_793), .Y(n_789) );
OAI21xp5_ASAP7_75t_SL g910 ( .A1(n_791), .A2(n_911), .B(n_912), .Y(n_910) );
NAND3xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_810), .C(n_814), .Y(n_794) );
BUFx2_ASAP7_75t_L g1405 ( .A(n_798), .Y(n_1405) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
AO22x2_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_998), .B1(n_1066), .B2(n_1067), .Y(n_817) );
INVx1_ASAP7_75t_L g1066 ( .A(n_818), .Y(n_1066) );
XNOR2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_946), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_887), .B1(n_944), .B2(n_945), .Y(n_819) );
INVx1_ASAP7_75t_L g945 ( .A(n_820), .Y(n_945) );
NAND3xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_880), .C(n_884), .Y(n_820) );
INVx1_ASAP7_75t_L g881 ( .A(n_822), .Y(n_881) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_830), .B1(n_831), .B2(n_832), .Y(n_826) );
INVx3_ASAP7_75t_L g1194 ( .A(n_828), .Y(n_1194) );
BUFx6f_ASAP7_75t_L g1273 ( .A(n_828), .Y(n_1273) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_846), .B1(n_847), .B2(n_848), .Y(n_834) );
INVx3_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx4_ASAP7_75t_L g955 ( .A(n_837), .Y(n_955) );
BUFx6f_ASAP7_75t_L g1059 ( .A(n_837), .Y(n_1059) );
INVx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g956 ( .A(n_839), .Y(n_956) );
AOI22xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_842), .B1(n_843), .B2(n_845), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_841), .A2(n_843), .B1(n_958), .B2(n_959), .Y(n_957) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
AOI222xp33_ASAP7_75t_L g874 ( .A1(n_845), .A2(n_875), .B1(n_876), .B2(n_877), .C1(n_878), .C2(n_879), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g953 ( .A1(n_846), .A2(n_847), .B1(n_954), .B2(n_960), .Y(n_953) );
INVx1_ASAP7_75t_L g882 ( .A(n_851), .Y(n_882) );
AND2x2_ASAP7_75t_L g851 ( .A(n_852), .B(n_863), .Y(n_851) );
INVx1_ASAP7_75t_L g1890 ( .A(n_858), .Y(n_1890) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g886 ( .A(n_867), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_873), .Y(n_867) );
NAND2x1_ASAP7_75t_L g868 ( .A(n_869), .B(n_872), .Y(n_868) );
INVx2_ASAP7_75t_SL g869 ( .A(n_870), .Y(n_869) );
INVx2_ASAP7_75t_L g1819 ( .A(n_871), .Y(n_1819) );
INVx1_ASAP7_75t_L g885 ( .A(n_874), .Y(n_885) );
AOI22xp5_ASAP7_75t_L g976 ( .A1(n_875), .A2(n_878), .B1(n_959), .B2(n_977), .Y(n_976) );
OAI21xp5_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_882), .B(n_883), .Y(n_880) );
OAI21xp33_ASAP7_75t_L g884 ( .A1(n_883), .A2(n_885), .B(n_886), .Y(n_884) );
INVx1_ASAP7_75t_L g944 ( .A(n_887), .Y(n_944) );
XNOR2xp5_ASAP7_75t_L g887 ( .A(n_888), .B(n_889), .Y(n_887) );
NOR2x1_ASAP7_75t_L g889 ( .A(n_890), .B(n_918), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_891), .B(n_894), .Y(n_890) );
OAI22xp5_ASAP7_75t_L g1817 ( .A1(n_899), .A2(n_1337), .B1(n_1792), .B2(n_1804), .Y(n_1817) );
OAI211xp5_ASAP7_75t_L g931 ( .A1(n_902), .A2(n_932), .B(n_934), .C(n_935), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_906), .A2(n_907), .B1(n_908), .B2(n_909), .Y(n_905) );
AOI22xp5_ASAP7_75t_L g924 ( .A1(n_915), .A2(n_925), .B1(n_926), .B2(n_927), .Y(n_924) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
NAND3xp33_ASAP7_75t_L g918 ( .A(n_919), .B(n_936), .C(n_940), .Y(n_918) );
NOR3xp33_ASAP7_75t_SL g919 ( .A(n_920), .B(n_928), .C(n_930), .Y(n_919) );
OAI21xp5_ASAP7_75t_SL g920 ( .A1(n_921), .A2(n_923), .B(n_924), .Y(n_920) );
INVx2_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_937), .B(n_938), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_941), .B(n_942), .Y(n_940) );
AOI21xp5_ASAP7_75t_L g948 ( .A1(n_949), .A2(n_974), .B(n_975), .Y(n_948) );
NAND4xp25_ASAP7_75t_L g949 ( .A(n_950), .B(n_953), .C(n_963), .D(n_968), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_951), .B(n_952), .Y(n_950) );
INVx1_ASAP7_75t_L g1197 ( .A(n_952), .Y(n_1197) );
AOI222xp33_ASAP7_75t_L g1407 ( .A1(n_952), .A2(n_1395), .B1(n_1396), .B2(n_1408), .C1(n_1409), .C2(n_1411), .Y(n_1407) );
OAI22xp5_ASAP7_75t_L g1867 ( .A1(n_961), .A2(n_1868), .B1(n_1869), .B2(n_1870), .Y(n_1867) );
OAI22xp5_ASAP7_75t_L g1880 ( .A1(n_961), .A2(n_1875), .B1(n_1881), .B2(n_1882), .Y(n_1880) );
INVx2_ASAP7_75t_L g1876 ( .A(n_962), .Y(n_1876) );
OAI211xp5_ASAP7_75t_L g968 ( .A1(n_969), .A2(n_970), .B(n_972), .C(n_973), .Y(n_968) );
OAI211xp5_ASAP7_75t_L g1372 ( .A1(n_970), .A2(n_1373), .B(n_1374), .C(n_1375), .Y(n_1372) );
OAI22xp5_ASAP7_75t_L g1796 ( .A1(n_970), .A2(n_1793), .B1(n_1797), .B2(n_1798), .Y(n_1796) );
INVx5_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_979), .A2(n_1255), .B1(n_1256), .B2(n_1257), .Y(n_1254) );
INVx2_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
INVx2_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
AOI33xp33_ASAP7_75t_L g1351 ( .A1(n_987), .A2(n_1012), .A3(n_1352), .B1(n_1353), .B2(n_1355), .B3(n_1358), .Y(n_1351) );
CKINVDCx5p33_ASAP7_75t_R g1392 ( .A(n_987), .Y(n_1392) );
INVx2_ASAP7_75t_L g1820 ( .A(n_987), .Y(n_1820) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_996), .B(n_997), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_997), .B(n_1009), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_997), .B(n_1259), .Y(n_1258) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_997), .B(n_1350), .Y(n_1349) );
INVx2_ASAP7_75t_L g1067 ( .A(n_998), .Y(n_1067) );
XOR2x2_ASAP7_75t_L g998 ( .A(n_999), .B(n_1065), .Y(n_998) );
NAND2xp5_ASAP7_75t_SL g999 ( .A(n_1000), .B(n_1031), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1011), .Y(n_1002) );
NOR2xp33_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1007), .Y(n_1003) );
NAND2xp5_ASAP7_75t_SL g1007 ( .A(n_1008), .B(n_1010), .Y(n_1007) );
NAND3xp33_ASAP7_75t_L g1173 ( .A(n_1010), .B(n_1174), .C(n_1176), .Y(n_1173) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1010), .Y(n_1340) );
NAND4xp25_ASAP7_75t_SL g1345 ( .A(n_1010), .B(n_1346), .C(n_1349), .D(n_1351), .Y(n_1345) );
AOI33xp33_ASAP7_75t_L g1011 ( .A1(n_1012), .A2(n_1013), .A3(n_1016), .B1(n_1019), .B2(n_1021), .B3(n_1022), .Y(n_1011) );
AOI33xp33_ASAP7_75t_L g1127 ( .A1(n_1012), .A2(n_1084), .A3(n_1128), .B1(n_1129), .B2(n_1132), .B3(n_1135), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1012), .B(n_1168), .Y(n_1167) );
AOI33xp33_ASAP7_75t_L g1211 ( .A1(n_1012), .A2(n_1212), .A3(n_1213), .B1(n_1214), .B2(n_1216), .B3(n_1217), .Y(n_1211) );
AOI33xp33_ASAP7_75t_L g1260 ( .A1(n_1012), .A2(n_1084), .A3(n_1261), .B1(n_1262), .B2(n_1264), .B3(n_1265), .Y(n_1260) );
AOI33xp33_ASAP7_75t_L g1385 ( .A1(n_1012), .A2(n_1386), .A3(n_1387), .B1(n_1390), .B2(n_1391), .B3(n_1393), .Y(n_1385) );
AOI33xp33_ASAP7_75t_L g1459 ( .A1(n_1012), .A2(n_1391), .A3(n_1460), .B1(n_1461), .B2(n_1462), .B3(n_1463), .Y(n_1459) );
INVx2_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx2_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx2_ASAP7_75t_R g1334 ( .A(n_1018), .Y(n_1334) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1018), .Y(n_1354) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
OAI21xp5_ASAP7_75t_L g1031 ( .A1(n_1032), .A2(n_1049), .B(n_1063), .Y(n_1031) );
NAND3xp33_ASAP7_75t_SL g1032 ( .A(n_1033), .B(n_1036), .C(n_1048), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_1034), .A2(n_1236), .B1(n_1237), .B2(n_1238), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1276 ( .A1(n_1034), .A2(n_1277), .B1(n_1278), .B2(n_1279), .Y(n_1276) );
INVx2_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
INVx2_ASAP7_75t_L g1186 ( .A(n_1039), .Y(n_1186) );
BUFx2_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1040), .Y(n_1110) );
BUFx3_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
INVx1_ASAP7_75t_SL g1045 ( .A(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_SL g1046 ( .A(n_1047), .Y(n_1046) );
BUFx3_ASAP7_75t_L g1234 ( .A(n_1047), .Y(n_1234) );
OAI221xp5_ASAP7_75t_L g1281 ( .A1(n_1052), .A2(n_1282), .B1(n_1283), .B2(n_1284), .C(n_1285), .Y(n_1281) );
INVx2_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx2_ASAP7_75t_L g1793 ( .A(n_1053), .Y(n_1793) );
INVx4_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_1057), .A2(n_1058), .B1(n_1060), .B2(n_1061), .Y(n_1056) );
OAI221xp5_ASAP7_75t_L g1095 ( .A1(n_1058), .A2(n_1061), .B1(n_1096), .B2(n_1097), .C(n_1098), .Y(n_1095) );
OAI221xp5_ASAP7_75t_L g1479 ( .A1(n_1058), .A2(n_1480), .B1(n_1481), .B2(n_1482), .C(n_1483), .Y(n_1479) );
INVx2_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
INVx2_ASAP7_75t_SL g1803 ( .A(n_1059), .Y(n_1803) );
OAI22xp33_ASAP7_75t_L g1784 ( .A1(n_1061), .A2(n_1785), .B1(n_1786), .B2(n_1790), .Y(n_1784) );
INVx5_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
AOI21xp5_ASAP7_75t_L g1397 ( .A1(n_1063), .A2(n_1398), .B(n_1412), .Y(n_1397) );
INVx2_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1064), .Y(n_1376) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1068), .Y(n_1152) );
XNOR2x1_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1115), .Y(n_1068) );
NAND3xp33_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1089), .C(n_1092), .Y(n_1070) );
NOR3xp33_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1086), .C(n_1088), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1076), .Y(n_1072) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
NOR3xp33_ASAP7_75t_L g1454 ( .A(n_1088), .B(n_1455), .C(n_1464), .Y(n_1454) );
NOR3xp33_ASAP7_75t_L g1487 ( .A(n_1088), .B(n_1488), .C(n_1499), .Y(n_1487) );
OAI21xp5_ASAP7_75t_L g1092 ( .A1(n_1093), .A2(n_1102), .B(n_1114), .Y(n_1092) );
BUFx2_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
INVx2_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
INVx2_ASAP7_75t_L g1231 ( .A(n_1101), .Y(n_1231) );
INVx2_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
AOI21xp5_ASAP7_75t_SL g1179 ( .A1(n_1114), .A2(n_1180), .B(n_1200), .Y(n_1179) );
O2A1O1Ixp5_ASAP7_75t_L g1267 ( .A1(n_1114), .A2(n_1268), .B(n_1280), .C(n_1289), .Y(n_1267) );
OAI21xp5_ASAP7_75t_L g1436 ( .A1(n_1114), .A2(n_1437), .B(n_1444), .Y(n_1436) );
OAI21xp5_ASAP7_75t_L g1503 ( .A1(n_1114), .A2(n_1504), .B(n_1513), .Y(n_1503) );
AND3x1_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1124), .C(n_1127), .Y(n_1120) );
INVx2_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
OAI21xp5_ASAP7_75t_L g1137 ( .A1(n_1138), .A2(n_1145), .B(n_1151), .Y(n_1137) );
INVx2_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx2_ASAP7_75t_L g1518 ( .A(n_1142), .Y(n_1518) );
INVxp67_ASAP7_75t_SL g1154 ( .A(n_1155), .Y(n_1154) );
AOI22xp5_ASAP7_75t_L g1155 ( .A1(n_1156), .A2(n_1157), .B1(n_1295), .B2(n_1520), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
HB1xp67_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
XNOR2xp5_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1251), .Y(n_1158) );
OAI22x1_ASAP7_75t_L g1159 ( .A1(n_1160), .A2(n_1161), .B1(n_1204), .B2(n_1250), .Y(n_1159) );
INVx2_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
XNOR2x1_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1163), .Y(n_1161) );
AND3x2_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1179), .C(n_1202), .Y(n_1163) );
NOR2xp33_ASAP7_75t_SL g1164 ( .A(n_1165), .B(n_1173), .Y(n_1164) );
OAI21xp5_ASAP7_75t_SL g1165 ( .A1(n_1166), .A2(n_1167), .B(n_1170), .Y(n_1165) );
NAND3xp33_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1184), .C(n_1190), .Y(n_1180) );
AOI31xp33_ASAP7_75t_L g1190 ( .A1(n_1191), .A2(n_1192), .A3(n_1195), .B(n_1196), .Y(n_1190) );
INVx2_ASAP7_75t_SL g1193 ( .A(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1198), .Y(n_1411) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1204), .Y(n_1250) );
NAND3xp33_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1220), .C(n_1223), .Y(n_1205) );
NOR3xp33_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1218), .C(n_1219), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1211), .Y(n_1207) );
OAI21xp5_ASAP7_75t_L g1223 ( .A1(n_1224), .A2(n_1240), .B(n_1248), .Y(n_1223) );
BUFx2_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1228), .Y(n_1473) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
HB1xp67_ASAP7_75t_L g1507 ( .A(n_1231), .Y(n_1507) );
AOI22xp33_ASAP7_75t_L g1475 ( .A1(n_1238), .A2(n_1401), .B1(n_1476), .B2(n_1477), .Y(n_1475) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1242), .B(n_1245), .Y(n_1241) );
OAI21xp5_ASAP7_75t_L g1468 ( .A1(n_1248), .A2(n_1469), .B(n_1478), .Y(n_1468) );
INVx2_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
XOR2x2_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1294), .Y(n_1251) );
NAND3x1_ASAP7_75t_SL g1252 ( .A(n_1253), .B(n_1267), .C(n_1292), .Y(n_1252) );
HB1xp67_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1295), .Y(n_1520) );
XOR2xp5_ASAP7_75t_L g1295 ( .A(n_1296), .B(n_1377), .Y(n_1295) );
HB1xp67_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
XNOR2x2_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1341), .Y(n_1297) );
NAND3xp33_ASAP7_75t_L g1299 ( .A(n_1300), .B(n_1322), .C(n_1325), .Y(n_1299) );
OAI31xp33_ASAP7_75t_L g1300 ( .A1(n_1301), .A2(n_1307), .A3(n_1319), .B(n_1320), .Y(n_1300) );
NAND2xp5_ASAP7_75t_L g1301 ( .A(n_1302), .B(n_1304), .Y(n_1301) );
OAI211xp5_ASAP7_75t_L g1308 ( .A1(n_1309), .A2(n_1310), .B(n_1311), .C(n_1312), .Y(n_1308) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
NOR3xp33_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1339), .C(n_1340), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1330), .Y(n_1326) );
INVx2_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
NOR3xp33_ASAP7_75t_L g1420 ( .A(n_1340), .B(n_1421), .C(n_1432), .Y(n_1420) );
XNOR2x2_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1343), .Y(n_1341) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1359 ( .A(n_1360), .B(n_1363), .Y(n_1359) );
OAI21xp33_ASAP7_75t_L g1363 ( .A1(n_1364), .A2(n_1371), .B(n_1376), .Y(n_1363) );
OAI22xp5_ASAP7_75t_L g1377 ( .A1(n_1378), .A2(n_1449), .B1(n_1450), .B2(n_1519), .Y(n_1377) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1378), .Y(n_1519) );
XNOR2xp5_ASAP7_75t_L g1378 ( .A(n_1379), .B(n_1417), .Y(n_1378) );
OAI22xp5_ASAP7_75t_L g1379 ( .A1(n_1380), .A2(n_1414), .B1(n_1415), .B2(n_1416), .Y(n_1379) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1380), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_1381), .B(n_1397), .Y(n_1380) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
NAND3xp33_ASAP7_75t_L g1398 ( .A(n_1399), .B(n_1403), .C(n_1407), .Y(n_1398) );
CKINVDCx5p33_ASAP7_75t_R g1414 ( .A(n_1415), .Y(n_1414) );
INVx2_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
NAND3xp33_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1433), .C(n_1436), .Y(n_1419) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_1422), .B(n_1425), .Y(n_1421) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
OAI22xp5_ASAP7_75t_L g1450 ( .A1(n_1451), .A2(n_1452), .B1(n_1484), .B2(n_1485), .Y(n_1450) );
INVx2_ASAP7_75t_SL g1451 ( .A(n_1452), .Y(n_1451) );
NAND3xp33_ASAP7_75t_L g1453 ( .A(n_1454), .B(n_1465), .C(n_1468), .Y(n_1453) );
NAND2xp5_ASAP7_75t_L g1455 ( .A(n_1456), .B(n_1459), .Y(n_1455) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
NAND3xp33_ASAP7_75t_L g1486 ( .A(n_1487), .B(n_1500), .C(n_1503), .Y(n_1486) );
NAND2xp5_ASAP7_75t_L g1488 ( .A(n_1489), .B(n_1492), .Y(n_1488) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
OAI221xp5_ASAP7_75t_SL g1521 ( .A1(n_1522), .A2(n_1740), .B1(n_1743), .B2(n_1853), .C(n_1856), .Y(n_1521) );
AOI21xp5_ASAP7_75t_L g1522 ( .A1(n_1523), .A2(n_1664), .B(n_1712), .Y(n_1522) );
NAND5xp2_ASAP7_75t_L g1523 ( .A(n_1524), .B(n_1586), .C(n_1627), .D(n_1642), .E(n_1657), .Y(n_1523) );
AOI211xp5_ASAP7_75t_SL g1524 ( .A1(n_1525), .A2(n_1550), .B(n_1568), .C(n_1579), .Y(n_1524) );
AND2x2_ASAP7_75t_L g1525 ( .A(n_1526), .B(n_1541), .Y(n_1525) );
OR2x2_ASAP7_75t_L g1649 ( .A(n_1526), .B(n_1551), .Y(n_1649) );
A2O1A1Ixp33_ASAP7_75t_SL g1657 ( .A1(n_1526), .A2(n_1641), .B(n_1658), .C(n_1661), .Y(n_1657) );
INVx2_ASAP7_75t_L g1662 ( .A(n_1526), .Y(n_1662) );
NAND2xp5_ASAP7_75t_SL g1668 ( .A(n_1526), .B(n_1600), .Y(n_1668) );
NAND2xp5_ASAP7_75t_L g1684 ( .A(n_1526), .B(n_1685), .Y(n_1684) );
INVx2_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
INVx3_ASAP7_75t_L g1578 ( .A(n_1527), .Y(n_1578) );
NOR2xp33_ASAP7_75t_L g1602 ( .A(n_1527), .B(n_1554), .Y(n_1602) );
NOR2xp33_ASAP7_75t_L g1606 ( .A(n_1527), .B(n_1607), .Y(n_1606) );
AND2x2_ASAP7_75t_L g1610 ( .A(n_1527), .B(n_1554), .Y(n_1610) );
NAND2xp5_ASAP7_75t_L g1678 ( .A(n_1527), .B(n_1629), .Y(n_1678) );
AND2x2_ASAP7_75t_L g1705 ( .A(n_1527), .B(n_1569), .Y(n_1705) );
AND2x2_ASAP7_75t_L g1527 ( .A(n_1528), .B(n_1536), .Y(n_1527) );
AND2x4_ASAP7_75t_L g1529 ( .A(n_1530), .B(n_1531), .Y(n_1529) );
AND2x6_ASAP7_75t_L g1534 ( .A(n_1530), .B(n_1535), .Y(n_1534) );
AND2x6_ASAP7_75t_L g1537 ( .A(n_1530), .B(n_1538), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_1530), .B(n_1540), .Y(n_1539) );
AND2x2_ASAP7_75t_L g1548 ( .A(n_1530), .B(n_1540), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1556 ( .A(n_1530), .B(n_1540), .Y(n_1556) );
AND2x2_ASAP7_75t_L g1531 ( .A(n_1532), .B(n_1533), .Y(n_1531) );
INVx2_ASAP7_75t_L g1742 ( .A(n_1534), .Y(n_1742) );
HB1xp67_ASAP7_75t_L g1923 ( .A(n_1535), .Y(n_1923) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1542), .Y(n_1541) );
OR2x2_ASAP7_75t_L g1588 ( .A(n_1542), .B(n_1569), .Y(n_1588) );
AOI21xp33_ASAP7_75t_L g1714 ( .A1(n_1542), .A2(n_1649), .B(n_1652), .Y(n_1714) );
OR2x2_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1546), .Y(n_1542) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1543), .Y(n_1577) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1543), .Y(n_1612) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1543), .Y(n_1629) );
AND2x2_ASAP7_75t_L g1673 ( .A(n_1543), .B(n_1546), .Y(n_1673) );
NAND2xp5_ASAP7_75t_L g1543 ( .A(n_1544), .B(n_1545), .Y(n_1543) );
OR2x2_ASAP7_75t_L g1585 ( .A(n_1546), .B(n_1577), .Y(n_1585) );
NAND2xp5_ASAP7_75t_L g1619 ( .A(n_1546), .B(n_1570), .Y(n_1619) );
AND2x2_ASAP7_75t_L g1641 ( .A(n_1546), .B(n_1569), .Y(n_1641) );
NAND2xp5_ASAP7_75t_L g1732 ( .A(n_1546), .B(n_1662), .Y(n_1732) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1547), .B(n_1549), .Y(n_1546) );
AND2x4_ASAP7_75t_L g1597 ( .A(n_1547), .B(n_1549), .Y(n_1597) );
NAND2xp5_ASAP7_75t_L g1550 ( .A(n_1551), .B(n_1565), .Y(n_1550) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1574 ( .A(n_1552), .B(n_1575), .Y(n_1574) );
AND2x2_ASAP7_75t_L g1552 ( .A(n_1553), .B(n_1558), .Y(n_1552) );
OR2x2_ASAP7_75t_L g1633 ( .A(n_1553), .B(n_1580), .Y(n_1633) );
AND2x2_ASAP7_75t_L g1645 ( .A(n_1553), .B(n_1646), .Y(n_1645) );
AND2x2_ASAP7_75t_L g1660 ( .A(n_1553), .B(n_1600), .Y(n_1660) );
AND2x2_ASAP7_75t_L g1663 ( .A(n_1553), .B(n_1621), .Y(n_1663) );
OR2x2_ASAP7_75t_L g1667 ( .A(n_1553), .B(n_1668), .Y(n_1667) );
AOI321xp33_ASAP7_75t_L g1697 ( .A1(n_1553), .A2(n_1698), .A3(n_1699), .B1(n_1700), .B2(n_1702), .C(n_1703), .Y(n_1697) );
AND2x2_ASAP7_75t_L g1723 ( .A(n_1553), .B(n_1628), .Y(n_1723) );
AND2x2_ASAP7_75t_L g1728 ( .A(n_1553), .B(n_1729), .Y(n_1728) );
CKINVDCx5p33_ASAP7_75t_R g1553 ( .A(n_1554), .Y(n_1553) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_1554), .B(n_1567), .Y(n_1566) );
AND2x2_ASAP7_75t_L g1624 ( .A(n_1554), .B(n_1625), .Y(n_1624) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1554), .B(n_1558), .Y(n_1685) );
OR2x2_ASAP7_75t_L g1691 ( .A(n_1554), .B(n_1626), .Y(n_1691) );
NAND2xp5_ASAP7_75t_L g1701 ( .A(n_1554), .B(n_1646), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1554 ( .A(n_1555), .B(n_1557), .Y(n_1554) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1555), .B(n_1557), .Y(n_1591) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1558), .Y(n_1607) );
NAND2xp5_ASAP7_75t_L g1721 ( .A(n_1558), .B(n_1662), .Y(n_1721) );
AND2x2_ASAP7_75t_L g1558 ( .A(n_1559), .B(n_1562), .Y(n_1558) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1559), .Y(n_1582) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1559), .Y(n_1646) );
NAND2xp5_ASAP7_75t_L g1559 ( .A(n_1560), .B(n_1561), .Y(n_1559) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1562), .Y(n_1567) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1562), .B(n_1582), .Y(n_1581) );
OR2x2_ASAP7_75t_L g1601 ( .A(n_1562), .B(n_1582), .Y(n_1601) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1562), .Y(n_1626) );
NAND2xp5_ASAP7_75t_L g1562 ( .A(n_1563), .B(n_1564), .Y(n_1562) );
CKINVDCx14_ASAP7_75t_R g1565 ( .A(n_1566), .Y(n_1565) );
A2O1A1Ixp33_ASAP7_75t_L g1713 ( .A1(n_1566), .A2(n_1656), .B(n_1698), .C(n_1714), .Y(n_1713) );
AND2x2_ASAP7_75t_L g1621 ( .A(n_1567), .B(n_1582), .Y(n_1621) );
NOR2xp33_ASAP7_75t_L g1568 ( .A(n_1569), .B(n_1573), .Y(n_1568) );
INVx3_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1570), .B(n_1605), .Y(n_1604) );
NOR2xp33_ASAP7_75t_L g1636 ( .A(n_1570), .B(n_1611), .Y(n_1636) );
INVx3_ASAP7_75t_L g1656 ( .A(n_1570), .Y(n_1656) );
AND2x2_ASAP7_75t_L g1686 ( .A(n_1570), .B(n_1629), .Y(n_1686) );
OR2x2_ASAP7_75t_L g1688 ( .A(n_1570), .B(n_1585), .Y(n_1688) );
AND2x2_ASAP7_75t_L g1696 ( .A(n_1570), .B(n_1611), .Y(n_1696) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1570), .B(n_1584), .Y(n_1702) );
AND2x2_ASAP7_75t_L g1727 ( .A(n_1570), .B(n_1673), .Y(n_1727) );
AND2x4_ASAP7_75t_SL g1570 ( .A(n_1571), .B(n_1572), .Y(n_1570) );
INVxp67_ASAP7_75t_L g1573 ( .A(n_1574), .Y(n_1573) );
AOI221xp5_ASAP7_75t_L g1665 ( .A1(n_1574), .A2(n_1585), .B1(n_1641), .B2(n_1666), .C(n_1671), .Y(n_1665) );
OAI21xp33_ASAP7_75t_L g1617 ( .A1(n_1575), .A2(n_1618), .B(n_1620), .Y(n_1617) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
NAND2xp5_ASAP7_75t_L g1576 ( .A(n_1577), .B(n_1578), .Y(n_1576) );
AND2x2_ASAP7_75t_L g1596 ( .A(n_1577), .B(n_1597), .Y(n_1596) );
NAND2xp5_ASAP7_75t_L g1583 ( .A(n_1578), .B(n_1584), .Y(n_1583) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1578), .Y(n_1593) );
NOR2xp33_ASAP7_75t_L g1628 ( .A(n_1578), .B(n_1601), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1578), .B(n_1581), .Y(n_1638) );
O2A1O1Ixp33_ASAP7_75t_L g1737 ( .A1(n_1578), .A2(n_1588), .B(n_1738), .C(n_1739), .Y(n_1737) );
NOR2xp33_ASAP7_75t_L g1579 ( .A(n_1580), .B(n_1583), .Y(n_1579) );
OR2x2_ASAP7_75t_L g1717 ( .A(n_1580), .B(n_1591), .Y(n_1717) );
INVx1_ASAP7_75t_L g1580 ( .A(n_1581), .Y(n_1580) );
NAND2xp5_ASAP7_75t_L g1592 ( .A(n_1581), .B(n_1593), .Y(n_1592) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_1581), .B(n_1602), .Y(n_1675) );
NAND3xp33_ASAP7_75t_L g1679 ( .A(n_1581), .B(n_1605), .C(n_1680), .Y(n_1679) );
AND2x2_ASAP7_75t_L g1734 ( .A(n_1581), .B(n_1610), .Y(n_1734) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1582), .Y(n_1729) );
NOR2xp33_ASAP7_75t_L g1622 ( .A(n_1583), .B(n_1623), .Y(n_1622) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1583), .Y(n_1648) );
AND2x2_ASAP7_75t_L g1698 ( .A(n_1584), .B(n_1593), .Y(n_1698) );
INVx2_ASAP7_75t_SL g1584 ( .A(n_1585), .Y(n_1584) );
AOI211xp5_ASAP7_75t_L g1586 ( .A1(n_1587), .A2(n_1589), .B(n_1594), .C(n_1622), .Y(n_1586) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
OR2x2_ASAP7_75t_L g1590 ( .A(n_1591), .B(n_1592), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_1591), .B(n_1621), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1653 ( .A(n_1591), .B(n_1600), .Y(n_1653) );
AOI32xp33_ASAP7_75t_L g1704 ( .A1(n_1591), .A2(n_1636), .A3(n_1705), .B1(n_1706), .B2(n_1708), .Y(n_1704) );
OAI211xp5_ASAP7_75t_L g1703 ( .A1(n_1592), .A2(n_1695), .B(n_1704), .C(n_1709), .Y(n_1703) );
AND2x2_ASAP7_75t_L g1680 ( .A(n_1593), .B(n_1681), .Y(n_1680) );
AND2x2_ASAP7_75t_L g1708 ( .A(n_1593), .B(n_1621), .Y(n_1708) );
OAI211xp5_ASAP7_75t_SL g1594 ( .A1(n_1595), .A2(n_1598), .B(n_1603), .C(n_1617), .Y(n_1594) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1596), .Y(n_1595) );
AOI221xp5_ASAP7_75t_L g1722 ( .A1(n_1596), .A2(n_1661), .B1(n_1702), .B2(n_1723), .C(n_1724), .Y(n_1722) );
INVx2_ASAP7_75t_L g1605 ( .A(n_1597), .Y(n_1605) );
CKINVDCx6p67_ASAP7_75t_R g1655 ( .A(n_1597), .Y(n_1655) );
NAND2xp5_ASAP7_75t_L g1676 ( .A(n_1597), .B(n_1677), .Y(n_1676) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1599), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1600), .B(n_1602), .Y(n_1599) );
NAND2xp5_ASAP7_75t_L g1609 ( .A(n_1600), .B(n_1610), .Y(n_1609) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1601), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1670 ( .A(n_1602), .B(n_1621), .Y(n_1670) );
INVx1_ASAP7_75t_L g1725 ( .A(n_1602), .Y(n_1725) );
AOI221xp5_ASAP7_75t_L g1603 ( .A1(n_1604), .A2(n_1606), .B1(n_1608), .B2(n_1611), .C(n_1613), .Y(n_1603) );
OAI22xp5_ASAP7_75t_L g1630 ( .A1(n_1604), .A2(n_1605), .B1(n_1631), .B2(n_1633), .Y(n_1630) );
INVx1_ASAP7_75t_L g1692 ( .A(n_1604), .Y(n_1692) );
OAI22xp5_ASAP7_75t_L g1666 ( .A1(n_1605), .A2(n_1654), .B1(n_1667), .B2(n_1669), .Y(n_1666) );
INVx1_ASAP7_75t_L g1739 ( .A(n_1606), .Y(n_1739) );
OAI22xp5_ASAP7_75t_L g1634 ( .A1(n_1607), .A2(n_1635), .B1(n_1637), .B2(n_1639), .Y(n_1634) );
NAND2xp5_ASAP7_75t_L g1706 ( .A(n_1607), .B(n_1707), .Y(n_1706) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1609), .Y(n_1608) );
NAND2xp5_ASAP7_75t_L g1632 ( .A(n_1609), .B(n_1629), .Y(n_1632) );
AND2x2_ASAP7_75t_L g1640 ( .A(n_1611), .B(n_1641), .Y(n_1640) );
AND2x2_ASAP7_75t_L g1733 ( .A(n_1611), .B(n_1734), .Y(n_1733) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1614), .Y(n_1613) );
INVx1_ASAP7_75t_L g1711 ( .A(n_1614), .Y(n_1711) );
AND2x2_ASAP7_75t_L g1614 ( .A(n_1615), .B(n_1616), .Y(n_1614) );
O2A1O1Ixp33_ASAP7_75t_L g1735 ( .A1(n_1618), .A2(n_1675), .B(n_1736), .C(n_1737), .Y(n_1735) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1619), .Y(n_1618) );
INVx1_ASAP7_75t_L g1738 ( .A(n_1620), .Y(n_1738) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1621), .Y(n_1707) );
NAND2xp5_ASAP7_75t_L g1658 ( .A(n_1623), .B(n_1659), .Y(n_1658) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
A2O1A1Ixp33_ASAP7_75t_L g1730 ( .A1(n_1624), .A2(n_1699), .B(n_1731), .C(n_1733), .Y(n_1730) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1626), .Y(n_1625) );
O2A1O1Ixp33_ASAP7_75t_L g1627 ( .A1(n_1628), .A2(n_1629), .B(n_1630), .C(n_1634), .Y(n_1627) );
NAND2xp5_ASAP7_75t_L g1651 ( .A(n_1628), .B(n_1629), .Y(n_1651) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1629), .Y(n_1681) );
INVxp67_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
NOR2xp33_ASAP7_75t_L g1694 ( .A(n_1633), .B(n_1695), .Y(n_1694) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
AOI21xp33_ASAP7_75t_L g1719 ( .A1(n_1639), .A2(n_1720), .B(n_1721), .Y(n_1719) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
AOI221xp5_ASAP7_75t_L g1715 ( .A1(n_1641), .A2(n_1677), .B1(n_1716), .B2(n_1718), .C(n_1719), .Y(n_1715) );
OAI21xp33_ASAP7_75t_L g1642 ( .A1(n_1643), .A2(n_1650), .B(n_1656), .Y(n_1642) );
OAI21xp33_ASAP7_75t_L g1643 ( .A1(n_1644), .A2(n_1647), .B(n_1649), .Y(n_1643) );
NOR2xp33_ASAP7_75t_L g1677 ( .A(n_1644), .B(n_1678), .Y(n_1677) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1645), .Y(n_1644) );
INVxp67_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
AOI21xp33_ASAP7_75t_SL g1650 ( .A1(n_1651), .A2(n_1652), .B(n_1654), .Y(n_1650) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1651), .Y(n_1736) );
CKINVDCx5p33_ASAP7_75t_R g1652 ( .A(n_1653), .Y(n_1652) );
CKINVDCx6p67_ASAP7_75t_R g1654 ( .A(n_1655), .Y(n_1654) );
INVx2_ASAP7_75t_L g1699 ( .A(n_1656), .Y(n_1699) );
OAI221xp5_ASAP7_75t_L g1687 ( .A1(n_1659), .A2(n_1688), .B1(n_1689), .B2(n_1692), .C(n_1693), .Y(n_1687) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1660), .Y(n_1659) );
AND2x2_ASAP7_75t_L g1661 ( .A(n_1662), .B(n_1663), .Y(n_1661) );
NOR2xp33_ASAP7_75t_L g1690 ( .A(n_1662), .B(n_1691), .Y(n_1690) );
NAND3xp33_ASAP7_75t_L g1664 ( .A(n_1665), .B(n_1682), .C(n_1697), .Y(n_1664) );
AOI211xp5_ASAP7_75t_L g1724 ( .A1(n_1668), .A2(n_1725), .B(n_1726), .C(n_1728), .Y(n_1724) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1670), .Y(n_1669) );
OAI211xp5_ASAP7_75t_L g1671 ( .A1(n_1672), .A2(n_1674), .B(n_1676), .C(n_1679), .Y(n_1671) );
CKINVDCx14_ASAP7_75t_R g1672 ( .A(n_1673), .Y(n_1672) );
INVx1_ASAP7_75t_L g1674 ( .A(n_1675), .Y(n_1674) );
O2A1O1Ixp33_ASAP7_75t_L g1682 ( .A1(n_1675), .A2(n_1683), .B(n_1686), .C(n_1687), .Y(n_1682) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1685), .Y(n_1720) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1688), .Y(n_1718) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
INVxp67_ASAP7_75t_SL g1693 ( .A(n_1694), .Y(n_1693) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1696), .Y(n_1695) );
INVx1_ASAP7_75t_L g1700 ( .A(n_1701), .Y(n_1700) );
INVx1_ASAP7_75t_L g1709 ( .A(n_1710), .Y(n_1709) );
INVx1_ASAP7_75t_L g1710 ( .A(n_1711), .Y(n_1710) );
NAND5xp2_ASAP7_75t_SL g1712 ( .A(n_1713), .B(n_1715), .C(n_1722), .D(n_1730), .E(n_1735), .Y(n_1712) );
INVx1_ASAP7_75t_L g1716 ( .A(n_1717), .Y(n_1716) );
INVx1_ASAP7_75t_L g1726 ( .A(n_1727), .Y(n_1726) );
INVx1_ASAP7_75t_L g1731 ( .A(n_1732), .Y(n_1731) );
CKINVDCx20_ASAP7_75t_R g1740 ( .A(n_1741), .Y(n_1740) );
CKINVDCx20_ASAP7_75t_R g1741 ( .A(n_1742), .Y(n_1741) );
INVx1_ASAP7_75t_L g1851 ( .A(n_1744), .Y(n_1851) );
OAI211xp5_ASAP7_75t_L g1744 ( .A1(n_1745), .A2(n_1751), .B(n_1780), .C(n_1822), .Y(n_1744) );
CKINVDCx14_ASAP7_75t_R g1745 ( .A(n_1746), .Y(n_1745) );
AND2x4_ASAP7_75t_L g1746 ( .A(n_1747), .B(n_1749), .Y(n_1746) );
AND2x2_ASAP7_75t_SL g1907 ( .A(n_1747), .B(n_1749), .Y(n_1907) );
INVx1_ASAP7_75t_SL g1747 ( .A(n_1748), .Y(n_1747) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1750), .Y(n_1749) );
NOR3xp33_ASAP7_75t_SL g1751 ( .A(n_1752), .B(n_1759), .C(n_1774), .Y(n_1751) );
INVx2_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
INVx2_ASAP7_75t_SL g1754 ( .A(n_1755), .Y(n_1754) );
INVx1_ASAP7_75t_L g1905 ( .A(n_1755), .Y(n_1905) );
INVx1_ASAP7_75t_L g1756 ( .A(n_1757), .Y(n_1756) );
INVx1_ASAP7_75t_L g1906 ( .A(n_1757), .Y(n_1906) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
CKINVDCx8_ASAP7_75t_R g1762 ( .A(n_1763), .Y(n_1762) );
AOI22xp33_ASAP7_75t_L g1764 ( .A1(n_1765), .A2(n_1769), .B1(n_1770), .B2(n_1773), .Y(n_1764) );
AOI22xp33_ASAP7_75t_L g1900 ( .A1(n_1765), .A2(n_1770), .B1(n_1901), .B2(n_1902), .Y(n_1900) );
BUFx3_ASAP7_75t_L g1765 ( .A(n_1766), .Y(n_1765) );
AND2x2_ASAP7_75t_L g1766 ( .A(n_1767), .B(n_1768), .Y(n_1766) );
AND2x4_ASAP7_75t_L g1771 ( .A(n_1767), .B(n_1772), .Y(n_1771) );
AOI22xp33_ASAP7_75t_L g1829 ( .A1(n_1769), .A2(n_1830), .B1(n_1833), .B2(n_1834), .Y(n_1829) );
BUFx6f_ASAP7_75t_L g1770 ( .A(n_1771), .Y(n_1770) );
BUFx2_ASAP7_75t_L g1775 ( .A(n_1776), .Y(n_1775) );
INVx2_ASAP7_75t_SL g1897 ( .A(n_1776), .Y(n_1897) );
INVx1_ASAP7_75t_L g1777 ( .A(n_1778), .Y(n_1777) );
INVx2_ASAP7_75t_L g1898 ( .A(n_1778), .Y(n_1898) );
INVx2_ASAP7_75t_L g1778 ( .A(n_1779), .Y(n_1778) );
NOR2xp33_ASAP7_75t_L g1780 ( .A(n_1781), .B(n_1808), .Y(n_1780) );
OAI33xp33_ASAP7_75t_L g1781 ( .A1(n_1782), .A2(n_1784), .A3(n_1791), .B1(n_1796), .B2(n_1799), .B3(n_1802), .Y(n_1781) );
BUFx6f_ASAP7_75t_L g1782 ( .A(n_1783), .Y(n_1782) );
OAI22xp33_ASAP7_75t_L g1811 ( .A1(n_1785), .A2(n_1797), .B1(n_1812), .B2(n_1815), .Y(n_1811) );
INVx1_ASAP7_75t_L g1786 ( .A(n_1787), .Y(n_1786) );
INVx1_ASAP7_75t_L g1787 ( .A(n_1788), .Y(n_1787) );
INVx1_ASAP7_75t_L g1788 ( .A(n_1789), .Y(n_1788) );
OAI22xp5_ASAP7_75t_L g1791 ( .A1(n_1792), .A2(n_1793), .B1(n_1794), .B2(n_1795), .Y(n_1791) );
HB1xp67_ASAP7_75t_L g1870 ( .A(n_1795), .Y(n_1870) );
OAI33xp33_ASAP7_75t_L g1866 ( .A1(n_1799), .A2(n_1867), .A3(n_1871), .B1(n_1872), .B2(n_1877), .B3(n_1880), .Y(n_1866) );
INVx2_ASAP7_75t_L g1799 ( .A(n_1800), .Y(n_1799) );
INVx1_ASAP7_75t_L g1800 ( .A(n_1801), .Y(n_1800) );
OAI22xp5_ASAP7_75t_L g1802 ( .A1(n_1803), .A2(n_1804), .B1(n_1805), .B2(n_1807), .Y(n_1802) );
BUFx3_ASAP7_75t_L g1805 ( .A(n_1806), .Y(n_1805) );
OAI33xp33_ASAP7_75t_L g1808 ( .A1(n_1809), .A2(n_1811), .A3(n_1817), .B1(n_1818), .B2(n_1820), .B3(n_1821), .Y(n_1808) );
BUFx3_ASAP7_75t_L g1809 ( .A(n_1810), .Y(n_1809) );
INVx2_ASAP7_75t_L g1812 ( .A(n_1813), .Y(n_1812) );
INVx1_ASAP7_75t_L g1813 ( .A(n_1814), .Y(n_1813) );
HB1xp67_ASAP7_75t_L g1815 ( .A(n_1816), .Y(n_1815) );
INVx1_ASAP7_75t_L g1887 ( .A(n_1816), .Y(n_1887) );
OAI31xp33_ASAP7_75t_L g1822 ( .A1(n_1823), .A2(n_1837), .A3(n_1845), .B(n_1848), .Y(n_1822) );
BUFx2_ASAP7_75t_L g1824 ( .A(n_1825), .Y(n_1824) );
INVx3_ASAP7_75t_L g1826 ( .A(n_1827), .Y(n_1826) );
AOI22xp33_ASAP7_75t_L g1919 ( .A1(n_1830), .A2(n_1834), .B1(n_1901), .B2(n_1920), .Y(n_1919) );
BUFx3_ASAP7_75t_L g1830 ( .A(n_1831), .Y(n_1830) );
INVx2_ASAP7_75t_L g1834 ( .A(n_1835), .Y(n_1834) );
INVx2_ASAP7_75t_L g1835 ( .A(n_1836), .Y(n_1835) );
INVx1_ASAP7_75t_L g1838 ( .A(n_1839), .Y(n_1838) );
INVx1_ASAP7_75t_L g1839 ( .A(n_1840), .Y(n_1839) );
HB1xp67_ASAP7_75t_L g1913 ( .A(n_1840), .Y(n_1913) );
HB1xp67_ASAP7_75t_L g1842 ( .A(n_1843), .Y(n_1842) );
BUFx2_ASAP7_75t_L g1843 ( .A(n_1844), .Y(n_1843) );
INVx1_ASAP7_75t_L g1917 ( .A(n_1844), .Y(n_1917) );
CKINVDCx16_ASAP7_75t_R g1846 ( .A(n_1847), .Y(n_1846) );
INVx3_ASAP7_75t_SL g1911 ( .A(n_1847), .Y(n_1911) );
OAI31xp33_ASAP7_75t_SL g1908 ( .A1(n_1848), .A2(n_1909), .A3(n_1912), .B(n_1918), .Y(n_1908) );
BUFx3_ASAP7_75t_L g1848 ( .A(n_1849), .Y(n_1848) );
INVx3_ASAP7_75t_L g1853 ( .A(n_1854), .Y(n_1853) );
HB1xp67_ASAP7_75t_L g1857 ( .A(n_1858), .Y(n_1857) );
BUFx3_ASAP7_75t_L g1858 ( .A(n_1859), .Y(n_1858) );
INVxp33_ASAP7_75t_SL g1860 ( .A(n_1861), .Y(n_1860) );
INVx1_ASAP7_75t_L g1862 ( .A(n_1863), .Y(n_1862) );
HB1xp67_ASAP7_75t_L g1863 ( .A(n_1864), .Y(n_1863) );
NAND3xp33_ASAP7_75t_L g1864 ( .A(n_1865), .B(n_1894), .C(n_1908), .Y(n_1864) );
NOR2xp33_ASAP7_75t_L g1865 ( .A(n_1866), .B(n_1883), .Y(n_1865) );
OAI22xp5_ASAP7_75t_L g1889 ( .A1(n_1869), .A2(n_1879), .B1(n_1890), .B2(n_1891), .Y(n_1889) );
OAI22xp33_ASAP7_75t_L g1884 ( .A1(n_1873), .A2(n_1881), .B1(n_1885), .B2(n_1886), .Y(n_1884) );
INVx2_ASAP7_75t_L g1875 ( .A(n_1876), .Y(n_1875) );
INVx2_ASAP7_75t_SL g1886 ( .A(n_1887), .Y(n_1886) );
BUFx6f_ASAP7_75t_L g1891 ( .A(n_1892), .Y(n_1891) );
OAI31xp33_ASAP7_75t_L g1894 ( .A1(n_1895), .A2(n_1899), .A3(n_1903), .B(n_1907), .Y(n_1894) );
INVx1_ASAP7_75t_L g1896 ( .A(n_1897), .Y(n_1896) );
INVx1_ASAP7_75t_L g1904 ( .A(n_1905), .Y(n_1904) );
INVx2_ASAP7_75t_L g1914 ( .A(n_1915), .Y(n_1914) );
INVx2_ASAP7_75t_L g1915 ( .A(n_1916), .Y(n_1915) );
INVx2_ASAP7_75t_L g1916 ( .A(n_1917), .Y(n_1916) );
HB1xp67_ASAP7_75t_L g1921 ( .A(n_1922), .Y(n_1921) );
OAI21xp5_ASAP7_75t_L g1922 ( .A1(n_1923), .A2(n_1924), .B(n_1925), .Y(n_1922) );
INVx1_ASAP7_75t_L g1925 ( .A(n_1926), .Y(n_1925) );
endmodule