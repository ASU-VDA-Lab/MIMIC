module fake_jpeg_13833_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_2),
.B(n_9),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_51),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_52),
.B(n_53),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_28),
.Y(n_56)
);

CKINVDCx12_ASAP7_75t_R g133 ( 
.A(n_56),
.Y(n_133)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_59),
.B(n_60),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_61),
.B(n_66),
.Y(n_146)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_63),
.Y(n_152)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_1),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_69),
.B(n_70),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_32),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_21),
.B(n_1),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_73),
.B(n_76),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_24),
.B(n_4),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_96),
.Y(n_118)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_32),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_34),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_82),
.B(n_93),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx5_ASAP7_75t_SL g122 ( 
.A(n_86),
.Y(n_122)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_16),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_41),
.B(n_6),
.Y(n_93)
);

INVx6_ASAP7_75t_SL g94 ( 
.A(n_34),
.Y(n_94)
);

INVx5_ASAP7_75t_SL g153 ( 
.A(n_94),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_95),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_43),
.B(n_10),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_16),
.B(n_14),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_100),
.B(n_101),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_27),
.B(n_35),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_49),
.B(n_12),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_102),
.B(n_13),
.Y(n_138)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_73),
.A2(n_49),
.B(n_39),
.C(n_42),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_123),
.B(n_138),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_64),
.A2(n_35),
.B(n_47),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_142),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_53),
.B(n_39),
.C(n_47),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_54),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_64),
.A2(n_42),
.B(n_13),
.Y(n_132)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_141),
.B(n_58),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_62),
.A2(n_19),
.B1(n_48),
.B2(n_33),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_19),
.B1(n_48),
.B2(n_81),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_88),
.A2(n_91),
.B1(n_72),
.B2(n_84),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_54),
.B(n_19),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_85),
.B(n_29),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_155),
.B(n_30),
.Y(n_196)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_157),
.Y(n_231)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_192),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_108),
.B(n_70),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_163),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_166),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_46),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_174),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_68),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_168),
.B(n_170),
.Y(n_229)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_169),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_77),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_171),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_150),
.A2(n_60),
.B1(n_33),
.B2(n_103),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_172),
.A2(n_133),
.B1(n_106),
.B2(n_143),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_114),
.B(n_120),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_178),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_120),
.B(n_80),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_85),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_179),
.B(n_191),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_58),
.B(n_99),
.C(n_51),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_180),
.A2(n_145),
.B(n_105),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_136),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_183),
.Y(n_207)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_136),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_187),
.Y(n_223)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_111),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_185),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_186),
.Y(n_228)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_129),
.B(n_46),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_189),
.Y(n_224)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

NAND2xp33_ASAP7_75t_SL g190 ( 
.A(n_130),
.B(n_63),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_190),
.A2(n_198),
.B(n_145),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_46),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_147),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_196),
.B(n_113),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_124),
.B(n_95),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_199),
.C(n_139),
.Y(n_208)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

AO22x1_ASAP7_75t_L g205 ( 
.A1(n_195),
.A2(n_197),
.B1(n_152),
.B2(n_122),
.Y(n_205)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_129),
.B(n_30),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_141),
.A2(n_55),
.B1(n_86),
.B2(n_137),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_200),
.A2(n_171),
.B1(n_168),
.B2(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_135),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_215),
.B1(n_222),
.B2(n_179),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_109),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_218),
.A2(n_180),
.B(n_165),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_173),
.A2(n_116),
.B1(n_149),
.B2(n_110),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_219),
.A2(n_232),
.B1(n_182),
.B2(n_185),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_190),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_186),
.A2(n_149),
.B1(n_128),
.B2(n_115),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_173),
.A2(n_113),
.B1(n_143),
.B2(n_127),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_238),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_SL g266 ( 
.A1(n_235),
.A2(n_249),
.B(n_232),
.C(n_205),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_236),
.A2(n_240),
.B1(n_254),
.B2(n_205),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_206),
.B(n_189),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_237),
.B(n_242),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_173),
.B1(n_179),
.B2(n_194),
.Y(n_240)
);

AND2x6_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_202),
.Y(n_241)
);

AOI322xp5_ASAP7_75t_L g268 ( 
.A1(n_241),
.A2(n_243),
.A3(n_244),
.B1(n_247),
.B2(n_240),
.C1(n_254),
.C2(n_255),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_191),
.Y(n_242)
);

A2O1A1O1Ixp25_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_233),
.B(n_249),
.C(n_221),
.D(n_246),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_229),
.A2(n_177),
.B1(n_192),
.B2(n_169),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_245),
.Y(n_259)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_157),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_253),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_218),
.A2(n_187),
.B1(n_158),
.B2(n_166),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_251),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_248),
.B(n_255),
.Y(n_271)
);

AO21x1_ASAP7_75t_L g249 ( 
.A1(n_219),
.A2(n_201),
.B(n_217),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_227),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_227),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_212),
.A2(n_164),
.B1(n_195),
.B2(n_197),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_184),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_252),
.B(n_213),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_184),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_212),
.A2(n_163),
.B1(n_175),
.B2(n_147),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_214),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_268),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_258),
.B(n_265),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

OAI32xp33_ASAP7_75t_L g263 ( 
.A1(n_233),
.A2(n_207),
.A3(n_208),
.B1(n_214),
.B2(n_224),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_255),
.Y(n_273)
);

NAND3xp33_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_270),
.C(n_239),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_223),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_266),
.A2(n_236),
.B1(n_245),
.B2(n_251),
.Y(n_281)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

A2O1A1O1Ixp25_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_226),
.B(n_223),
.C(n_204),
.D(n_220),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_273),
.B(n_223),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_274),
.A2(n_282),
.B1(n_256),
.B2(n_263),
.Y(n_288)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_283),
.B1(n_272),
.B2(n_266),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_238),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_259),
.A2(n_209),
.B1(n_222),
.B2(n_226),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_284),
.Y(n_286)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_280),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_287),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_290),
.B(n_294),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_273),
.A2(n_258),
.B(n_259),
.Y(n_290)
);

AOI21x1_ASAP7_75t_SL g291 ( 
.A1(n_275),
.A2(n_272),
.B(n_266),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_291),
.A2(n_295),
.B1(n_283),
.B2(n_225),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_293),
.A2(n_281),
.B1(n_284),
.B2(n_275),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_278),
.A2(n_266),
.B(n_271),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_271),
.B1(n_209),
.B2(n_257),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_285),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_277),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_298),
.B(n_302),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_301),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_276),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g303 ( 
.A(n_287),
.B(n_279),
.CI(n_276),
.CON(n_303),
.SN(n_303)
);

OA21x2_ASAP7_75t_SL g307 ( 
.A1(n_303),
.A2(n_296),
.B(n_292),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_304),
.A2(n_291),
.B(n_292),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_294),
.B(n_293),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_308),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_300),
.Y(n_311)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_303),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_310),
.Y(n_312)
);

OAI21x1_ASAP7_75t_SL g316 ( 
.A1(n_311),
.A2(n_298),
.B(n_286),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_309),
.B(n_302),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_313),
.A2(n_306),
.B1(n_305),
.B2(n_304),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_317),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_316),
.A2(n_310),
.B(n_314),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_312),
.A2(n_297),
.B1(n_303),
.B2(n_286),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_317),
.Y(n_318)
);

AOI322xp5_ASAP7_75t_L g322 ( 
.A1(n_318),
.A2(n_319),
.A3(n_225),
.B1(n_230),
.B2(n_231),
.C1(n_289),
.C2(n_317),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_289),
.B(n_301),
.C(n_220),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_321),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_322),
.Y(n_324)
);


endmodule