module fake_netlist_1_8317_n_709 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_709);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_709;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_17), .Y(n_78) );
INVxp67_ASAP7_75t_SL g79 ( .A(n_30), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_40), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_42), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_59), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_16), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_1), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_10), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_29), .Y(n_86) );
INVxp67_ASAP7_75t_L g87 ( .A(n_28), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_9), .Y(n_88) );
INVxp67_ASAP7_75t_L g89 ( .A(n_61), .Y(n_89) );
BUFx3_ASAP7_75t_L g90 ( .A(n_51), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_46), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_52), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_71), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_53), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_14), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_2), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_38), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_8), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_24), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_14), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_0), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_72), .Y(n_102) );
INVxp67_ASAP7_75t_L g103 ( .A(n_19), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_49), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_15), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_4), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_32), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_69), .Y(n_108) );
INVxp33_ASAP7_75t_L g109 ( .A(n_58), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_16), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_64), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_55), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_44), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_23), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_63), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_70), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_74), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_65), .Y(n_118) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_31), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_18), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_5), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g122 ( .A(n_43), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_60), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_36), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_37), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_111), .Y(n_126) );
INVx5_ASAP7_75t_L g127 ( .A(n_111), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_83), .B(n_0), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_80), .B(n_1), .Y(n_129) );
NOR2xp67_ASAP7_75t_L g130 ( .A(n_83), .B(n_2), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_122), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_78), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_78), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_125), .B(n_3), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_122), .B(n_3), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_80), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_109), .B(n_4), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_93), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_107), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_93), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_111), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_91), .B(n_5), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_91), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_117), .Y(n_146) );
AND2x2_ASAP7_75t_SL g147 ( .A(n_92), .B(n_97), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_100), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_100), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_108), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_125), .B(n_6), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_88), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_88), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_92), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_108), .B(n_6), .Y(n_155) );
INVx5_ASAP7_75t_L g156 ( .A(n_111), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_95), .B(n_7), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_97), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_99), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_99), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_102), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_124), .B(n_7), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_84), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_95), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_98), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_98), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_96), .Y(n_167) );
INVx6_ASAP7_75t_L g168 ( .A(n_115), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_126), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_147), .B(n_89), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_127), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_131), .B(n_87), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_127), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_163), .B(n_110), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_127), .Y(n_175) );
INVx1_ASAP7_75t_SL g176 ( .A(n_163), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_147), .B(n_106), .Y(n_177) );
OR2x2_ASAP7_75t_L g178 ( .A(n_131), .B(n_121), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_127), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_141), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_139), .B(n_110), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_128), .A2(n_105), .B1(n_101), .B2(n_85), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_167), .B(n_103), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_164), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_164), .Y(n_185) );
BUFx10_ASAP7_75t_L g186 ( .A(n_167), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_127), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_127), .Y(n_188) );
OR2x2_ASAP7_75t_L g189 ( .A(n_137), .B(n_101), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_164), .Y(n_190) );
INVx5_ASAP7_75t_L g191 ( .A(n_168), .Y(n_191) );
OR2x2_ASAP7_75t_L g192 ( .A(n_137), .B(n_105), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_165), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_132), .B(n_123), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_128), .B(n_115), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_165), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_132), .B(n_82), .Y(n_197) );
NAND3x1_ASAP7_75t_L g198 ( .A(n_139), .B(n_124), .C(n_120), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_128), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_165), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_168), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_156), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_156), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_138), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_138), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_168), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_152), .B(n_115), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_140), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_126), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_168), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_140), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_133), .B(n_94), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_153), .B(n_90), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_133), .B(n_104), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_134), .B(n_120), .Y(n_215) );
INVx4_ASAP7_75t_L g216 ( .A(n_157), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_157), .B(n_118), .Y(n_217) );
INVx1_ASAP7_75t_SL g218 ( .A(n_146), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_142), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_157), .A2(n_118), .B1(n_113), .B2(n_102), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_141), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_142), .Y(n_222) );
AND2x6_ASAP7_75t_L g223 ( .A(n_134), .B(n_113), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_135), .A2(n_90), .B1(n_116), .B2(n_112), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_150), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_150), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_135), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_145), .A2(n_116), .B1(n_112), .B2(n_114), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_156), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_156), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_145), .B(n_111), .Y(n_231) );
AND2x2_ASAP7_75t_SL g232 ( .A(n_154), .B(n_119), .Y(n_232) );
INVx2_ASAP7_75t_SL g233 ( .A(n_195), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_199), .A2(n_159), .B(n_154), .Y(n_234) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_176), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_206), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_216), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_227), .B(n_161), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_184), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_216), .Y(n_240) );
BUFx12f_ASAP7_75t_L g241 ( .A(n_186), .Y(n_241) );
OR2x6_ASAP7_75t_SL g242 ( .A(n_180), .B(n_158), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_227), .B(n_161), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_194), .B(n_158), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_184), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_197), .B(n_159), .Y(n_246) );
AND2x6_ASAP7_75t_L g247 ( .A(n_217), .B(n_160), .Y(n_247) );
INVx1_ASAP7_75t_SL g248 ( .A(n_218), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_186), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_212), .B(n_160), .Y(n_250) );
AOI211xp5_ASAP7_75t_L g251 ( .A1(n_170), .A2(n_166), .B(n_162), .C(n_136), .Y(n_251) );
AND2x6_ASAP7_75t_SL g252 ( .A(n_221), .B(n_151), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_232), .A2(n_144), .B1(n_155), .B2(n_129), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_214), .B(n_149), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_172), .B(n_148), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_213), .B(n_130), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_185), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_216), .B(n_81), .Y(n_258) );
BUFx12f_ASAP7_75t_L g259 ( .A(n_186), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_232), .A2(n_223), .B1(n_217), .B2(n_199), .Y(n_260) );
BUFx3_ASAP7_75t_L g261 ( .A(n_206), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_185), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_181), .B(n_79), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_190), .Y(n_264) );
INVxp67_ASAP7_75t_L g265 ( .A(n_178), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_213), .B(n_156), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_199), .B(n_156), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_232), .A2(n_143), .B1(n_126), .B2(n_10), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_183), .B(n_45), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_178), .Y(n_270) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_174), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_190), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_217), .B(n_126), .Y(n_273) );
OAI22xp5_ASAP7_75t_SL g274 ( .A1(n_180), .A2(n_8), .B1(n_9), .B2(n_11), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_181), .B(n_143), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_223), .A2(n_143), .B1(n_126), .B2(n_13), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_223), .A2(n_143), .B1(n_12), .B2(n_13), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_220), .B(n_143), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_193), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_174), .B(n_11), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_193), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_189), .B(n_12), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_196), .Y(n_283) );
INVxp67_ASAP7_75t_L g284 ( .A(n_189), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_223), .Y(n_285) );
NOR3xp33_ASAP7_75t_SL g286 ( .A(n_177), .B(n_15), .C(n_20), .Y(n_286) );
INVx2_ASAP7_75t_SL g287 ( .A(n_192), .Y(n_287) );
OAI21xp5_ASAP7_75t_L g288 ( .A1(n_196), .A2(n_200), .B(n_195), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_207), .B(n_21), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_210), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_200), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_204), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g293 ( .A1(n_198), .A2(n_22), .B1(n_25), .B2(n_26), .Y(n_293) );
INVx2_ASAP7_75t_SL g294 ( .A(n_192), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_207), .B(n_27), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_222), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_195), .B(n_33), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_223), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_195), .B(n_34), .Y(n_299) );
BUFx4f_ASAP7_75t_L g300 ( .A(n_223), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_260), .A2(n_198), .B1(n_182), .B2(n_226), .Y(n_301) );
INVx4_ASAP7_75t_L g302 ( .A(n_247), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_235), .B(n_208), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_L g304 ( .A1(n_284), .A2(n_215), .B(n_204), .C(n_226), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_300), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_L g306 ( .A1(n_244), .A2(n_219), .B(n_208), .C(n_225), .Y(n_306) );
INVxp67_ASAP7_75t_L g307 ( .A(n_247), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_300), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_237), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_SL g310 ( .A1(n_299), .A2(n_231), .B(n_225), .C(n_219), .Y(n_310) );
INVx1_ASAP7_75t_SL g311 ( .A(n_248), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_247), .B(n_223), .Y(n_312) );
INVx4_ASAP7_75t_L g313 ( .A(n_247), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_247), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_241), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_234), .A2(n_228), .B(n_224), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_280), .A2(n_222), .B1(n_205), .B2(n_211), .Y(n_317) );
NAND2x1p5_ASAP7_75t_L g318 ( .A(n_233), .B(n_222), .Y(n_318) );
INVxp67_ASAP7_75t_L g319 ( .A(n_247), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_287), .B(n_205), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_270), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_237), .Y(n_322) );
BUFx2_ASAP7_75t_SL g323 ( .A(n_294), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_265), .B(n_201), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_241), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_280), .A2(n_211), .B1(n_201), .B2(n_210), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_285), .B(n_201), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_280), .A2(n_230), .B1(n_229), .B2(n_171), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_298), .Y(n_329) );
OR2x6_ASAP7_75t_L g330 ( .A(n_259), .B(n_230), .Y(n_330) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_246), .A2(n_229), .B(n_203), .C(n_202), .Y(n_331) );
INVx4_ASAP7_75t_L g332 ( .A(n_259), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_285), .Y(n_333) );
OR2x6_ASAP7_75t_L g334 ( .A(n_282), .B(n_187), .Y(n_334) );
BUFx4f_ASAP7_75t_L g335 ( .A(n_263), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_250), .A2(n_187), .B(n_203), .Y(n_336) );
INVx6_ASAP7_75t_L g337 ( .A(n_236), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_233), .Y(n_338) );
BUFx2_ASAP7_75t_L g339 ( .A(n_242), .Y(n_339) );
OAI221xp5_ASAP7_75t_L g340 ( .A1(n_253), .A2(n_179), .B1(n_202), .B2(n_188), .C(n_171), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_249), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_249), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_275), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_237), .Y(n_344) );
NOR2x1_ASAP7_75t_L g345 ( .A(n_263), .B(n_188), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_245), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_240), .Y(n_347) );
OAI21x1_ASAP7_75t_L g348 ( .A1(n_288), .A2(n_179), .B(n_175), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_263), .A2(n_175), .B1(n_173), .B2(n_191), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_240), .Y(n_350) );
A2O1A1Ixp33_ASAP7_75t_L g351 ( .A1(n_255), .A2(n_173), .B(n_191), .C(n_209), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_262), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_346), .Y(n_353) );
AO31x2_ASAP7_75t_L g354 ( .A1(n_326), .A2(n_297), .A3(n_292), .B(n_295), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_348), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_352), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_335), .A2(n_271), .B1(n_258), .B2(n_268), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_302), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_331), .A2(n_299), .B(n_289), .Y(n_359) );
OAI21x1_ASAP7_75t_L g360 ( .A1(n_331), .A2(n_278), .B(n_293), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_303), .B(n_254), .Y(n_361) );
OAI21x1_ASAP7_75t_L g362 ( .A1(n_306), .A2(n_278), .B(n_238), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_343), .Y(n_363) );
AO21x2_ASAP7_75t_L g364 ( .A1(n_351), .A2(n_286), .B(n_256), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_317), .A2(n_251), .B1(n_291), .B2(n_272), .Y(n_365) );
BUFx3_ASAP7_75t_L g366 ( .A(n_302), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_335), .A2(n_258), .B1(n_240), .B2(n_274), .Y(n_367) );
OA21x2_ASAP7_75t_L g368 ( .A1(n_336), .A2(n_264), .B(n_281), .Y(n_368) );
OAI21x1_ASAP7_75t_L g369 ( .A1(n_306), .A2(n_243), .B(n_238), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_313), .Y(n_370) );
CKINVDCx10_ASAP7_75t_R g371 ( .A(n_330), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_320), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_301), .B(n_243), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_336), .A2(n_257), .B(n_239), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_326), .A2(n_269), .B(n_283), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_321), .A2(n_279), .B1(n_296), .B2(n_273), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_301), .A2(n_273), .B1(n_239), .B2(n_283), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_309), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_322), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_344), .Y(n_380) );
CKINVDCx12_ASAP7_75t_R g381 ( .A(n_330), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_350), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_311), .Y(n_383) );
AO32x2_ASAP7_75t_L g384 ( .A1(n_313), .A2(n_296), .A3(n_252), .B1(n_277), .B2(n_266), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_383), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_361), .B(n_311), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_374), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_367), .A2(n_339), .B1(n_323), .B2(n_334), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_363), .Y(n_389) );
AO21x2_ASAP7_75t_L g390 ( .A1(n_355), .A2(n_310), .B(n_316), .Y(n_390) );
AOI222xp33_ASAP7_75t_L g391 ( .A1(n_361), .A2(n_342), .B1(n_341), .B2(n_315), .C1(n_332), .C2(n_325), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g392 ( .A1(n_372), .A2(n_334), .B1(n_332), .B2(n_330), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_365), .A2(n_334), .B1(n_328), .B2(n_345), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_377), .A2(n_307), .B1(n_319), .B2(n_318), .Y(n_394) );
AOI22xp33_ASAP7_75t_SL g395 ( .A1(n_372), .A2(n_324), .B1(n_314), .B2(n_319), .Y(n_395) );
OA21x2_ASAP7_75t_L g396 ( .A1(n_355), .A2(n_316), .B(n_340), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_365), .A2(n_363), .B1(n_357), .B2(n_373), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_353), .A2(n_304), .B1(n_340), .B2(n_349), .C(n_338), .Y(n_398) );
OAI22xp33_ASAP7_75t_L g399 ( .A1(n_371), .A2(n_307), .B1(n_314), .B2(n_312), .Y(n_399) );
OA21x2_ASAP7_75t_L g400 ( .A1(n_355), .A2(n_276), .B(n_257), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_353), .Y(n_401) );
INVxp67_ASAP7_75t_L g402 ( .A(n_356), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_373), .A2(n_356), .B1(n_364), .B2(n_376), .Y(n_403) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_366), .Y(n_404) );
OAI22xp33_ASAP7_75t_L g405 ( .A1(n_371), .A2(n_312), .B1(n_318), .B2(n_329), .Y(n_405) );
INVxp67_ASAP7_75t_SL g406 ( .A(n_377), .Y(n_406) );
OAI21xp33_ASAP7_75t_SL g407 ( .A1(n_374), .A2(n_296), .B(n_347), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_368), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_358), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_379), .B(n_347), .Y(n_410) );
NOR2x1_ASAP7_75t_SL g411 ( .A(n_366), .B(n_305), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_379), .B(n_304), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_389), .B(n_378), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_404), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_397), .B(n_401), .Y(n_415) );
AO21x2_ASAP7_75t_L g416 ( .A1(n_387), .A2(n_375), .B(n_360), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_401), .B(n_378), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_386), .Y(n_418) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_403), .B(n_368), .C(n_382), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_389), .Y(n_420) );
INVx2_ASAP7_75t_SL g421 ( .A(n_404), .Y(n_421) );
OAI21xp5_ASAP7_75t_SL g422 ( .A1(n_391), .A2(n_358), .B(n_370), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_408), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_385), .B(n_354), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_408), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_387), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_396), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_412), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_410), .B(n_378), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_385), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_402), .Y(n_431) );
CKINVDCx11_ASAP7_75t_R g432 ( .A(n_409), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_410), .Y(n_433) );
INVxp67_ASAP7_75t_L g434 ( .A(n_411), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_396), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_406), .B(n_382), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_396), .B(n_354), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_393), .B(n_380), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_396), .Y(n_439) );
BUFx2_ASAP7_75t_SL g440 ( .A(n_404), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_393), .B(n_380), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_390), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_390), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_392), .B(n_384), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_390), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_404), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_404), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_407), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_431), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_418), .B(n_388), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_433), .B(n_405), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_437), .A2(n_407), .B(n_375), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_433), .B(n_354), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_431), .Y(n_454) );
AND2x4_ASAP7_75t_L g455 ( .A(n_428), .B(n_411), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_420), .B(n_398), .Y(n_456) );
NOR2xp67_ASAP7_75t_L g457 ( .A(n_434), .B(n_381), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_420), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_430), .B(n_354), .Y(n_459) );
OAI22xp33_ASAP7_75t_L g460 ( .A1(n_422), .A2(n_394), .B1(n_399), .B2(n_370), .Y(n_460) );
NOR2xp33_ASAP7_75t_SL g461 ( .A(n_434), .B(n_381), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_413), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_423), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_413), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_423), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_429), .B(n_354), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_417), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_429), .B(n_384), .Y(n_468) );
OAI31xp33_ASAP7_75t_L g469 ( .A1(n_422), .A2(n_366), .A3(n_384), .B(n_267), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_417), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_428), .A2(n_364), .B1(n_395), .B2(n_267), .C(n_384), .Y(n_471) );
INVx4_ASAP7_75t_L g472 ( .A(n_414), .Y(n_472) );
INVx4_ASAP7_75t_L g473 ( .A(n_414), .Y(n_473) );
AOI221xp5_ASAP7_75t_L g474 ( .A1(n_415), .A2(n_364), .B1(n_384), .B2(n_261), .C(n_290), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_423), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_425), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_425), .Y(n_477) );
OR2x6_ASAP7_75t_L g478 ( .A(n_440), .B(n_375), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_425), .Y(n_479) );
OR2x6_ASAP7_75t_L g480 ( .A(n_440), .B(n_368), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_446), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_417), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_424), .B(n_354), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_424), .B(n_368), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_414), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_427), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_417), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_427), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_444), .A2(n_364), .B1(n_360), .B2(n_369), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_432), .B(n_384), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_427), .Y(n_491) );
OR2x6_ASAP7_75t_L g492 ( .A(n_444), .B(n_362), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_436), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_415), .B(n_369), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_436), .B(n_369), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_438), .B(n_362), .Y(n_496) );
INVx3_ASAP7_75t_L g497 ( .A(n_447), .Y(n_497) );
NAND4xp25_ASAP7_75t_L g498 ( .A(n_438), .B(n_441), .C(n_419), .D(n_448), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_441), .B(n_359), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_426), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_486), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_478), .B(n_448), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_466), .B(n_439), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_466), .B(n_439), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_486), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_459), .B(n_437), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_453), .B(n_435), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_484), .B(n_435), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_458), .Y(n_509) );
NAND3xp33_ASAP7_75t_L g510 ( .A(n_469), .B(n_419), .C(n_445), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_460), .B(n_421), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_485), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_453), .B(n_435), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_493), .B(n_421), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_488), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_483), .B(n_426), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_495), .B(n_426), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_488), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_492), .B(n_445), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_463), .B(n_443), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_492), .B(n_443), .Y(n_521) );
INVx2_ASAP7_75t_SL g522 ( .A(n_481), .Y(n_522) );
OAI33xp33_ASAP7_75t_L g523 ( .A1(n_460), .A2(n_442), .A3(n_447), .B1(n_327), .B2(n_47), .B3(n_48), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_449), .B(n_447), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_492), .B(n_442), .Y(n_525) );
OAI33xp33_ASAP7_75t_L g526 ( .A1(n_454), .A2(n_35), .A3(n_39), .B1(n_41), .B2(n_50), .B3(n_54), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_491), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_491), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_463), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_475), .B(n_416), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_475), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_462), .B(n_416), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_476), .B(n_416), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_464), .B(n_416), .Y(n_534) );
BUFx3_ASAP7_75t_L g535 ( .A(n_481), .Y(n_535) );
INVxp67_ASAP7_75t_L g536 ( .A(n_461), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_476), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_477), .Y(n_538) );
NOR3xp33_ASAP7_75t_L g539 ( .A(n_490), .B(n_359), .C(n_290), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_477), .Y(n_540) );
INVxp67_ASAP7_75t_L g541 ( .A(n_455), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_465), .Y(n_542) );
OAI221xp5_ASAP7_75t_L g543 ( .A1(n_471), .A2(n_337), .B1(n_236), .B2(n_261), .C(n_329), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_450), .B(n_400), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_468), .B(n_400), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_496), .B(n_400), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_498), .A2(n_337), .B1(n_400), .B2(n_329), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_500), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_455), .A2(n_337), .B1(n_333), .B2(n_308), .Y(n_549) );
NAND5xp2_ASAP7_75t_L g550 ( .A(n_474), .B(n_56), .C(n_57), .D(n_62), .E(n_66), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_465), .Y(n_551) );
INVx4_ASAP7_75t_L g552 ( .A(n_480), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_455), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_478), .B(n_67), .Y(n_554) );
BUFx2_ASAP7_75t_L g555 ( .A(n_480), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_479), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_479), .B(n_68), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_480), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_467), .B(n_73), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_497), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_503), .B(n_499), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_503), .B(n_478), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_504), .B(n_456), .Y(n_563) );
INVx2_ASAP7_75t_SL g564 ( .A(n_535), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_502), .B(n_487), .Y(n_565) );
AOI32xp33_ASAP7_75t_L g566 ( .A1(n_512), .A2(n_451), .A3(n_473), .B1(n_472), .B2(n_489), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_504), .B(n_482), .Y(n_567) );
NAND2x1p5_ASAP7_75t_L g568 ( .A(n_554), .B(n_457), .Y(n_568) );
OR2x6_ASAP7_75t_L g569 ( .A(n_552), .B(n_452), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_509), .B(n_470), .Y(n_570) );
OR2x6_ASAP7_75t_L g571 ( .A(n_552), .B(n_473), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_507), .B(n_489), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_535), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_509), .B(n_494), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_522), .B(n_473), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_507), .B(n_497), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_548), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_513), .B(n_497), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_513), .B(n_472), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_501), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_506), .B(n_472), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_506), .B(n_75), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_522), .B(n_76), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_519), .B(n_77), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_514), .B(n_169), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_519), .B(n_521), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_501), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_521), .B(n_169), .Y(n_588) );
NAND2x1_ASAP7_75t_L g589 ( .A(n_552), .B(n_305), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_550), .A2(n_333), .B1(n_305), .B2(n_308), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_516), .B(n_169), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_516), .B(n_169), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_525), .B(n_169), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_525), .B(n_209), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_548), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_546), .B(n_209), .Y(n_596) );
OAI31xp33_ASAP7_75t_L g597 ( .A1(n_536), .A2(n_333), .A3(n_308), .B(n_191), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_508), .B(n_209), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_546), .B(n_209), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_505), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_551), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_524), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_545), .B(n_191), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_529), .B(n_191), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_545), .B(n_191), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_502), .B(n_558), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_529), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_508), .B(n_517), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_531), .B(n_538), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_531), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_537), .B(n_538), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_502), .B(n_558), .Y(n_612) );
INVx3_ASAP7_75t_L g613 ( .A(n_502), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_610), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_581), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_609), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_563), .B(n_511), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_581), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_573), .B(n_523), .Y(n_619) );
OAI221xp5_ASAP7_75t_L g620 ( .A1(n_566), .A2(n_555), .B1(n_547), .B2(n_541), .C(n_510), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_611), .Y(n_621) );
OAI221xp5_ASAP7_75t_SL g622 ( .A1(n_569), .A2(n_555), .B1(n_553), .B2(n_510), .C(n_539), .Y(n_622) );
AOI211xp5_ASAP7_75t_SL g623 ( .A1(n_582), .A2(n_554), .B(n_544), .C(n_534), .Y(n_623) );
INVxp33_ASAP7_75t_L g624 ( .A(n_568), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_572), .B(n_537), .Y(n_625) );
NAND4xp25_ASAP7_75t_L g626 ( .A(n_584), .B(n_532), .C(n_549), .D(n_554), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_607), .Y(n_627) );
AO22x1_ASAP7_75t_L g628 ( .A1(n_564), .A2(n_554), .B1(n_540), .B2(n_551), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_586), .B(n_540), .Y(n_629) );
AOI21xp33_ASAP7_75t_L g630 ( .A1(n_564), .A2(n_520), .B(n_559), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_572), .B(n_530), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_562), .A2(n_526), .B1(n_533), .B2(n_530), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_561), .B(n_533), .Y(n_633) );
O2A1O1Ixp5_ASAP7_75t_SL g634 ( .A1(n_613), .A2(n_556), .B(n_543), .C(n_559), .Y(n_634) );
OAI31xp33_ASAP7_75t_L g635 ( .A1(n_568), .A2(n_517), .A3(n_557), .B(n_520), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g636 ( .A1(n_568), .A2(n_560), .B1(n_556), .B2(n_518), .C(n_527), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_602), .A2(n_560), .B1(n_515), .B2(n_518), .C(n_527), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_577), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_608), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_577), .Y(n_640) );
NAND2x1_ASAP7_75t_SL g641 ( .A(n_613), .B(n_557), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_586), .B(n_505), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_561), .B(n_515), .Y(n_643) );
NOR4xp25_ASAP7_75t_SL g644 ( .A(n_595), .B(n_528), .C(n_542), .D(n_601), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_571), .A2(n_528), .B1(n_542), .B2(n_582), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_562), .A2(n_584), .B1(n_565), .B2(n_579), .Y(n_646) );
AOI222xp33_ASAP7_75t_L g647 ( .A1(n_567), .A2(n_612), .B1(n_606), .B2(n_574), .C1(n_578), .C2(n_576), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_567), .Y(n_648) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_608), .Y(n_649) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_579), .Y(n_650) );
XNOR2x2_ASAP7_75t_SL g651 ( .A(n_646), .B(n_606), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_649), .B(n_612), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_628), .A2(n_589), .B(n_571), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_649), .B(n_647), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_614), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_617), .B(n_576), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_650), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_650), .Y(n_658) );
INVxp67_ASAP7_75t_SL g659 ( .A(n_619), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_629), .B(n_613), .Y(n_660) );
NOR3x1_ASAP7_75t_L g661 ( .A(n_626), .B(n_589), .C(n_575), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_639), .B(n_578), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_617), .B(n_601), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_619), .A2(n_570), .B1(n_565), .B2(n_596), .C(n_599), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_616), .B(n_565), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_621), .B(n_596), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_648), .B(n_599), .Y(n_667) );
NAND2xp33_ASAP7_75t_L g668 ( .A(n_624), .B(n_583), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_622), .A2(n_588), .B1(n_594), .B2(n_593), .C(n_604), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_624), .A2(n_571), .B1(n_569), .B2(n_580), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_627), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_638), .Y(n_672) );
INVx1_ASAP7_75t_SL g673 ( .A(n_615), .Y(n_673) );
NAND2xp33_ASAP7_75t_SL g674 ( .A(n_654), .B(n_641), .Y(n_674) );
AOI32xp33_ASAP7_75t_L g675 ( .A1(n_659), .A2(n_623), .A3(n_645), .B1(n_618), .B2(n_642), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_664), .B(n_632), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_672), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_652), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_669), .A2(n_620), .B1(n_625), .B2(n_642), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_657), .B(n_631), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_665), .A2(n_636), .B1(n_643), .B2(n_633), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_671), .Y(n_682) );
AOI22x1_ASAP7_75t_L g683 ( .A1(n_653), .A2(n_605), .B1(n_603), .B2(n_644), .Y(n_683) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_658), .Y(n_684) );
AO22x1_ASAP7_75t_L g685 ( .A1(n_661), .A2(n_635), .B1(n_571), .B2(n_640), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g686 ( .A(n_656), .Y(n_686) );
XNOR2xp5_ASAP7_75t_L g687 ( .A(n_651), .B(n_637), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_682), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_685), .A2(n_670), .B(n_668), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_675), .A2(n_663), .B1(n_655), .B2(n_665), .C(n_658), .Y(n_690) );
OAI211xp5_ASAP7_75t_SL g691 ( .A1(n_676), .A2(n_668), .B(n_597), .C(n_666), .Y(n_691) );
NOR2x1_ASAP7_75t_L g692 ( .A(n_687), .B(n_673), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_674), .A2(n_667), .B1(n_630), .B2(n_662), .C(n_660), .Y(n_693) );
NAND4xp25_ASAP7_75t_SL g694 ( .A(n_679), .B(n_634), .C(n_662), .D(n_590), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_678), .A2(n_588), .B1(n_593), .B2(n_594), .C(n_603), .Y(n_695) );
INVxp67_ASAP7_75t_L g696 ( .A(n_692), .Y(n_696) );
NAND3xp33_ASAP7_75t_SL g697 ( .A(n_690), .B(n_686), .C(n_683), .Y(n_697) );
NOR2x1_ASAP7_75t_L g698 ( .A(n_689), .B(n_677), .Y(n_698) );
OAI211xp5_ASAP7_75t_L g699 ( .A1(n_693), .A2(n_681), .B(n_684), .C(n_680), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_696), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_698), .B(n_688), .Y(n_701) );
XNOR2xp5_ASAP7_75t_L g702 ( .A(n_697), .B(n_695), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_700), .Y(n_703) );
OA22x2_ASAP7_75t_L g704 ( .A1(n_702), .A2(n_699), .B1(n_694), .B2(n_684), .Y(n_704) );
OAI22xp5_ASAP7_75t_SL g705 ( .A1(n_703), .A2(n_701), .B1(n_691), .B2(n_569), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_705), .A2(n_704), .B(n_585), .Y(n_706) );
AOI222xp33_ASAP7_75t_SL g707 ( .A1(n_706), .A2(n_569), .B1(n_580), .B2(n_587), .C1(n_600), .C2(n_605), .Y(n_707) );
OA22x2_ASAP7_75t_L g708 ( .A1(n_707), .A2(n_591), .B1(n_592), .B2(n_587), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_708), .A2(n_598), .B1(n_600), .B2(n_697), .Y(n_709) );
endmodule