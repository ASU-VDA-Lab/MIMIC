module fake_jpeg_13480_n_517 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g148 ( 
.A(n_55),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_57),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_58),
.B(n_68),
.Y(n_140)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

CKINVDCx12_ASAP7_75t_R g125 ( 
.A(n_63),
.Y(n_125)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_0),
.C(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_67),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_33),
.B(n_1),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_1),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_75),
.Y(n_104)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_74),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_17),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_17),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_83),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_38),
.B(n_2),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_85),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_17),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_18),
.B(n_3),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_86),
.B(n_48),
.Y(n_155)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_91),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_18),
.B(n_14),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_3),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_17),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_100),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_38),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_105),
.B(n_112),
.Y(n_159)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_65),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_109),
.A2(n_30),
.B1(n_50),
.B2(n_46),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_23),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_80),
.B(n_21),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_23),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_124),
.B(n_155),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_74),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_82),
.B(n_32),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_151),
.Y(n_177)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_56),
.Y(n_142)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_142),
.Y(n_201)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_53),
.Y(n_144)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_88),
.B(n_40),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_60),
.B(n_35),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_158),
.Y(n_180)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_63),
.B(n_21),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_156),
.B(n_88),
.Y(n_185)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_64),
.Y(n_157)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_60),
.B(n_35),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_114),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_160),
.B(n_164),
.Y(n_223)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_103),
.A2(n_37),
.B1(n_93),
.B2(n_90),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_165),
.Y(n_220)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_166),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_135),
.A2(n_92),
.B1(n_69),
.B2(n_76),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_167),
.A2(n_170),
.B1(n_197),
.B2(n_205),
.Y(n_243)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_135),
.A2(n_92),
.B1(n_69),
.B2(n_76),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_173),
.A2(n_46),
.B1(n_50),
.B2(n_111),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_175),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_110),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_199),
.Y(n_211)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_42),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_181),
.B(n_182),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_115),
.B(n_42),
.Y(n_182)
);

CKINVDCx12_ASAP7_75t_R g183 ( 
.A(n_148),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_183),
.Y(n_219)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_185),
.B(n_186),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_113),
.B(n_55),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_115),
.B(n_66),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_150),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_106),
.B(n_43),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_192),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_151),
.A2(n_62),
.B1(n_30),
.B2(n_87),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_202),
.C(n_139),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_119),
.B(n_43),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_143),
.B(n_104),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_194),
.B(n_206),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_133),
.A2(n_44),
.B1(n_34),
.B2(n_54),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_141),
.B(n_44),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_120),
.B(n_34),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_200),
.B(n_204),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_127),
.B(n_55),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_133),
.A2(n_37),
.B1(n_97),
.B2(n_79),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g244 ( 
.A1(n_203),
.A2(n_126),
.B1(n_149),
.B2(n_111),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_145),
.B(n_142),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_145),
.A2(n_25),
.B1(n_47),
.B2(n_49),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_129),
.B(n_47),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_210),
.A2(n_108),
.B1(n_101),
.B2(n_121),
.Y(n_261)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_214),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_215),
.B(n_218),
.Y(n_285)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_204),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_225),
.B(n_231),
.Y(n_281)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_230),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_190),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_232),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_202),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_234),
.A2(n_179),
.B(n_196),
.Y(n_280)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_169),
.Y(n_238)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_180),
.B(n_174),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_181),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_134),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_241),
.B(n_211),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_244),
.A2(n_150),
.B1(n_201),
.B2(n_137),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_189),
.B(n_148),
.C(n_149),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_182),
.Y(n_258)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_198),
.Y(n_246)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_248),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_200),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_249),
.B(n_265),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_257),
.Y(n_292)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_217),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_251),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_247),
.A2(n_173),
.B1(n_177),
.B2(n_191),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_253),
.A2(n_262),
.B1(n_285),
.B2(n_268),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_254),
.B(n_264),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_242),
.B(n_171),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_258),
.B(n_285),
.C(n_262),
.Y(n_305)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_217),
.Y(n_260)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_261),
.A2(n_273),
.B1(n_278),
.B2(n_178),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_223),
.A2(n_218),
.B1(n_245),
.B2(n_243),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_199),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_159),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_161),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_268),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_213),
.B(n_208),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_267),
.B(n_269),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_165),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_165),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_270),
.B(n_272),
.Y(n_316)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_212),
.Y(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_172),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_210),
.A2(n_201),
.B1(n_131),
.B2(n_121),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_226),
.B(n_168),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_276),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_227),
.B(n_168),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_229),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_277),
.B(n_279),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_215),
.B(n_29),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_280),
.B(n_179),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_220),
.A2(n_216),
.B1(n_222),
.B2(n_238),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_282),
.A2(n_263),
.B1(n_255),
.B2(n_224),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_220),
.A2(n_134),
.B(n_138),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_283),
.A2(n_240),
.B(n_102),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_274),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_287),
.B(n_294),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_236),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_290),
.B(n_295),
.C(n_305),
.Y(n_322)
);

XNOR2x2_ASAP7_75t_L g291 ( 
.A(n_249),
.B(n_209),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_291),
.A2(n_264),
.B(n_254),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_276),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_228),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_296),
.A2(n_310),
.B1(n_311),
.B2(n_317),
.Y(n_333)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_297),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_267),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_299),
.B(n_312),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_SL g332 ( 
.A1(n_300),
.A2(n_301),
.B(n_102),
.C(n_138),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_283),
.A2(n_240),
.B(n_219),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_252),
.Y(n_302)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_302),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_281),
.A2(n_244),
.B1(n_248),
.B2(n_246),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_303),
.A2(n_304),
.B1(n_319),
.B2(n_284),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_266),
.A2(n_244),
.B1(n_126),
.B2(n_131),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_269),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_306),
.B(n_29),
.Y(n_353)
);

OAI32xp33_ASAP7_75t_L g308 ( 
.A1(n_272),
.A2(n_232),
.A3(n_230),
.B1(n_214),
.B2(n_222),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_280),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_253),
.A2(n_250),
.B1(n_277),
.B2(n_265),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_275),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_252),
.Y(n_313)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_313),
.Y(n_342)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_315),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_279),
.A2(n_244),
.B1(n_216),
.B2(n_237),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_318),
.B(n_74),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_321),
.B(n_323),
.Y(n_370)
);

AND2x6_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_296),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_301),
.A2(n_263),
.B(n_256),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_324),
.A2(n_332),
.B(n_107),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_325),
.B(n_52),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_329),
.B(n_338),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_304),
.A2(n_257),
.B1(n_251),
.B2(n_260),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_330),
.A2(n_336),
.B1(n_344),
.B2(n_346),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_306),
.A2(n_256),
.B1(n_255),
.B2(n_284),
.Y(n_331)
);

OAI21xp33_ASAP7_75t_L g373 ( 
.A1(n_331),
.A2(n_136),
.B(n_49),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_314),
.Y(n_334)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_334),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_259),
.Y(n_335)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_335),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_303),
.A2(n_251),
.B1(n_260),
.B2(n_273),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_294),
.Y(n_337)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_337),
.Y(n_382)
);

AO22x2_ASAP7_75t_L g338 ( 
.A1(n_287),
.A2(n_291),
.B1(n_317),
.B2(n_308),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_290),
.B(n_295),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_343),
.C(n_316),
.Y(n_360)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_289),
.Y(n_340)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_320),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_341),
.B(n_352),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_311),
.B(n_259),
.C(n_196),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_289),
.A2(n_255),
.B1(n_261),
.B2(n_237),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_297),
.A2(n_221),
.B1(n_184),
.B2(n_162),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_302),
.A2(n_221),
.B1(n_207),
.B2(n_50),
.Y(n_347)
);

OA22x2_ASAP7_75t_L g387 ( 
.A1(n_347),
.A2(n_336),
.B1(n_344),
.B2(n_346),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_293),
.B(n_207),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_353),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_349),
.B(n_117),
.Y(n_378)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_313),
.Y(n_350)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_350),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_292),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_293),
.B(n_48),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_354),
.B(n_3),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_325),
.B(n_288),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_369),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_333),
.A2(n_300),
.B1(n_298),
.B2(n_286),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_356),
.A2(n_365),
.B(n_385),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_292),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_357),
.B(n_362),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_324),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_375),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_321),
.A2(n_286),
.B1(n_307),
.B2(n_315),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_359),
.A2(n_329),
.B1(n_330),
.B2(n_348),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_360),
.B(n_374),
.C(n_361),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_322),
.B(n_318),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_361),
.B(n_363),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_334),
.B(n_307),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_322),
.B(n_166),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_195),
.Y(n_364)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_364),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_343),
.B(n_195),
.Y(n_366)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_351),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_373),
.A2(n_41),
.B1(n_50),
.B2(n_17),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_136),
.C(n_117),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_331),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_376),
.B(n_381),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_335),
.B(n_136),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_378),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_337),
.Y(n_381)
);

FAx1_ASAP7_75t_SL g384 ( 
.A(n_323),
.B(n_57),
.CI(n_107),
.CON(n_384),
.SN(n_384)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_387),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_390),
.A2(n_379),
.B1(n_387),
.B2(n_384),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_385),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_393),
.B(n_394),
.Y(n_421)
);

NOR3xp33_ASAP7_75t_SL g394 ( 
.A(n_386),
.B(n_332),
.C(n_327),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_396),
.B(n_406),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_356),
.A2(n_338),
.B1(n_332),
.B2(n_340),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_397),
.A2(n_379),
.B1(n_387),
.B2(n_384),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_360),
.B(n_349),
.C(n_328),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_398),
.B(n_403),
.C(n_404),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_358),
.A2(n_338),
.B(n_332),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_400),
.B(n_405),
.Y(n_431)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_367),
.Y(n_402)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_402),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_342),
.C(n_345),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_338),
.C(n_347),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_375),
.A2(n_4),
.B(n_5),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_368),
.B(n_378),
.Y(n_406)
);

INVxp33_ASAP7_75t_L g420 ( 
.A(n_407),
.Y(n_420)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_367),
.Y(n_410)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_410),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_380),
.B(n_382),
.Y(n_411)
);

CKINVDCx14_ASAP7_75t_R g438 ( 
.A(n_411),
.Y(n_438)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_383),
.Y(n_413)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_413),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_377),
.B(n_370),
.C(n_359),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_414),
.B(n_370),
.C(n_372),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_371),
.B(n_25),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_415),
.B(n_39),
.Y(n_430)
);

OA21x2_ASAP7_75t_L g416 ( 
.A1(n_371),
.A2(n_4),
.B(n_5),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_416),
.B(n_11),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_390),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_422),
.A2(n_425),
.B1(n_400),
.B2(n_393),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_396),
.B(n_365),
.C(n_372),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_424),
.B(n_432),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_389),
.B(n_376),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_430),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_401),
.A2(n_387),
.B1(n_41),
.B2(n_25),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_429),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_391),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_389),
.B(n_39),
.C(n_24),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_433),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_39),
.C(n_8),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_436),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_403),
.B(n_7),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_435),
.B(n_437),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_11),
.C(n_12),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_404),
.B(n_392),
.C(n_406),
.Y(n_437)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_439),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_440),
.B(n_457),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_431),
.B(n_399),
.Y(n_441)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_441),
.Y(n_460)
);

INVx13_ASAP7_75t_L g445 ( 
.A(n_438),
.Y(n_445)
);

INVx11_ASAP7_75t_L g473 ( 
.A(n_445),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_392),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_448),
.B(n_427),
.Y(n_467)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_417),
.Y(n_449)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_449),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_421),
.Y(n_452)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_452),
.Y(n_468)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_423),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_453),
.A2(n_441),
.B1(n_420),
.B2(n_446),
.Y(n_474)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_426),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_458),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_455),
.A2(n_397),
.B1(n_409),
.B2(n_388),
.Y(n_464)
);

INVx13_ASAP7_75t_L g456 ( 
.A(n_420),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_456),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_422),
.A2(n_409),
.B(n_399),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_424),
.B(n_412),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_418),
.C(n_428),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_465),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_464),
.B(n_470),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_418),
.C(n_419),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_443),
.A2(n_411),
.B1(n_408),
.B2(n_395),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_472),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_467),
.B(n_447),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_388),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_446),
.Y(n_471)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_471),
.Y(n_486)
);

BUFx24_ASAP7_75t_SL g472 ( 
.A(n_442),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_474),
.B(n_475),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_447),
.B(n_434),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_441),
.C(n_457),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_482),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_450),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_463),
.A2(n_451),
.B(n_444),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_478),
.A2(n_480),
.B(n_484),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_469),
.Y(n_479)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_479),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_465),
.A2(n_468),
.B(n_473),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_415),
.C(n_443),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_460),
.A2(n_473),
.B(n_464),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_459),
.A2(n_445),
.B(n_394),
.Y(n_488)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_488),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_461),
.B(n_436),
.C(n_456),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_489),
.B(n_14),
.C(n_11),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_485),
.B(n_433),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_490),
.B(n_491),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_482),
.B(n_416),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_492),
.B(n_483),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_479),
.A2(n_453),
.B1(n_405),
.B2(n_416),
.Y(n_494)
);

CKINVDCx14_ASAP7_75t_R g503 ( 
.A(n_494),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_481),
.A2(n_407),
.B(n_12),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_495),
.A2(n_498),
.B(n_489),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_500),
.B(n_506),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_502),
.B(n_505),
.Y(n_509)
);

NOR2xp67_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_476),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_504),
.A2(n_493),
.B(n_499),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_496),
.A2(n_488),
.B(n_486),
.Y(n_505)
);

BUFx24_ASAP7_75t_SL g506 ( 
.A(n_496),
.Y(n_506)
);

AOI21x1_ASAP7_75t_L g511 ( 
.A1(n_508),
.A2(n_501),
.B(n_498),
.Y(n_511)
);

AOI211xp5_ASAP7_75t_L g510 ( 
.A1(n_503),
.A2(n_497),
.B(n_487),
.C(n_491),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_510),
.B(n_487),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_511),
.A2(n_512),
.B(n_509),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_513),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_514),
.A2(n_507),
.B(n_490),
.Y(n_515)
);

O2A1O1Ixp33_ASAP7_75t_SL g516 ( 
.A1(n_515),
.A2(n_13),
.B(n_512),
.C(n_481),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_516),
.Y(n_517)
);


endmodule