module real_aes_3176_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_287;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_987;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_979;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_974;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_884;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_983;
wire n_767;
wire n_138;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_961;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_981;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_976;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_984;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_962;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_164;
wire n_671;
wire n_973;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_617;
wire n_402;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_972;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_928;
wire n_243;
wire n_899;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_926;
wire n_922;
wire n_149;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_134;
wire n_946;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_982;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_968;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx1_ASAP7_75t_L g672 ( .A(n_0), .Y(n_672) );
INVx1_ASAP7_75t_L g168 ( .A(n_1), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_2), .A2(n_17), .B1(n_215), .B2(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g320 ( .A(n_3), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_4), .B(n_591), .Y(n_636) );
INVx1_ASAP7_75t_SL g184 ( .A(n_5), .Y(n_184) );
INVxp67_ASAP7_75t_L g121 ( .A(n_6), .Y(n_121) );
BUFx2_ASAP7_75t_L g574 ( .A(n_6), .Y(n_574) );
INVx1_ASAP7_75t_L g979 ( .A(n_6), .Y(n_979) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_7), .B(n_204), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_8), .A2(n_40), .B1(n_590), .B2(n_595), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_9), .A2(n_46), .B1(n_271), .B2(n_618), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_10), .A2(n_69), .B1(n_621), .B2(n_680), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_11), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_12), .B(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g667 ( .A(n_13), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_14), .A2(n_56), .B1(n_203), .B2(n_204), .Y(n_202) );
INVx1_ASAP7_75t_L g670 ( .A(n_15), .Y(n_670) );
OA21x2_ASAP7_75t_L g147 ( .A1(n_16), .A2(n_73), .B(n_148), .Y(n_147) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_16), .A2(n_73), .B(n_148), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_18), .A2(n_71), .B1(n_621), .B2(n_680), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_19), .B(n_170), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_20), .A2(n_85), .B1(n_315), .B2(n_316), .Y(n_314) );
INVx2_ASAP7_75t_L g276 ( .A(n_21), .Y(n_276) );
INVx1_ASAP7_75t_L g664 ( .A(n_22), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_23), .A2(n_27), .B1(n_183), .B2(n_240), .Y(n_253) );
BUFx3_ASAP7_75t_L g113 ( .A(n_24), .Y(n_113) );
O2A1O1Ixp5_ASAP7_75t_L g270 ( .A1(n_25), .A2(n_158), .B(n_271), .C(n_273), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_26), .A2(n_66), .B1(n_272), .B2(n_292), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_28), .Y(n_241) );
AO22x1_ASAP7_75t_L g633 ( .A1(n_29), .A2(n_83), .B1(n_192), .B2(n_634), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_30), .Y(n_604) );
AND2x2_ASAP7_75t_L g695 ( .A(n_31), .B(n_618), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_32), .B(n_192), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_33), .A2(n_86), .B1(n_211), .B2(n_214), .Y(n_210) );
INVx1_ASAP7_75t_L g126 ( .A(n_34), .Y(n_126) );
INVx1_ASAP7_75t_L g266 ( .A(n_35), .Y(n_266) );
AOI22x1_ASAP7_75t_L g620 ( .A1(n_36), .A2(n_102), .B1(n_588), .B2(n_621), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_37), .A2(n_565), .B1(n_566), .B2(n_570), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_37), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_38), .B(n_559), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_39), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_39), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g986 ( .A(n_41), .B(n_987), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_42), .B(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g274 ( .A(n_43), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_44), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_45), .B(n_647), .Y(n_702) );
INVx2_ASAP7_75t_L g293 ( .A(n_47), .Y(n_293) );
NAND3xp33_ASAP7_75t_SL g137 ( .A(n_48), .B(n_138), .C(n_395), .Y(n_137) );
INVx1_ASAP7_75t_L g544 ( .A(n_48), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_49), .B(n_156), .Y(n_155) );
INVx1_ASAP7_75t_SL g191 ( .A(n_50), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_51), .B(n_183), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g974 ( .A(n_52), .Y(n_974) );
INVx1_ASAP7_75t_L g235 ( .A(n_53), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_54), .B(n_268), .Y(n_607) );
INVx1_ASAP7_75t_L g148 ( .A(n_55), .Y(n_148) );
AND2x4_ASAP7_75t_L g174 ( .A(n_57), .B(n_175), .Y(n_174) );
AND2x4_ASAP7_75t_L g230 ( .A(n_57), .B(n_175), .Y(n_230) );
XNOR2xp5_ASAP7_75t_L g566 ( .A(n_58), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g197 ( .A(n_59), .Y(n_197) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_60), .Y(n_159) );
INVx2_ASAP7_75t_L g682 ( .A(n_61), .Y(n_682) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_62), .A2(n_128), .B1(n_129), .B2(n_130), .Y(n_127) );
INVx1_ASAP7_75t_L g129 ( .A(n_62), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_63), .A2(n_79), .B1(n_588), .B2(n_590), .Y(n_587) );
CKINVDCx14_ASAP7_75t_R g640 ( .A(n_64), .Y(n_640) );
AND2x2_ASAP7_75t_L g700 ( .A(n_65), .B(n_192), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_67), .B(n_186), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_68), .B(n_156), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_70), .B(n_145), .Y(n_643) );
NAND2x1p5_ASAP7_75t_L g703 ( .A(n_72), .B(n_613), .Y(n_703) );
CKINVDCx14_ASAP7_75t_R g624 ( .A(n_74), .Y(n_624) );
AOI22x1_ASAP7_75t_SL g567 ( .A1(n_75), .A2(n_97), .B1(n_568), .B2(n_569), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_75), .Y(n_568) );
OAI22x1_ASAP7_75t_SL g550 ( .A1(n_76), .A2(n_89), .B1(n_551), .B2(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g552 ( .A(n_76), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_77), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_78), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_80), .B(n_591), .Y(n_648) );
OR2x6_ASAP7_75t_L g123 ( .A(n_81), .B(n_124), .Y(n_123) );
AND3x1_ASAP7_75t_L g985 ( .A(n_81), .B(n_574), .C(n_986), .Y(n_985) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_82), .B(n_153), .Y(n_193) );
INVx1_ASAP7_75t_L g125 ( .A(n_84), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_84), .B(n_126), .Y(n_984) );
INVx1_ASAP7_75t_L g987 ( .A(n_87), .Y(n_987) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_88), .Y(n_154) );
BUFx5_ASAP7_75t_L g157 ( .A(n_88), .Y(n_157) );
INVx1_ASAP7_75t_L g188 ( .A(n_88), .Y(n_188) );
INVx1_ASAP7_75t_L g551 ( .A(n_89), .Y(n_551) );
INVx2_ASAP7_75t_L g674 ( .A(n_90), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_91), .B(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g296 ( .A(n_92), .Y(n_296) );
AOI32xp33_ASAP7_75t_L g105 ( .A1(n_93), .A2(n_106), .A3(n_562), .B1(n_980), .B2(n_988), .Y(n_105) );
INVx1_ASAP7_75t_L g300 ( .A(n_94), .Y(n_300) );
NAND2xp33_ASAP7_75t_L g697 ( .A(n_95), .B(n_589), .Y(n_697) );
INVx2_ASAP7_75t_L g244 ( .A(n_96), .Y(n_244) );
INVx1_ASAP7_75t_L g569 ( .A(n_97), .Y(n_569) );
INVx2_ASAP7_75t_SL g175 ( .A(n_98), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_99), .B(n_233), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_100), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_101), .B(n_145), .Y(n_144) );
AO32x2_ASAP7_75t_L g249 ( .A1(n_103), .A2(n_220), .A3(n_250), .B1(n_255), .B2(n_256), .Y(n_249) );
AO22x2_ASAP7_75t_L g328 ( .A1(n_103), .A2(n_250), .B1(n_329), .B2(n_331), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_104), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_114), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g971 ( .A(n_109), .Y(n_971) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
BUFx8_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
CKINVDCx6p67_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI21x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_131), .B(n_554), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_127), .Y(n_116) );
INVx2_ASAP7_75t_L g556 ( .A(n_117), .Y(n_556) );
BUFx4f_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx12f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx8_ASAP7_75t_L g561 ( .A(n_119), .Y(n_561) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
INVx8_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_123), .A2(n_563), .B(n_970), .Y(n_562) );
OR2x6_ASAP7_75t_L g978 ( .A(n_123), .B(n_979), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_127), .B(n_556), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_128), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_SL g554 ( .A1(n_133), .A2(n_555), .B(n_557), .Y(n_554) );
OAI22x1_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_135), .B1(n_550), .B2(n_553), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_135), .A2(n_572), .B(n_575), .Y(n_571) );
OR2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_541), .Y(n_135) );
NOR2x1_ASAP7_75t_L g136 ( .A(n_137), .B(n_458), .Y(n_136) );
INVx1_ASAP7_75t_L g543 ( .A(n_138), .Y(n_543) );
NOR4xp75_ASAP7_75t_L g138 ( .A(n_139), .B(n_321), .C(n_358), .D(n_381), .Y(n_138) );
OAI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_245), .B(n_277), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OAI21xp33_ASAP7_75t_L g522 ( .A1(n_141), .A2(n_515), .B(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_198), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_176), .Y(n_142) );
INVx1_ASAP7_75t_L g305 ( .A(n_143), .Y(n_305) );
INVx2_ASAP7_75t_L g335 ( .A(n_143), .Y(n_335) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_143), .Y(n_340) );
INVx1_ASAP7_75t_L g402 ( .A(n_143), .Y(n_402) );
AND2x2_ASAP7_75t_L g442 ( .A(n_143), .B(n_200), .Y(n_442) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_149), .Y(n_143) );
NOR2x1_ASAP7_75t_L g653 ( .A(n_145), .B(n_654), .Y(n_653) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx3_ASAP7_75t_L g255 ( .A(n_146), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_146), .B(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_146), .B(n_320), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_146), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx4_ASAP7_75t_L g180 ( .A(n_147), .Y(n_180) );
BUFx3_ASAP7_75t_L g285 ( .A(n_147), .Y(n_285) );
OAI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_160), .B(n_171), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_155), .B(n_158), .Y(n_150) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g183 ( .A(n_153), .Y(n_183) );
INVx1_ASAP7_75t_L g204 ( .A(n_153), .Y(n_204) );
INVx2_ASAP7_75t_L g316 ( .A(n_153), .Y(n_316) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx6_ASAP7_75t_L g170 ( .A(n_154), .Y(n_170) );
INVx2_ASAP7_75t_L g213 ( .A(n_154), .Y(n_213) );
INVx2_ASAP7_75t_L g215 ( .A(n_154), .Y(n_215) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g165 ( .A(n_157), .Y(n_165) );
INVx2_ASAP7_75t_L g192 ( .A(n_157), .Y(n_192) );
INVx2_ASAP7_75t_L g203 ( .A(n_157), .Y(n_203) );
INVx2_ASAP7_75t_L g240 ( .A(n_157), .Y(n_240) );
INVx2_ASAP7_75t_L g591 ( .A(n_157), .Y(n_591) );
INVx4_ASAP7_75t_L g238 ( .A(n_158), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_158), .A2(n_251), .B1(n_253), .B2(n_254), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_158), .B(n_586), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_158), .A2(n_590), .B1(n_602), .B2(n_605), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_158), .A2(n_646), .B(n_648), .Y(n_645) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx4_ASAP7_75t_L g163 ( .A(n_159), .Y(n_163) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_159), .Y(n_189) );
INVx3_ASAP7_75t_L g194 ( .A(n_159), .Y(n_194) );
INVx1_ASAP7_75t_L g217 ( .A(n_159), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_159), .B(n_664), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_159), .B(n_667), .Y(n_666) );
INVxp67_ASAP7_75t_L g698 ( .A(n_159), .Y(n_698) );
OAI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_164), .B(n_166), .Y(n_160) );
AND2x2_ASAP7_75t_L g263 ( .A(n_162), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g265 ( .A(n_162), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_163), .B(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_SL g669 ( .A(n_163), .B(n_670), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_163), .B(n_672), .Y(n_671) );
NAND3xp33_ASAP7_75t_SL g677 ( .A(n_163), .B(n_660), .C(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_169), .Y(n_166) );
OAI22xp33_ASAP7_75t_L g239 ( .A1(n_169), .A2(n_240), .B1(n_241), .B2(n_242), .Y(n_239) );
INVx2_ASAP7_75t_L g618 ( .A(n_169), .Y(n_618) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_SL g252 ( .A(n_170), .Y(n_252) );
INVx2_ASAP7_75t_L g262 ( .A(n_170), .Y(n_262) );
INVx1_ASAP7_75t_L g292 ( .A(n_170), .Y(n_292) );
INVx1_ASAP7_75t_L g589 ( .A(n_170), .Y(n_589) );
INVx1_ASAP7_75t_L g647 ( .A(n_170), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
INVx1_ASAP7_75t_L g196 ( .A(n_172), .Y(n_196) );
NOR2xp67_ASAP7_75t_L g206 ( .A(n_172), .B(n_173), .Y(n_206) );
BUFx3_ASAP7_75t_L g208 ( .A(n_172), .Y(n_208) );
INVx1_ASAP7_75t_L g221 ( .A(n_172), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_172), .B(n_173), .Y(n_298) );
INVx1_ASAP7_75t_L g330 ( .A(n_172), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_172), .B(n_173), .Y(n_586) );
INVx2_ASAP7_75t_L g660 ( .A(n_172), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_173), .B(n_179), .Y(n_178) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_174), .Y(n_256) );
AND2x2_ASAP7_75t_L g311 ( .A(n_174), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g329 ( .A(n_174), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g631 ( .A(n_174), .Y(n_631) );
INVx3_ASAP7_75t_L g654 ( .A(n_174), .Y(n_654) );
INVx1_ASAP7_75t_L g380 ( .A(n_176), .Y(n_380) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
OR2x2_ASAP7_75t_L g282 ( .A(n_177), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g306 ( .A(n_177), .Y(n_306) );
AND2x2_ASAP7_75t_L g336 ( .A(n_177), .B(n_218), .Y(n_336) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_177), .Y(n_389) );
INVx2_ASAP7_75t_L g405 ( .A(n_177), .Y(n_405) );
INVx1_ASAP7_75t_L g411 ( .A(n_177), .Y(n_411) );
AO31x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_181), .A3(n_190), .B(n_195), .Y(n_177) );
INVx2_ASAP7_75t_L g312 ( .A(n_179), .Y(n_312) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx3_ASAP7_75t_L g613 ( .A(n_180), .Y(n_613) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_184), .B(n_185), .C(n_189), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g272 ( .A(n_187), .Y(n_272) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g227 ( .A(n_188), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_189), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g254 ( .A(n_189), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g295 ( .A1(n_189), .A2(n_226), .B(n_296), .C(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g317 ( .A(n_189), .Y(n_317) );
INVxp67_ASAP7_75t_L g609 ( .A(n_189), .Y(n_609) );
INVx2_ASAP7_75t_SL g638 ( .A(n_189), .Y(n_638) );
INVx1_ASAP7_75t_L g652 ( .A(n_189), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_193), .C(n_194), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_192), .A2(n_268), .B1(n_669), .B2(n_671), .Y(n_668) );
INVx3_ASAP7_75t_L g231 ( .A(n_194), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_194), .A2(n_291), .B(n_293), .C(n_294), .Y(n_290) );
NOR2xp33_ASAP7_75t_SL g195 ( .A(n_196), .B(n_197), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_196), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g597 ( .A(n_196), .Y(n_597) );
AND2x2_ASAP7_75t_L g421 ( .A(n_198), .B(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g478 ( .A(n_198), .B(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_218), .Y(n_198) );
AND2x2_ASAP7_75t_L g341 ( .A(n_199), .B(n_342), .Y(n_341) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_199), .Y(n_351) );
BUFx2_ASAP7_75t_L g367 ( .A(n_199), .Y(n_367) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g281 ( .A(n_200), .Y(n_281) );
AND2x2_ASAP7_75t_L g334 ( .A(n_200), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g430 ( .A(n_200), .Y(n_430) );
NAND2x1p5_ASAP7_75t_L g200 ( .A(n_201), .B(n_209), .Y(n_200) );
AND2x2_ASAP7_75t_SL g304 ( .A(n_201), .B(n_209), .Y(n_304) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_205), .B(n_207), .Y(n_201) );
INVx2_ASAP7_75t_L g621 ( .A(n_203), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_206), .B(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_216), .Y(n_209) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g233 ( .A(n_213), .Y(n_233) );
INVxp67_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g268 ( .A(n_215), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_217), .B(n_586), .Y(n_593) );
INVx1_ASAP7_75t_L g619 ( .A(n_217), .Y(n_619) );
OR2x2_ASAP7_75t_L g353 ( .A(n_218), .B(n_335), .Y(n_353) );
AND2x2_ASAP7_75t_L g463 ( .A(n_218), .B(n_464), .Y(n_463) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_222), .B(n_243), .Y(n_218) );
INVxp67_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_221), .B(n_244), .Y(n_243) );
AO21x2_ASAP7_75t_L g283 ( .A1(n_222), .A2(n_243), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_236), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_228), .B1(n_232), .B2(n_234), .Y(n_223) );
NOR2xp67_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g315 ( .A(n_227), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_231), .Y(n_228) );
NOR3xp33_ASAP7_75t_L g234 ( .A(n_229), .B(n_231), .C(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_229), .B(n_238), .Y(n_237) );
AOI221x1_ASAP7_75t_L g259 ( .A1(n_229), .A2(n_260), .B1(n_263), .B2(n_265), .C(n_267), .Y(n_259) );
INVx4_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_231), .A2(n_314), .B1(n_317), .B2(n_318), .Y(n_313) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_231), .B(n_660), .C(n_678), .Y(n_684) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_239), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_238), .B(n_603), .Y(n_602) );
OAI22x1_ASAP7_75t_L g616 ( .A1(n_238), .A2(n_617), .B1(n_619), .B2(n_620), .Y(n_616) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVxp67_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g324 ( .A(n_247), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_257), .Y(n_247) );
AND2x2_ASAP7_75t_L g373 ( .A(n_248), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_248), .B(n_417), .Y(n_416) );
AND2x4_ASAP7_75t_L g486 ( .A(n_248), .B(n_288), .Y(n_486) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
BUFx8_ASAP7_75t_L g301 ( .A(n_249), .Y(n_301) );
AND2x2_ASAP7_75t_L g433 ( .A(n_249), .B(n_417), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_252), .B(n_274), .Y(n_273) );
AO31x2_ASAP7_75t_L g258 ( .A1(n_255), .A2(n_259), .A3(n_269), .B(n_275), .Y(n_258) );
INVx2_ASAP7_75t_L g331 ( .A(n_255), .Y(n_331) );
OAI21x1_ASAP7_75t_L g600 ( .A1(n_256), .A2(n_601), .B(n_606), .Y(n_600) );
AO31x2_ASAP7_75t_L g615 ( .A1(n_256), .A2(n_616), .A3(n_622), .B(n_623), .Y(n_615) );
AO31x2_ASAP7_75t_L g691 ( .A1(n_256), .A2(n_616), .A3(n_622), .B(n_623), .Y(n_691) );
AND2x2_ASAP7_75t_L g308 ( .A(n_257), .B(n_309), .Y(n_308) );
BUFx3_ASAP7_75t_L g355 ( .A(n_257), .Y(n_355) );
INVx2_ASAP7_75t_SL g374 ( .A(n_257), .Y(n_374) );
INVx1_ASAP7_75t_L g392 ( .A(n_257), .Y(n_392) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g287 ( .A(n_258), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_258), .B(n_326), .Y(n_346) );
OR2x2_ASAP7_75t_L g363 ( .A(n_258), .B(n_326), .Y(n_363) );
AND2x2_ASAP7_75t_L g407 ( .A(n_258), .B(n_357), .Y(n_407) );
INVx1_ASAP7_75t_L g425 ( .A(n_258), .Y(n_425) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_268), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_286), .B1(n_302), .B2(n_307), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_278), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
AND2x2_ASAP7_75t_L g388 ( .A(n_280), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g435 ( .A(n_280), .Y(n_435) );
AND2x2_ASAP7_75t_L g507 ( .A(n_280), .B(n_336), .Y(n_507) );
AND2x4_ASAP7_75t_L g518 ( .A(n_280), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g527 ( .A(n_282), .Y(n_527) );
INVx2_ASAP7_75t_L g342 ( .A(n_283), .Y(n_342) );
BUFx2_ASAP7_75t_L g394 ( .A(n_283), .Y(n_394) );
AND2x2_ASAP7_75t_L g404 ( .A(n_283), .B(n_405), .Y(n_404) );
NOR2xp67_ASAP7_75t_SL g623 ( .A(n_284), .B(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g639 ( .A(n_284), .B(n_640), .Y(n_639) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OA21x2_ASAP7_75t_L g599 ( .A1(n_285), .A2(n_600), .B(n_610), .Y(n_599) );
OA21x2_ASAP7_75t_L g725 ( .A1(n_285), .A2(n_600), .B(n_610), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_286), .B(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g506 ( .A(n_286), .B(n_480), .Y(n_506) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_301), .Y(n_286) );
INVx2_ASAP7_75t_L g415 ( .A(n_287), .Y(n_415) );
NAND2x1p5_ASAP7_75t_L g470 ( .A(n_287), .B(n_370), .Y(n_470) );
AND2x2_ASAP7_75t_L g494 ( .A(n_287), .B(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g511 ( .A(n_287), .Y(n_511) );
BUFx3_ASAP7_75t_L g332 ( .A(n_288), .Y(n_332) );
INVx1_ASAP7_75t_L g348 ( .A(n_288), .Y(n_348) );
INVx2_ASAP7_75t_L g357 ( .A(n_288), .Y(n_357) );
AND2x4_ASAP7_75t_L g424 ( .A(n_288), .B(n_425), .Y(n_424) );
INVx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AO31x2_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_295), .A3(n_298), .B(n_299), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g307 ( .A(n_301), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g364 ( .A(n_301), .B(n_365), .Y(n_364) );
INVxp67_ASAP7_75t_SL g383 ( .A(n_301), .Y(n_383) );
AND2x2_ASAP7_75t_L g406 ( .A(n_301), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_SL g423 ( .A(n_301), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g452 ( .A(n_301), .Y(n_452) );
AND2x2_ASAP7_75t_L g467 ( .A(n_301), .B(n_374), .Y(n_467) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_303), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g378 ( .A(n_304), .Y(n_378) );
INVx2_ASAP7_75t_L g464 ( .A(n_304), .Y(n_464) );
AND2x2_ASAP7_75t_L g514 ( .A(n_304), .B(n_305), .Y(n_514) );
INVx1_ASAP7_75t_L g386 ( .A(n_305), .Y(n_386) );
AND2x2_ASAP7_75t_L g422 ( .A(n_306), .B(n_402), .Y(n_422) );
OAI31xp67_ASAP7_75t_L g322 ( .A1(n_307), .A2(n_323), .A3(n_327), .B(n_333), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_308), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g485 ( .A(n_308), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g481 ( .A(n_309), .Y(n_481) );
AND2x2_ASAP7_75t_L g502 ( .A(n_309), .B(n_357), .Y(n_502) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g326 ( .A(n_310), .Y(n_326) );
INVx1_ASAP7_75t_L g372 ( .A(n_310), .Y(n_372) );
AOI21x1_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_313), .B(n_319), .Y(n_310) );
AOI21xp33_ASAP7_75t_SL g705 ( .A1(n_312), .A2(n_678), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g634 ( .A(n_315), .Y(n_634) );
INVx1_ASAP7_75t_L g595 ( .A(n_316), .Y(n_595) );
INVx1_ASAP7_75t_L g680 ( .A(n_316), .Y(n_680) );
AOI21x1_ASAP7_75t_L g632 ( .A1(n_317), .A2(n_633), .B(n_635), .Y(n_632) );
NAND2x1_ASAP7_75t_L g321 ( .A(n_322), .B(n_337), .Y(n_321) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_324), .B(n_344), .Y(n_343) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g473 ( .A(n_327), .B(n_474), .Y(n_473) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_332), .Y(n_327) );
INVx1_ASAP7_75t_L g349 ( .A(n_328), .Y(n_349) );
AND2x4_ASAP7_75t_L g356 ( .A(n_328), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g495 ( .A(n_328), .Y(n_495) );
INVx2_ASAP7_75t_SL g391 ( .A(n_332), .Y(n_391) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
AND2x2_ASAP7_75t_L g408 ( .A(n_334), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g449 ( .A(n_334), .B(n_379), .Y(n_449) );
NAND2xp67_ASAP7_75t_L g526 ( .A(n_334), .B(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g538 ( .A(n_334), .Y(n_538) );
AND2x2_ASAP7_75t_L g366 ( .A(n_336), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g441 ( .A(n_336), .B(n_442), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_343), .B1(n_350), .B2(n_354), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
INVx1_ASAP7_75t_L g490 ( .A(n_339), .Y(n_490) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g479 ( .A(n_340), .B(n_410), .Y(n_479) );
AND2x4_ASAP7_75t_L g379 ( .A(n_342), .B(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g457 ( .A(n_342), .B(n_402), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g365 ( .A(n_346), .Y(n_365) );
AND2x2_ASAP7_75t_L g398 ( .A(n_347), .B(n_355), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_347), .B(n_440), .Y(n_487) );
AND2x2_ASAP7_75t_L g515 ( .A(n_347), .B(n_481), .Y(n_515) );
AND2x4_ASAP7_75t_SL g347 ( .A(n_348), .B(n_349), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_350), .B(n_501), .Y(n_500) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVxp67_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g431 ( .A(n_353), .Y(n_431) );
INVxp67_ASAP7_75t_L g519 ( .A(n_353), .Y(n_519) );
OR2x6_ASAP7_75t_L g529 ( .A(n_353), .B(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
AND2x2_ASAP7_75t_L g501 ( .A(n_355), .B(n_502), .Y(n_501) );
INVx4_ASAP7_75t_L g361 ( .A(n_356), .Y(n_361) );
AND2x2_ASAP7_75t_L g375 ( .A(n_356), .B(n_371), .Y(n_375) );
AND2x4_ASAP7_75t_L g439 ( .A(n_356), .B(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_SL g466 ( .A(n_356), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_368), .Y(n_358) );
OAI21xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_364), .B(n_366), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_362), .A2(n_428), .B1(n_432), .B2(n_434), .Y(n_427) );
AND2x2_ASAP7_75t_L g469 ( .A(n_362), .B(n_391), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_362), .B(n_390), .Y(n_533) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g440 ( .A(n_363), .Y(n_440) );
OR2x2_ASAP7_75t_L g451 ( .A(n_363), .B(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g517 ( .A(n_365), .B(n_495), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_375), .B(n_376), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_369), .A2(n_423), .B1(n_525), .B2(n_528), .Y(n_524) );
AND2x4_ASAP7_75t_L g369 ( .A(n_370), .B(n_373), .Y(n_369) );
AND2x2_ASAP7_75t_L g523 ( .A(n_370), .B(n_424), .Y(n_523) );
INVx4_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g446 ( .A(n_371), .B(n_407), .Y(n_446) );
AND2x2_ASAP7_75t_L g454 ( .A(n_371), .B(n_424), .Y(n_454) );
INVx2_ASAP7_75t_L g474 ( .A(n_371), .Y(n_474) );
BUFx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g417 ( .A(n_372), .Y(n_417) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_379), .B(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_L g476 ( .A(n_379), .B(n_401), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_379), .A2(n_492), .B(n_497), .Y(n_491) );
AND2x2_ASAP7_75t_L g513 ( .A(n_379), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g535 ( .A(n_379), .Y(n_535) );
OAI21xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B(n_387), .Y(n_381) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND5xp2_ASAP7_75t_L g387 ( .A(n_386), .B(n_388), .C(n_390), .D(n_392), .E(n_393), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_SL g445 ( .A(n_392), .B(n_433), .Y(n_445) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NOR3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_426), .C(n_443), .Y(n_395) );
INVxp67_ASAP7_75t_L g547 ( .A(n_396), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_412), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B1(n_406), .B2(n_408), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_400), .B(n_403), .Y(n_399) );
AND2x2_ASAP7_75t_L g447 ( .A(n_400), .B(n_404), .Y(n_447) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_403), .B(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_405), .Y(n_437) );
INVxp67_ASAP7_75t_SL g530 ( .A(n_405), .Y(n_530) );
OR2x2_ASAP7_75t_L g537 ( .A(n_405), .B(n_481), .Y(n_537) );
AND2x2_ASAP7_75t_L g432 ( .A(n_407), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g455 ( .A(n_407), .B(n_452), .Y(n_455) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_410), .Y(n_420) );
AND2x2_ASAP7_75t_L g429 ( .A(n_410), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_418), .B1(n_421), .B2(n_423), .Y(n_412) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
NOR2xp67_ASAP7_75t_L g536 ( .A(n_415), .B(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_421), .A2(n_455), .B1(n_517), .B2(n_518), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_421), .B(n_533), .Y(n_532) );
AND2x4_ASAP7_75t_L g462 ( .A(n_422), .B(n_463), .Y(n_462) );
INVxp67_ASAP7_75t_SL g549 ( .A(n_426), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_438), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_428), .A2(n_510), .B1(n_513), .B2(n_515), .Y(n_509) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
NOR2xp33_ASAP7_75t_SL g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NOR2xp67_ASAP7_75t_L g456 ( .A(n_437), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_439), .B(n_441), .Y(n_438) );
INVxp67_ASAP7_75t_L g548 ( .A(n_443), .Y(n_548) );
NAND3xp33_ASAP7_75t_SL g443 ( .A(n_444), .B(n_448), .C(n_453), .Y(n_443) );
OAI21xp5_ASAP7_75t_SL g444 ( .A1(n_445), .A2(n_446), .B(n_447), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_445), .A2(n_535), .B(n_536), .C(n_538), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_455), .B(n_456), .Y(n_453) );
NOR2xp67_ASAP7_75t_SL g499 ( .A(n_457), .B(n_464), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_503), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI21xp33_ASAP7_75t_L g545 ( .A1(n_460), .A2(n_544), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_491), .Y(n_460) );
AOI211xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_465), .B(n_471), .C(n_482), .Y(n_461) );
INVx2_ASAP7_75t_L g483 ( .A(n_462), .Y(n_483) );
NAND3xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .C(n_470), .Y(n_465) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx3_ASAP7_75t_L g540 ( .A(n_470), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_475), .B1(n_477), .B2(n_480), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g496 ( .A(n_480), .Y(n_496) );
BUFx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B1(n_487), .B2(n_488), .Y(n_482) );
INVx2_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_496), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_500), .Y(n_497) );
INVx1_ASAP7_75t_L g512 ( .A(n_502), .Y(n_512) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OAI21xp33_ASAP7_75t_L g542 ( .A1(n_504), .A2(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_520), .Y(n_504) );
AOI21xp5_ASAP7_75t_SL g505 ( .A1(n_506), .A2(n_507), .B(n_508), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_516), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_511), .B(n_512), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_531), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_524), .Y(n_521) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVxp67_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .C(n_539), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_545), .Y(n_541) );
NAND3xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .C(n_549), .Y(n_546) );
INVxp67_ASAP7_75t_R g553 ( .A(n_550), .Y(n_553) );
CKINVDCx14_ASAP7_75t_R g557 ( .A(n_558), .Y(n_557) );
NAND3xp33_ASAP7_75t_L g970 ( .A(n_558), .B(n_971), .C(n_972), .Y(n_970) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
XNOR2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_571), .Y(n_563) );
INVx1_ASAP7_75t_L g570 ( .A(n_566), .Y(n_570) );
NOR2x1_ASAP7_75t_L g575 ( .A(n_572), .B(n_576), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_573), .Y(n_572) );
BUFx8_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g576 ( .A(n_577), .B(n_863), .Y(n_576) );
NOR3xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_775), .C(n_811), .Y(n_577) );
NAND3xp33_ASAP7_75t_SL g578 ( .A(n_579), .B(n_708), .C(n_753), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_625), .B1(n_686), .B2(n_689), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g966 ( .A(n_581), .Y(n_966) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_598), .Y(n_581) );
INVx2_ASAP7_75t_L g728 ( .A(n_582), .Y(n_728) );
INVx2_ASAP7_75t_L g855 ( .A(n_582), .Y(n_855) );
INVx2_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g707 ( .A(n_583), .B(n_599), .Y(n_707) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_592), .Y(n_583) );
NAND2x1p5_ASAP7_75t_L g723 ( .A(n_584), .B(n_592), .Y(n_723) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OA21x2_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B(n_596), .Y(n_592) );
INVx1_ASAP7_75t_L g622 ( .A(n_597), .Y(n_622) );
OR2x2_ASAP7_75t_L g803 ( .A(n_598), .B(n_804), .Y(n_803) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_598), .Y(n_951) );
NAND2x1_ASAP7_75t_L g598 ( .A(n_599), .B(n_614), .Y(n_598) );
AND2x2_ASAP7_75t_L g749 ( .A(n_599), .B(n_723), .Y(n_749) );
AND2x2_ASAP7_75t_L g895 ( .A(n_599), .B(n_731), .Y(n_895) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B(n_609), .Y(n_606) );
OR2x2_ASAP7_75t_L g630 ( .A(n_611), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g681 ( .A(n_612), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g721 ( .A(n_614), .Y(n_721) );
INVx1_ASAP7_75t_L g740 ( .A(n_614), .Y(n_740) );
AND2x2_ASAP7_75t_L g748 ( .A(n_614), .B(n_693), .Y(n_748) );
AND2x2_ASAP7_75t_L g884 ( .A(n_614), .B(n_764), .Y(n_884) );
INVx3_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g756 ( .A(n_615), .B(n_724), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_618), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g960 ( .A(n_626), .Y(n_960) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_655), .Y(n_626) );
OR2x2_ASAP7_75t_L g814 ( .A(n_627), .B(n_734), .Y(n_814) );
OR2x2_ASAP7_75t_SL g924 ( .A(n_627), .B(n_925), .Y(n_924) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g686 ( .A(n_628), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g868 ( .A(n_628), .B(n_827), .Y(n_868) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_641), .Y(n_628) );
INVx2_ASAP7_75t_SL g746 ( .A(n_629), .Y(n_746) );
AND2x2_ASAP7_75t_L g752 ( .A(n_629), .B(n_642), .Y(n_752) );
OAI21x1_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .B(n_639), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g715 ( .A1(n_630), .A2(n_632), .B(n_639), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_631), .B(n_659), .Y(n_658) );
AOI21x1_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B(n_638), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_638), .B(n_703), .Y(n_704) );
INVx1_ASAP7_75t_L g790 ( .A(n_641), .Y(n_790) );
AND2x2_ASAP7_75t_L g874 ( .A(n_641), .B(n_675), .Y(n_874) );
INVx3_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g712 ( .A(n_642), .Y(n_712) );
AND2x2_ASAP7_75t_L g745 ( .A(n_642), .B(n_746), .Y(n_745) );
AND2x4_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
OAI21x1_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_649), .B(n_653), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B(n_652), .Y(n_649) );
INVx2_ASAP7_75t_L g678 ( .A(n_654), .Y(n_678) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g751 ( .A(n_656), .B(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_656), .B(n_852), .Y(n_851) );
NAND2x1_ASAP7_75t_SL g889 ( .A(n_656), .B(n_745), .Y(n_889) );
HB1xp67_ASAP7_75t_L g900 ( .A(n_656), .Y(n_900) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_675), .Y(n_656) );
INVx1_ASAP7_75t_L g688 ( .A(n_657), .Y(n_688) );
INVxp67_ASAP7_75t_L g711 ( .A(n_657), .Y(n_711) );
OR2x2_ASAP7_75t_L g736 ( .A(n_657), .B(n_715), .Y(n_736) );
INVx1_ASAP7_75t_L g798 ( .A(n_657), .Y(n_798) );
INVx1_ASAP7_75t_L g810 ( .A(n_657), .Y(n_810) );
AND2x2_ASAP7_75t_L g845 ( .A(n_657), .B(n_746), .Y(n_845) );
AO21x2_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_661), .B(n_673), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND3xp33_ASAP7_75t_SL g661 ( .A(n_662), .B(n_665), .C(n_668), .Y(n_661) );
AND2x2_ASAP7_75t_L g687 ( .A(n_675), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g716 ( .A(n_675), .Y(n_716) );
INVx1_ASAP7_75t_L g734 ( .A(n_675), .Y(n_734) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_675), .Y(n_779) );
NOR2x1_ASAP7_75t_L g809 ( .A(n_675), .B(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g828 ( .A(n_675), .Y(n_828) );
INVx1_ASAP7_75t_L g831 ( .A(n_675), .Y(n_831) );
OR2x6_ASAP7_75t_L g675 ( .A(n_676), .B(n_683), .Y(n_675) );
OAI21x1_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_679), .B(n_681), .Y(n_676) );
NOR2xp67_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
AND2x2_ASAP7_75t_L g827 ( .A(n_688), .B(n_828), .Y(n_827) );
AND2x4_ASAP7_75t_L g689 ( .A(n_690), .B(n_707), .Y(n_689) );
BUFx3_ASAP7_75t_L g758 ( .A(n_690), .Y(n_758) );
INVx3_ASAP7_75t_L g856 ( .A(n_690), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_690), .B(n_762), .Y(n_956) );
AND2x4_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
OR2x2_ASAP7_75t_L g730 ( .A(n_691), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g774 ( .A(n_691), .B(n_731), .Y(n_774) );
INVx1_ASAP7_75t_L g860 ( .A(n_691), .Y(n_860) );
INVx1_ASAP7_75t_L g850 ( .A(n_692), .Y(n_850) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVxp67_ASAP7_75t_L g761 ( .A(n_693), .Y(n_761) );
INVx1_ASAP7_75t_L g842 ( .A(n_693), .Y(n_842) );
AO21x2_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_699), .B(n_705), .Y(n_693) );
AO21x2_ASAP7_75t_L g731 ( .A1(n_694), .A2(n_699), .B(n_705), .Y(n_731) );
OAI21x1_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B(n_698), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI21x1_ASAP7_75t_SL g699 ( .A1(n_700), .A2(n_701), .B(n_704), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g706 ( .A(n_703), .Y(n_706) );
INVx1_ASAP7_75t_L g767 ( .A(n_707), .Y(n_767) );
AND2x2_ASAP7_75t_L g880 ( .A(n_707), .B(n_881), .Y(n_880) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_707), .Y(n_913) );
NOR2xp67_ASAP7_75t_SL g918 ( .A(n_707), .B(n_856), .Y(n_918) );
INVx1_ASAP7_75t_L g946 ( .A(n_707), .Y(n_946) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_717), .B1(n_726), .B2(n_732), .C(n_737), .Y(n_708) );
INVx2_ASAP7_75t_L g888 ( .A(n_709), .Y(n_888) );
AND2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_713), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_711), .Y(n_800) );
AND2x2_ASAP7_75t_L g733 ( .A(n_712), .B(n_734), .Y(n_733) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_712), .Y(n_771) );
INVx2_ASAP7_75t_L g852 ( .A(n_712), .Y(n_852) );
OR2x2_ASAP7_75t_L g869 ( .A(n_712), .B(n_736), .Y(n_869) );
AND2x2_ASAP7_75t_L g952 ( .A(n_713), .B(n_953), .Y(n_952) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .Y(n_713) );
BUFx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_716), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_716), .B(n_845), .Y(n_969) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .Y(n_719) );
AND2x2_ASAP7_75t_L g786 ( .A(n_720), .B(n_741), .Y(n_786) );
INVx1_ASAP7_75t_L g892 ( .A(n_720), .Y(n_892) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g921 ( .A(n_721), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_722), .Y(n_922) );
INVx2_ASAP7_75t_L g964 ( .A(n_722), .Y(n_964) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx2_ASAP7_75t_L g764 ( .A(n_723), .Y(n_764) );
INVx1_ASAP7_75t_L g785 ( .A(n_723), .Y(n_785) );
INVx1_ASAP7_75t_L g819 ( .A(n_723), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_723), .B(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g762 ( .A(n_724), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_724), .B(n_764), .Y(n_908) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g742 ( .A(n_725), .Y(n_742) );
OAI31xp33_ASAP7_75t_L g948 ( .A1(n_726), .A2(n_949), .A3(n_950), .B(n_952), .Y(n_948) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND2x1_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
AND3x2_ASAP7_75t_L g760 ( .A(n_728), .B(n_761), .C(n_762), .Y(n_760) );
AND2x2_ASAP7_75t_L g773 ( .A(n_728), .B(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g781 ( .A(n_730), .B(n_762), .Y(n_781) );
INVx2_ASAP7_75t_L g881 ( .A(n_730), .Y(n_881) );
AND2x4_ASAP7_75t_L g741 ( .A(n_731), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g768 ( .A(n_732), .Y(n_768) );
AND2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_735), .Y(n_732) );
NAND2x2_ASAP7_75t_L g843 ( .A(n_733), .B(n_844), .Y(n_843) );
AND2x2_ASAP7_75t_L g744 ( .A(n_734), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g770 ( .A(n_735), .B(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g780 ( .A(n_736), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_743), .B1(n_747), .B2(n_750), .Y(n_737) );
INVx2_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
NAND2xp67_ASAP7_75t_L g816 ( .A(n_739), .B(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g822 ( .A(n_739), .Y(n_822) );
AND2x4_ASAP7_75t_SL g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g837 ( .A(n_740), .Y(n_837) );
AND2x2_ASAP7_75t_L g943 ( .A(n_740), .B(n_749), .Y(n_943) );
AND2x2_ASAP7_75t_L g763 ( .A(n_741), .B(n_764), .Y(n_763) );
BUFx3_ASAP7_75t_L g797 ( .A(n_741), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_741), .B(n_884), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_742), .B(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g865 ( .A1(n_744), .A2(n_763), .B1(n_866), .B2(n_870), .C(n_871), .Y(n_865) );
INVx1_ASAP7_75t_L g791 ( .A(n_746), .Y(n_791) );
INVx1_ASAP7_75t_L g931 ( .A(n_746), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
AND2x2_ASAP7_75t_L g832 ( .A(n_749), .B(n_761), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_749), .B(n_837), .Y(n_836) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_751), .Y(n_765) );
INVx2_ASAP7_75t_L g806 ( .A(n_752), .Y(n_806) );
AND2x2_ASAP7_75t_L g902 ( .A(n_752), .B(n_903), .Y(n_902) );
O2A1O1Ixp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_763), .B(n_765), .C(n_766), .Y(n_753) );
NAND3xp33_ASAP7_75t_SL g754 ( .A(n_755), .B(n_757), .C(n_759), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2x1p5_ASAP7_75t_L g848 ( .A(n_756), .B(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g804 ( .A(n_761), .Y(n_804) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_761), .Y(n_915) );
OR2x2_ASAP7_75t_L g911 ( .A(n_762), .B(n_841), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_768), .B1(n_769), .B2(n_772), .Y(n_766) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g929 ( .A(n_771), .B(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g958 ( .A(n_774), .Y(n_958) );
OAI221xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_781), .B1(n_782), .B2(n_787), .C(n_792), .Y(n_775) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
AND2x2_ASAP7_75t_L g830 ( .A(n_780), .B(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g875 ( .A(n_780), .Y(n_875) );
AOI21xp33_ASAP7_75t_L g926 ( .A1(n_781), .A2(n_927), .B(n_928), .Y(n_926) );
INVxp67_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_784), .B(n_786), .Y(n_783) );
AND2x2_ASAP7_75t_L g793 ( .A(n_784), .B(n_794), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_784), .B(n_858), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_784), .A2(n_855), .B1(n_867), .B2(n_869), .Y(n_866) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g898 ( .A(n_788), .Y(n_898) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NOR2xp67_ASAP7_75t_SL g834 ( .A(n_789), .B(n_798), .Y(n_834) );
OR2x2_ASAP7_75t_L g861 ( .A(n_789), .B(n_862), .Y(n_861) );
OR2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
INVx1_ASAP7_75t_L g794 ( .A(n_790), .Y(n_794) );
INVxp67_ASAP7_75t_SL g825 ( .A(n_791), .Y(n_825) );
A2O1A1Ixp33_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_795), .B(n_798), .C(n_799), .Y(n_792) );
INVx1_ASAP7_75t_L g940 ( .A(n_794), .Y(n_940) );
INVxp67_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_796), .B(n_872), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g910 ( .A1(n_796), .A2(n_843), .B1(n_901), .B2(n_911), .Y(n_910) );
INVx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g879 ( .A(n_798), .Y(n_879) );
AND2x2_ASAP7_75t_L g930 ( .A(n_798), .B(n_931), .Y(n_930) );
AND2x2_ASAP7_75t_L g953 ( .A(n_798), .B(n_852), .Y(n_953) );
AOI21xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_801), .B(n_807), .Y(n_799) );
INVx1_ASAP7_75t_L g903 ( .A(n_800), .Y(n_903) );
NAND2xp5_ASAP7_75t_SL g801 ( .A(n_802), .B(n_805), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
AOI221xp5_ASAP7_75t_L g876 ( .A1(n_806), .A2(n_877), .B1(n_882), .B2(n_885), .C(n_887), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_807), .B(n_852), .Y(n_942) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
OR2x2_ASAP7_75t_L g886 ( .A(n_808), .B(n_852), .Y(n_886) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
NAND3xp33_ASAP7_75t_SL g811 ( .A(n_812), .B(n_820), .C(n_833), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_815), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_817), .B(n_847), .Y(n_934) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
AOI21x1_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_823), .B(n_829), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
OR2x2_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
AND2x2_ASAP7_75t_L g829 ( .A(n_830), .B(n_832), .Y(n_829) );
AOI221xp5_ASAP7_75t_L g954 ( .A1(n_830), .A2(n_955), .B1(n_957), .B2(n_960), .C(n_961), .Y(n_954) );
INVx2_ASAP7_75t_L g925 ( .A(n_831), .Y(n_925) );
AOI211xp5_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_835), .B(n_838), .C(n_853), .Y(n_833) );
INVxp67_ASAP7_75t_SL g835 ( .A(n_836), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_839), .A2(n_843), .B1(n_846), .B2(n_851), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
BUFx3_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
AND2x4_ASAP7_75t_L g947 ( .A(n_845), .B(n_874), .Y(n_947) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
AOI211xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_856), .B(n_857), .C(n_861), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
OR2x2_ASAP7_75t_L g927 ( .A(n_855), .B(n_894), .Y(n_927) );
AND2x2_ASAP7_75t_L g949 ( .A(n_855), .B(n_895), .Y(n_949) );
INVx1_ASAP7_75t_L g870 ( .A(n_857), .Y(n_870) );
INVx2_ASAP7_75t_SL g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g909 ( .A(n_860), .Y(n_909) );
NOR2xp67_ASAP7_75t_L g863 ( .A(n_864), .B(n_916), .Y(n_863) );
NAND3xp33_ASAP7_75t_L g864 ( .A(n_865), .B(n_876), .C(n_896), .Y(n_864) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
OR2x2_ASAP7_75t_L g872 ( .A(n_873), .B(n_875), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_881), .B(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
AOI21xp33_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .B(n_890), .Y(n_887) );
NOR3xp33_ASAP7_75t_L g912 ( .A(n_888), .B(n_913), .C(n_914), .Y(n_912) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_892), .B(n_893), .Y(n_891) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
NOR3xp33_ASAP7_75t_L g896 ( .A(n_897), .B(n_910), .C(n_912), .Y(n_896) );
O2A1O1Ixp33_ASAP7_75t_L g897 ( .A1(n_898), .A2(n_899), .B(n_901), .C(n_904), .Y(n_897) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_907), .B(n_909), .Y(n_906) );
INVxp67_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
NAND4xp25_ASAP7_75t_SL g916 ( .A(n_917), .B(n_932), .C(n_948), .D(n_954), .Y(n_916) );
O2A1O1Ixp33_ASAP7_75t_SL g917 ( .A1(n_918), .A2(n_919), .B(n_923), .C(n_926), .Y(n_917) );
INVxp67_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
OR2x2_ASAP7_75t_L g920 ( .A(n_921), .B(n_922), .Y(n_920) );
OR2x2_ASAP7_75t_L g945 ( .A(n_921), .B(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx2_ASAP7_75t_L g938 ( .A(n_925), .Y(n_938) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
AOI222xp33_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_935), .B1(n_941), .B2(n_943), .C1(n_944), .C2(n_947), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
NOR2xp33_ASAP7_75t_L g935 ( .A(n_936), .B(n_939), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g959 ( .A(n_943), .Y(n_959) );
INVx2_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVxp67_ASAP7_75t_SL g950 ( .A(n_951), .Y(n_950) );
INVxp67_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_958), .B(n_959), .Y(n_957) );
AOI21xp33_ASAP7_75t_L g961 ( .A1(n_962), .A2(n_965), .B(n_967), .Y(n_961) );
INVx2_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
NOR2xp33_ASAP7_75t_L g973 ( .A(n_974), .B(n_975), .Y(n_973) );
BUFx2_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
BUFx2_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
BUFx3_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
BUFx4_ASAP7_75t_SL g980 ( .A(n_981), .Y(n_980) );
BUFx3_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
BUFx3_ASAP7_75t_L g990 ( .A(n_982), .Y(n_990) );
AND2x4_ASAP7_75t_L g982 ( .A(n_983), .B(n_985), .Y(n_982) );
CKINVDCx20_ASAP7_75t_R g983 ( .A(n_984), .Y(n_983) );
CKINVDCx6p67_ASAP7_75t_R g988 ( .A(n_989), .Y(n_988) );
BUFx2_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
endmodule