module fake_jpeg_14978_n_116 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_116);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_28),
.Y(n_40)
);

NOR2xp67_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_2),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_3),
.B(n_4),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_28),
.Y(n_42)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_3),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_13),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_15),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_42),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_26),
.A2(n_15),
.B1(n_24),
.B2(n_25),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_45),
.B1(n_24),
.B2(n_12),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_26),
.A2(n_18),
.B1(n_13),
.B2(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_49),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_32),
.B1(n_30),
.B2(n_12),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_36),
.B1(n_44),
.B2(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_40),
.B(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_48),
.B(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_18),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_31),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_54),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_60),
.B1(n_16),
.B2(n_23),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_30),
.B1(n_32),
.B2(n_36),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_33),
.B1(n_19),
.B2(n_6),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_33),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_21),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_33),
.B(n_5),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_68),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_73),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_74),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_57),
.B(n_60),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_53),
.B1(n_52),
.B2(n_54),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_52),
.C(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_51),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_69),
.B1(n_21),
.B2(n_6),
.Y(n_90)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_59),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_62),
.B(n_66),
.Y(n_87)
);

A2O1A1O1Ixp25_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_61),
.B(n_21),
.C(n_17),
.D(n_7),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_3),
.B(n_5),
.Y(n_94)
);

OAI321xp33_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_62),
.A3(n_66),
.B1(n_71),
.B2(n_70),
.C(n_65),
.Y(n_86)
);

NOR3xp33_ASAP7_75t_SL g96 ( 
.A(n_86),
.B(n_91),
.C(n_84),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_75),
.C(n_82),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_94),
.B(n_6),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_69),
.C(n_9),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_92),
.B(n_82),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_88),
.C(n_83),
.Y(n_101)
);

OAI221xp5_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_94),
.C(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_99),
.Y(n_103)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_10),
.C(n_8),
.Y(n_107)
);

XNOR2x1_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_87),
.Y(n_102)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_102),
.B(n_85),
.CI(n_8),
.CON(n_106),
.SN(n_106)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_104),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_103),
.B(n_104),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_10),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_109),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

AOI21x1_ASAP7_75t_L g113 ( 
.A1(n_111),
.A2(n_108),
.B(n_106),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_107),
.C(n_8),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_114),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_110),
.Y(n_116)
);


endmodule