module real_jpeg_5611_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_1),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_2),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_2),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_2),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_2),
.B(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_2),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_2),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_2),
.B(n_389),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_3),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_3),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_3),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_3),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_3),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_4),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_4),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_4),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_4),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_4),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_4),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_5),
.B(n_90),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_5),
.A2(n_115),
.B(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_5),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_5),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_5),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_5),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_5),
.B(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_5),
.B(n_369),
.Y(n_396)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_7),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_7),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_7),
.Y(n_306)
);

BUFx5_ASAP7_75t_L g369 ( 
.A(n_7),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_8),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_8),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_8),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_8),
.B(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_8),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_8),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_8),
.B(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_9),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_9),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_9),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_9),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_9),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_9),
.B(n_358),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_9),
.B(n_393),
.Y(n_392)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_10),
.Y(n_116)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_10),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g300 ( 
.A(n_10),
.Y(n_300)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_12),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_12),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_12),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_12),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_12),
.B(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_12),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_12),
.B(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_12),
.B(n_410),
.Y(n_409)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_13),
.Y(n_121)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_13),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_13),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_14),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_14),
.Y(n_358)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_14),
.Y(n_413)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_15),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_15),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_15),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_15),
.B(n_85),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_15),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_204),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_202),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_169),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_19),
.B(n_169),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_97),
.C(n_125),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_20),
.B(n_97),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_59),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_41),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_22),
.B(n_41),
.C(n_59),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.C(n_39),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_23),
.B(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_26),
.C(n_31),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_24),
.B(n_51),
.C(n_55),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_24),
.A2(n_55),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_24),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_24),
.A2(n_31),
.B1(n_93),
.B2(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_24),
.A2(n_93),
.B1(n_371),
.B2(n_373),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_24),
.B(n_373),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_26),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_26),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_26),
.A2(n_128),
.B1(n_197),
.B2(n_201),
.Y(n_196)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_30),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_30),
.Y(n_229)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_30),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_31),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_31),
.B(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_31),
.A2(n_131),
.B1(n_265),
.B2(n_266),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_32),
.Y(n_365)
);

INVx8_ASAP7_75t_L g387 ( 
.A(n_32),
.Y(n_387)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g395 ( 
.A(n_33),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_34),
.A2(n_39),
.B1(n_49),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_34),
.Y(n_168)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_38),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_43),
.B1(n_44),
.B2(n_49),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_50),
.B1(n_57),
.B2(n_58),
.Y(n_41)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_44),
.B(n_49),
.C(n_58),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_47),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_47),
.Y(n_219)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_48),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_48),
.Y(n_312)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_51),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_51),
.B(n_227),
.C(n_230),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_51),
.A2(n_95),
.B1(n_227),
.B2(n_295),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_79),
.C(n_91),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_60),
.B(n_79),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_66),
.B2(n_67),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_69),
.C(n_74),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_61),
.A2(n_62),
.B1(n_120),
.B2(n_122),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_61),
.B(n_120),
.C(n_124),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_61),
.A2(n_62),
.B1(n_146),
.B2(n_147),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_62),
.B(n_147),
.Y(n_303)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_74),
.B2(n_78),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_71),
.Y(n_160)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx6_ASAP7_75t_L g331 ( 
.A(n_72),
.Y(n_331)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_73),
.Y(n_178)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_73),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_73),
.Y(n_355)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.C(n_87),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_80),
.B(n_143),
.Y(n_142)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_84),
.B(n_87),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_86),
.Y(n_243)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_91),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_117),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_99),
.B(n_100),
.C(n_117),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_111),
.B2(n_112),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_105),
.B1(n_109),
.B2(n_110),
.Y(n_102)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_105),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_105),
.B(n_109),
.C(n_112),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_105),
.B(n_134),
.Y(n_213)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_133),
.C(n_138),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_116),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_123),
.B2(n_124),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_120),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_123),
.A2(n_124),
.B1(n_181),
.B2(n_184),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_123),
.B(n_257),
.C(n_261),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_123),
.A2(n_124),
.B1(n_261),
.B2(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_125),
.B(n_286),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_144),
.C(n_166),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_126),
.B(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_132),
.C(n_142),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_127),
.Y(n_250)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_132),
.B(n_142),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_138),
.B(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_144),
.B(n_166),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_159),
.C(n_161),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_145),
.B(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_152),
.C(n_158),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_146),
.A2(n_147),
.B1(n_158),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_151),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_152),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_152),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_157),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_158),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_159),
.A2(n_161),
.B1(n_162),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_159),
.Y(n_248)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_165),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g447 ( 
.A(n_169),
.Y(n_447)
);

FAx1_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_171),
.CI(n_185),
.CON(n_169),
.SN(n_169)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_215),
.C(n_220),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_176),
.A2(n_177),
.B1(n_215),
.B2(n_216),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_181),
.Y(n_184)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI221xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_344),
.B1(n_439),
.B2(n_444),
.C(n_445),
.Y(n_205)
);

NOR3xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_283),
.C(n_287),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_207),
.A2(n_440),
.B(n_443),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_276),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_208),
.B(n_276),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_249),
.C(n_252),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_209),
.B(n_249),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_234),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_210),
.B(n_235),
.C(n_246),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.C(n_225),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_212),
.B(n_226),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_214),
.B(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_220),
.B(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g372 ( 
.A(n_224),
.Y(n_372)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_230),
.B(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_246),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_241),
.C(n_244),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_275),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_236),
.A2(n_237),
.B(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_244),
.Y(n_275)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_243),
.B(n_298),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_252),
.B(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_269),
.C(n_274),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_253),
.B(n_291),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.C(n_263),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_254),
.B(n_340),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_256),
.A2(n_263),
.B1(n_264),
.B2(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_256),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_257),
.B(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_261),
.Y(n_324)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_274),
.Y(n_291)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_280),
.C(n_282),
.Y(n_284)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_283),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_284),
.B(n_285),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_317),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_288),
.A2(n_441),
.B(n_442),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_315),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_289),
.B(n_315),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.C(n_313),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_290),
.B(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_313),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_296),
.C(n_301),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_296),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.C(n_307),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_302),
.A2(n_303),
.B1(n_427),
.B2(n_428),
.Y(n_426)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_304),
.A2(n_305),
.B1(n_307),
.B2(n_308),
.Y(n_427)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_312),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_342),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_318),
.B(n_342),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_321),
.C(n_339),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_319),
.B(n_437),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_321),
.B(n_339),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_325),
.C(n_337),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_322),
.B(n_430),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_325),
.A2(n_337),
.B1(n_338),
.B2(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_325),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.C(n_332),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_326),
.A2(n_327),
.B1(n_332),
.B2(n_333),
.Y(n_419)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_329),
.B(n_419),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_330),
.B(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_331),
.Y(n_380)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_345),
.A2(n_434),
.B(n_438),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_421),
.B(n_433),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_405),
.B(n_420),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_381),
.B(n_404),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_349),
.B(n_374),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_349),
.B(n_374),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_361),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_350),
.B(n_362),
.C(n_370),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_356),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_351),
.B(n_357),
.C(n_359),
.Y(n_417)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_359),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_370),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_366),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_366),
.Y(n_375)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_371),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.C(n_377),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_401),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_376),
.A2(n_377),
.B1(n_378),
.B2(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_376),
.Y(n_402)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_398),
.B(n_403),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_391),
.B(n_397),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_390),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_384),
.B(n_390),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_388),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_385),
.B(n_388),
.Y(n_399)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_396),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_394),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_400),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_407),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_416),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_408),
.A2(n_424),
.B1(n_425),
.B2(n_426),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_408),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_408),
.B(n_417),
.C(n_418),
.Y(n_432)
);

FAx1_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_414),
.CI(n_415),
.CON(n_408),
.SN(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_422),
.B(n_432),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_422),
.B(n_432),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_429),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_426),
.C(n_429),
.Y(n_435)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_427),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_436),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_435),
.B(n_436),
.Y(n_438)
);


endmodule