module real_jpeg_12137_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_97;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_3),
.A2(n_25),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_3),
.A2(n_31),
.B1(n_43),
.B2(n_44),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_5),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_109),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_109),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_5),
.A2(n_25),
.B1(n_32),
.B2(n_109),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_7),
.A2(n_62),
.B1(n_63),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_7),
.A2(n_57),
.B1(n_58),
.B2(n_67),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_67),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_7),
.A2(n_25),
.B1(n_32),
.B2(n_67),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_8),
.A2(n_56),
.B(n_62),
.C(n_101),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_8),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_8),
.A2(n_62),
.B1(n_63),
.B2(n_102),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_8),
.B(n_131),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_8),
.B(n_57),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_SL g201 ( 
.A1(n_8),
.A2(n_57),
.B(n_187),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_8),
.B(n_25),
.C(n_39),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_102),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_8),
.A2(n_24),
.B1(n_27),
.B2(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_8),
.B(n_80),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_9),
.A2(n_62),
.B1(n_63),
.B2(n_69),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_9),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_9),
.A2(n_57),
.B1(n_58),
.B2(n_69),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_69),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_9),
.A2(n_25),
.B1(n_32),
.B2(n_69),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_10),
.A2(n_25),
.B1(n_32),
.B2(n_46),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_10),
.A2(n_46),
.B1(n_57),
.B2(n_58),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_13),
.A2(n_25),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_13),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_13),
.A2(n_36),
.B1(n_57),
.B2(n_58),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_14),
.A2(n_57),
.B1(n_58),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_14),
.A2(n_25),
.B1(n_32),
.B2(n_72),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_14),
.A2(n_62),
.B1(n_63),
.B2(n_72),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_72),
.Y(n_152)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_137),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_110),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_20),
.B(n_110),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.C(n_94),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_21),
.B(n_82),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_51),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_22),
.B(n_52),
.C(n_81),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_23),
.B(n_37),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B(n_33),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_24),
.B(n_35),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_24),
.A2(n_27),
.B(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_24),
.A2(n_27),
.B1(n_216),
.B2(n_224),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_24),
.A2(n_86),
.B(n_218),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_25),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_32),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_27),
.B(n_102),
.Y(n_222)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_28),
.B(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_28),
.A2(n_30),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_28),
.A2(n_88),
.B(n_98),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_28),
.A2(n_97),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_32),
.B(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_34),
.A2(n_87),
.B(n_97),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B(n_47),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_38),
.B(n_102),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_42),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_43),
.A2(n_44),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_SL g188 ( 
.A(n_43),
.B(n_58),
.C(n_75),
.Y(n_188)
);

INVx5_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_44),
.A2(n_76),
.B(n_186),
.C(n_188),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_44),
.B(n_210),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_48),
.B(n_91),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_49),
.A2(n_92),
.B(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_49),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_49),
.A2(n_91),
.B1(n_181),
.B2(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_49),
.A2(n_91),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_49),
.A2(n_91),
.B1(n_203),
.B2(n_213),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_70),
.B2(n_81),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_66),
.B2(n_68),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_54),
.A2(n_55),
.B1(n_66),
.B2(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_54),
.A2(n_68),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_54),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_61),
.Y(n_54)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_56),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_58),
.B1(n_75),
.B2(n_76),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_57),
.A2(n_60),
.B(n_102),
.Y(n_101)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_73),
.B(n_78),
.Y(n_70)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_73),
.A2(n_74),
.B1(n_104),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_73),
.A2(n_74),
.B1(n_147),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_73),
.A2(n_74),
.B1(n_163),
.B2(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_74),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_79),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_89),
.B2(n_93),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_93),
.Y(n_122)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_91),
.B(n_152),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_94),
.B(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_103),
.C(n_107),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_95),
.B(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_96),
.A2(n_99),
.B1(n_100),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_103),
.B(n_107),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_108),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_135),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_120),
.B1(n_133),
.B2(n_134),
.Y(n_111)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_119),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_131),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_170),
.B(n_249),
.C(n_253),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_164),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_139),
.B(n_164),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_154),
.C(n_157),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_148),
.C(n_153),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_148),
.B1(n_149),
.B2(n_153),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_150),
.A2(n_180),
.B(n_182),
.Y(n_179)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_162),
.B(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_165),
.B(n_168),
.C(n_169),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_247),
.B(n_248),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_191),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_173),
.B(n_176),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.C(n_183),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_179),
.A2(n_183),
.B1(n_184),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_189),
.B1(n_190),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_204),
.B(n_246),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_193),
.B(n_196),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.C(n_202),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_240),
.B(n_245),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_230),
.B(n_239),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_219),
.B(n_229),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_214),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_214),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_211),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_225),
.B(n_228),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_227),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_232),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_235),
.C(n_238),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_237),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_244),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_252),
.Y(n_253)
);


endmodule