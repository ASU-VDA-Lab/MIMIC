module fake_jpeg_13060_n_397 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_397);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_397;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_43),
.B(n_48),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_44),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_47),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_49),
.B(n_50),
.Y(n_120)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_51),
.Y(n_131)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_52),
.B(n_54),
.Y(n_121)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_17),
.B(n_14),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_17),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_55),
.B(n_57),
.Y(n_123)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_1),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_61),
.B(n_63),
.Y(n_94)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

BUFx12f_ASAP7_75t_SL g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_67),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_68),
.Y(n_96)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_18),
.B(n_13),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_69),
.B(n_70),
.Y(n_124)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_71),
.Y(n_87)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_72),
.B(n_73),
.Y(n_95)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_74),
.B(n_76),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_25),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_79),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_80),
.Y(n_92)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_38),
.B1(n_34),
.B2(n_28),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_25),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_83),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_24),
.Y(n_82)
);

HAxp5_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_40),
.CON(n_102),
.SN(n_102)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_24),
.B(n_1),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_5),
.C(n_6),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_37),
.B1(n_23),
.B2(n_41),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_86),
.A2(n_103),
.B1(n_104),
.B2(n_113),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_41),
.B1(n_20),
.B2(n_37),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_107),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_41),
.B1(n_40),
.B2(n_39),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_51),
.A2(n_41),
.B1(n_28),
.B2(n_38),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_98),
.A2(n_100),
.B1(n_116),
.B2(n_94),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_102),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_63),
.A2(n_34),
.B1(n_27),
.B2(n_22),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_72),
.A2(n_29),
.B1(n_27),
.B2(n_22),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_66),
.A2(n_29),
.B1(n_27),
.B2(n_22),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_105),
.A2(n_107),
.B1(n_90),
.B2(n_126),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_39),
.B1(n_36),
.B2(n_33),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_76),
.A2(n_36),
.B1(n_33),
.B2(n_32),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_110),
.A2(n_119),
.B1(n_127),
.B2(n_87),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_32),
.B1(n_29),
.B2(n_4),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_111),
.A2(n_115),
.B1(n_126),
.B2(n_131),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_56),
.A2(n_62),
.B1(n_47),
.B2(n_70),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_83),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_114),
.A2(n_125),
.B1(n_129),
.B2(n_100),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_82),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_115)
);

HAxp5_ASAP7_75t_SL g117 ( 
.A(n_52),
.B(n_44),
.CON(n_117),
.SN(n_117)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_117),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_60),
.B(n_2),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_119),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_71),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_88),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_71),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_44),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_60),
.A2(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_64),
.B(n_7),
.C(n_67),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_124),
.C(n_118),
.Y(n_136)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_135),
.B(n_140),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_136),
.B(n_160),
.C(n_169),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_163),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_138),
.A2(n_146),
.B1(n_151),
.B2(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_120),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_141),
.B(n_150),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_142),
.B(n_144),
.Y(n_187)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_92),
.B(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_124),
.B(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_145),
.B(n_91),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_122),
.A2(n_133),
.B1(n_95),
.B2(n_93),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_97),
.Y(n_150)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_95),
.A2(n_93),
.B1(n_105),
.B2(n_97),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_96),
.A2(n_91),
.B(n_94),
.C(n_100),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_156),
.B(n_169),
.Y(n_216)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_159),
.A2(n_174),
.B1(n_135),
.B2(n_149),
.Y(n_206)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_101),
.B(n_112),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_178),
.C(n_100),
.Y(n_186)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_85),
.Y(n_163)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_85),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_98),
.A2(n_127),
.B1(n_96),
.B2(n_108),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_172),
.B1(n_138),
.B2(n_155),
.Y(n_200)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_87),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_171),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_116),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_89),
.B1(n_99),
.B2(n_111),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_116),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_176),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_128),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_110),
.B(n_91),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_196),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_189),
.B(n_190),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_116),
.Y(n_190)
);

MAJx2_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_136),
.C(n_144),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_195),
.C(n_219),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_139),
.B(n_99),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_207),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_100),
.C(n_99),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_171),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_166),
.B1(n_134),
.B2(n_167),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_206),
.A2(n_201),
.B1(n_217),
.B2(n_216),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_146),
.B(n_148),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_153),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_211),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_175),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_165),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_177),
.Y(n_254)
);

AO22x1_ASAP7_75t_SL g217 ( 
.A1(n_168),
.A2(n_164),
.B1(n_156),
.B2(n_172),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_205),
.Y(n_241)
);

AOI32xp33_ASAP7_75t_L g218 ( 
.A1(n_164),
.A2(n_157),
.A3(n_174),
.B1(n_173),
.B2(n_143),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_206),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_188),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_222),
.B(n_240),
.Y(n_272)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_226),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_192),
.A2(n_167),
.B1(n_152),
.B2(n_158),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_187),
.B(n_162),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_227),
.B(n_244),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_192),
.A2(n_147),
.B1(n_179),
.B2(n_173),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_228),
.B(n_229),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_207),
.A2(n_173),
.B1(n_217),
.B2(n_214),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_230),
.A2(n_241),
.B1(n_231),
.B2(n_220),
.Y(n_263)
);

AO21x1_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_189),
.B(n_184),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_231),
.A2(n_232),
.B(n_230),
.Y(n_278)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_180),
.A2(n_216),
.B1(n_201),
.B2(n_211),
.Y(n_236)
);

INVxp33_ASAP7_75t_SL g271 ( 
.A(n_236),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_196),
.A2(n_183),
.B(n_187),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_237),
.A2(n_239),
.B(n_235),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_180),
.A2(n_194),
.B1(n_219),
.B2(n_191),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_238),
.A2(n_243),
.B1(n_245),
.B2(n_253),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_197),
.A2(n_204),
.B(n_195),
.Y(n_239)
);

OAI32xp33_ASAP7_75t_L g240 ( 
.A1(n_205),
.A2(n_185),
.A3(n_209),
.B1(n_210),
.B2(n_203),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_209),
.A2(n_202),
.B1(n_210),
.B2(n_182),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_185),
.B(n_203),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_202),
.A2(n_182),
.B1(n_213),
.B2(n_199),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_213),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_248),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_198),
.C(n_193),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_249),
.C(n_232),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_193),
.B(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_187),
.B(n_214),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_250),
.B(n_251),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_187),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_181),
.Y(n_252)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_200),
.A2(n_218),
.B1(n_192),
.B2(n_207),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_242),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_235),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_258),
.B(n_267),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_238),
.C(n_251),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_259),
.B(n_265),
.C(n_268),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_260),
.B(n_275),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_274),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_239),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_278),
.C(n_284),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_220),
.C(n_229),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_244),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_237),
.C(n_253),
.Y(n_268)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_246),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_241),
.A2(n_221),
.B(n_254),
.Y(n_276)
);

AO21x1_ASAP7_75t_L g300 ( 
.A1(n_276),
.A2(n_252),
.B(n_233),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_243),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_279),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_248),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_222),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_281),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_221),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_283),
.B(n_247),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_260),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_287),
.B(n_301),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_228),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_290),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_261),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_302),
.Y(n_314)
);

XOR2x1_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_268),
.Y(n_294)
);

XNOR2x1_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_309),
.Y(n_329)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_256),
.Y(n_296)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_256),
.Y(n_297)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_297),
.Y(n_315)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_262),
.Y(n_298)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_298),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_259),
.B(n_227),
.C(n_226),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_264),
.C(n_278),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_279),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_272),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_223),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_276),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_258),
.B(n_234),
.Y(n_305)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_305),
.Y(n_324)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_262),
.Y(n_306)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_306),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_308),
.B(n_284),
.Y(n_313)
);

NAND2x1_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_224),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_266),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_310),
.A2(n_266),
.B1(n_280),
.B2(n_269),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_311),
.B(n_316),
.C(n_321),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_313),
.B(n_326),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_273),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_301),
.A2(n_257),
.B1(n_271),
.B2(n_274),
.Y(n_320)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_320),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_273),
.C(n_282),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_289),
.A2(n_267),
.B1(n_255),
.B2(n_277),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_322),
.A2(n_289),
.B1(n_303),
.B2(n_290),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_323),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_282),
.C(n_257),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_299),
.C(n_302),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_327),
.B(n_330),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_328),
.A2(n_300),
.B(n_295),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_280),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_290),
.A2(n_255),
.B1(n_270),
.B2(n_269),
.Y(n_331)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_331),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_295),
.Y(n_332)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_332),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_334),
.A2(n_348),
.B(n_349),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_291),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_335),
.B(n_340),
.Y(n_354)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_336),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_320),
.Y(n_339)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_339),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_328),
.A2(n_287),
.B1(n_304),
.B2(n_290),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_303),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_343),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_305),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_346),
.Y(n_358)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

AOI322xp5_ASAP7_75t_L g346 ( 
.A1(n_319),
.A2(n_292),
.A3(n_294),
.B1(n_308),
.B2(n_300),
.C1(n_302),
.C2(n_309),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_331),
.B(n_293),
.Y(n_348)
);

AO221x1_ASAP7_75t_L g349 ( 
.A1(n_312),
.A2(n_318),
.B1(n_315),
.B2(n_325),
.C(n_306),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_337),
.B(n_316),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_350),
.B(n_362),
.Y(n_364)
);

FAx1_ASAP7_75t_SL g355 ( 
.A(n_343),
.B(n_314),
.CI(n_327),
.CON(n_355),
.SN(n_355)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_355),
.B(n_314),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_330),
.C(n_311),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_359),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_321),
.C(n_313),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_341),
.B(n_294),
.C(n_329),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_333),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_334),
.B(n_329),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_363),
.A2(n_358),
.B(n_360),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_362),
.B(n_357),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_366),
.B(n_368),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_339),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_361),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_359),
.B(n_292),
.C(n_345),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_369),
.B(n_370),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_286),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_353),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_371),
.B(n_353),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_286),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_372),
.B(n_373),
.Y(n_379)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_358),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_364),
.B(n_350),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_364),
.C(n_366),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_377),
.B(n_380),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_378),
.A2(n_381),
.B(n_367),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_371),
.A2(n_351),
.B(n_356),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_340),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_382),
.B(n_351),
.Y(n_387)
);

NAND4xp25_ASAP7_75t_L g390 ( 
.A(n_384),
.B(n_352),
.C(n_332),
.D(n_338),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_379),
.A2(n_376),
.B(n_377),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_388),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_386),
.B(n_387),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_373),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_383),
.B(n_380),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_389),
.B(n_336),
.Y(n_394)
);

AOI322xp5_ASAP7_75t_L g393 ( 
.A1(n_390),
.A2(n_338),
.A3(n_342),
.B1(n_296),
.B2(n_297),
.C1(n_298),
.C2(n_310),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_393),
.B(n_394),
.Y(n_395)
);

OAI21xp33_ASAP7_75t_L g396 ( 
.A1(n_395),
.A2(n_391),
.B(n_392),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_396),
.B(n_392),
.Y(n_397)
);


endmodule