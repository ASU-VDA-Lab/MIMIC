module fake_jpeg_6973_n_298 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_182;
wire n_19;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_38),
.Y(n_51)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_45),
.A2(n_64),
.B1(n_28),
.B2(n_25),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_61),
.B1(n_30),
.B2(n_25),
.Y(n_78)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_52),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_71),
.B(n_19),
.C(n_17),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_56),
.B(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_59),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_23),
.B1(n_33),
.B2(n_20),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_18),
.B1(n_33),
.B2(n_20),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_34),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_70),
.B(n_39),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_37),
.B(n_31),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_37),
.A3(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_78),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_80),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_37),
.B1(n_41),
.B2(n_44),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_18),
.C(n_24),
.Y(n_82)
);

AO21x1_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_95),
.B(n_70),
.Y(n_107)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_19),
.B1(n_40),
.B2(n_37),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_56),
.A2(n_44),
.B1(n_31),
.B2(n_30),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_44),
.B1(n_40),
.B2(n_31),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_30),
.B1(n_28),
.B2(n_25),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_28),
.B1(n_66),
.B2(n_69),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_98),
.B(n_102),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_58),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_111),
.Y(n_148)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_107),
.Y(n_130)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_77),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_47),
.C(n_51),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_19),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_71),
.Y(n_106)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_52),
.Y(n_108)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_68),
.Y(n_109)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_63),
.Y(n_110)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_51),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_49),
.Y(n_113)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_91),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_114),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_61),
.Y(n_115)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_67),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_86),
.B1(n_87),
.B2(n_79),
.Y(n_147)
);

AO21x1_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_67),
.B(n_40),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_120),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_85),
.Y(n_121)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_85),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_118),
.C(n_103),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_53),
.B1(n_65),
.B2(n_55),
.Y(n_125)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_121),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_133),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_98),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_131),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_101),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_69),
.B1(n_66),
.B2(n_62),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_134),
.B(n_144),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_69),
.B1(n_66),
.B2(n_72),
.Y(n_140)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_19),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_141),
.A2(n_106),
.B(n_110),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_146),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_119),
.B1(n_75),
.B2(n_120),
.Y(n_171)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_150),
.Y(n_159)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

BUFx8_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_151),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_123),
.B(n_136),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_111),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_156),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_108),
.Y(n_156)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_172),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_139),
.A2(n_105),
.B(n_114),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_127),
.B(n_137),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_164),
.C(n_175),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_163),
.B(n_169),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_118),
.C(n_105),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_118),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_167),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_109),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_104),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_173),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_171),
.A2(n_123),
.B1(n_136),
.B2(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_104),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_128),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_174),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_113),
.C(n_79),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_179),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_128),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_177),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_107),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_141),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_132),
.B(n_107),
.Y(n_179)
);

AOI221xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_190),
.B1(n_151),
.B2(n_17),
.C(n_27),
.Y(n_214)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_186),
.Y(n_224)
);

AOI321xp33_ASAP7_75t_L g213 ( 
.A1(n_182),
.A2(n_156),
.A3(n_168),
.B1(n_17),
.B2(n_151),
.C(n_21),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_183),
.A2(n_17),
.B(n_21),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_135),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_184),
.A2(n_193),
.B(n_73),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_175),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_173),
.A2(n_127),
.B1(n_135),
.B2(n_132),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_165),
.Y(n_189)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_177),
.C(n_176),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_141),
.B1(n_129),
.B2(n_145),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_191),
.A2(n_196),
.B1(n_154),
.B2(n_163),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_161),
.A2(n_137),
.B(n_131),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_155),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_195),
.B(n_197),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_158),
.A2(n_129),
.B1(n_149),
.B2(n_120),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_153),
.Y(n_208)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_184),
.A2(n_164),
.A3(n_162),
.B1(n_166),
.B2(n_152),
.C1(n_154),
.C2(n_165),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_210),
.Y(n_238)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_216),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_169),
.B1(n_172),
.B2(n_171),
.Y(n_211)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_215),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_186),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_223),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_160),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_144),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_122),
.C(n_73),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_225),
.C(n_198),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_89),
.B1(n_97),
.B2(n_100),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_222),
.Y(n_241)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_203),
.A2(n_89),
.B1(n_97),
.B2(n_60),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_60),
.C(n_97),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_197),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_21),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_208),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_224),
.A2(n_204),
.B1(n_200),
.B2(n_196),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_232),
.A2(n_243),
.B1(n_246),
.B2(n_0),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_216),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_218),
.Y(n_248)
);

A2O1A1O1Ixp25_ASAP7_75t_L g234 ( 
.A1(n_226),
.A2(n_184),
.B(n_182),
.C(n_194),
.D(n_201),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_234),
.B(n_21),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_21),
.C(n_1),
.Y(n_256)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_220),
.A2(n_191),
.B1(n_199),
.B2(n_180),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_187),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_0),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_181),
.B1(n_192),
.B2(n_189),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_252),
.Y(n_262)
);

XNOR2x1_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_215),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_231),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_250),
.A2(n_260),
.B(n_247),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_225),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_217),
.B1(n_210),
.B2(n_213),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_257),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_236),
.A2(n_227),
.B(n_223),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_258),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_241),
.C(n_230),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_7),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_237),
.Y(n_271)
);

OAI31xp33_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_6),
.A3(n_13),
.B(n_2),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_243),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_239),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_266),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_270),
.B(n_272),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_269),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_238),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_230),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

INVxp33_ASAP7_75t_SL g274 ( 
.A(n_267),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_274),
.A2(n_281),
.B(n_4),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_264),
.A2(n_261),
.B1(n_229),
.B2(n_240),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_280),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_254),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_5),
.Y(n_285)
);

AO21x1_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_256),
.B(n_254),
.Y(n_280)
);

OAI21x1_ASAP7_75t_SL g281 ( 
.A1(n_272),
.A2(n_8),
.B(n_3),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_278),
.A2(n_262),
.B(n_1),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_9),
.C(n_11),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_277),
.A2(n_3),
.B(n_4),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_283),
.A2(n_285),
.B(n_9),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_287),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_L g286 ( 
.A1(n_277),
.A2(n_6),
.B(n_8),
.Y(n_286)
);

AOI21x1_ASAP7_75t_L g289 ( 
.A1(n_286),
.A2(n_9),
.B(n_11),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_8),
.Y(n_287)
);

AOI221xp5_ASAP7_75t_SL g295 ( 
.A1(n_289),
.A2(n_291),
.B1(n_12),
.B2(n_13),
.C(n_16),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_288),
.A2(n_279),
.B1(n_11),
.B2(n_12),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_12),
.C(n_13),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_16),
.C(n_292),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_294),
.A2(n_295),
.B(n_296),
.Y(n_297)
);

XNOR2x2_ASAP7_75t_SL g298 ( 
.A(n_297),
.B(n_16),
.Y(n_298)
);


endmodule