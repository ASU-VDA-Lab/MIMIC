module fake_ariane_180_n_1292 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_345, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_221, n_321, n_86, n_361, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_359, n_155, n_127, n_1292);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_345;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_359;
input n_155;
input n_127;

output n_1292;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_868;
wire n_884;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_365;
wire n_1013;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1230;
wire n_612;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_461;
wire n_1121;
wire n_490;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_444;
wire n_851;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_1178;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_746;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_965;
wire n_934;
wire n_1220;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_776;
wire n_424;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1134;
wire n_647;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_845;
wire n_888;
wire n_551;
wire n_417;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1266;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1243;
wire n_608;
wire n_1037;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_1204;
wire n_994;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_1057;
wire n_1011;
wire n_978;
wire n_828;
wire n_558;
wire n_653;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_679;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_997;
wire n_635;
wire n_694;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1148;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_371;
wire n_1114;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_895;
wire n_583;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_548;
wire n_523;
wire n_457;
wire n_782;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_153),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_227),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_19),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_14),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_253),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_131),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_180),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_150),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_247),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_198),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_310),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_15),
.Y(n_376)
);

BUFx10_ASAP7_75t_L g377 ( 
.A(n_240),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_157),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_162),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_66),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_279),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_202),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_68),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_278),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_119),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_132),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_158),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_141),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_294),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_126),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_223),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_98),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_348),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_103),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_134),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_89),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_333),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_261),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_260),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_332),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_315),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_356),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_49),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_118),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_358),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_273),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_283),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_228),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_274),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_231),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_179),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_205),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_133),
.Y(n_414)
);

BUFx5_ASAP7_75t_L g415 ( 
.A(n_1),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_308),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_200),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_284),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_208),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_363),
.Y(n_420)
);

BUFx10_ASAP7_75t_L g421 ( 
.A(n_112),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_282),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_15),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_77),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_187),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_182),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_258),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_144),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_85),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_276),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_136),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_335),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_189),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_297),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_347),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_212),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_111),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_129),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_192),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_31),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_147),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_113),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_17),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_222),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_287),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_52),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_152),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_103),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_4),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_277),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_306),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_351),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_203),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_201),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_164),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_56),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_300),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_216),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_262),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_211),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_196),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_83),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_121),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_171),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_142),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_185),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_204),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_352),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_361),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_81),
.Y(n_470)
);

BUFx10_ASAP7_75t_L g471 ( 
.A(n_165),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_281),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g473 ( 
.A(n_298),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_174),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_143),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_345),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_52),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_219),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_17),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_115),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_275),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_346),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_357),
.Y(n_483)
);

NOR2xp67_ASAP7_75t_L g484 ( 
.A(n_194),
.B(n_176),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_210),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_69),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_175),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_123),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_183),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_326),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_138),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_159),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_265),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_236),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_266),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_72),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_256),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_209),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_13),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_26),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_106),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_109),
.Y(n_502)
);

BUFx10_ASAP7_75t_L g503 ( 
.A(n_327),
.Y(n_503)
);

BUFx10_ASAP7_75t_L g504 ( 
.A(n_197),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_50),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_69),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_76),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_148),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_214),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_12),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_244),
.Y(n_511)
);

BUFx10_ASAP7_75t_L g512 ( 
.A(n_321),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_181),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_97),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_84),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_49),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_93),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_130),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_43),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_289),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_226),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_225),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_122),
.Y(n_523)
);

NOR2xp67_ASAP7_75t_L g524 ( 
.A(n_304),
.B(n_213),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_268),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_167),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_229),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_13),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_169),
.B(n_269),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_245),
.Y(n_530)
);

BUFx10_ASAP7_75t_L g531 ( 
.A(n_292),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_376),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_456),
.B(n_0),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_415),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_369),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_415),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_415),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_376),
.B(n_2),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_409),
.Y(n_539)
);

BUFx8_ASAP7_75t_L g540 ( 
.A(n_403),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_474),
.B(n_415),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_409),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_384),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_384),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_391),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_444),
.A2(n_482),
.B(n_475),
.Y(n_546)
);

OAI21x1_ASAP7_75t_L g547 ( 
.A1(n_444),
.A2(n_116),
.B(n_114),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_409),
.Y(n_548)
);

BUFx12f_ASAP7_75t_L g549 ( 
.A(n_377),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_386),
.Y(n_550)
);

INVx5_ASAP7_75t_L g551 ( 
.A(n_409),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_528),
.B(n_487),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_475),
.A2(n_120),
.B(n_117),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_486),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_419),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_419),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_419),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_415),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_415),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_497),
.B(n_375),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_386),
.Y(n_561)
);

INVx5_ASAP7_75t_L g562 ( 
.A(n_377),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_379),
.B(n_7),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_368),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_365),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_394),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_421),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_394),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_412),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_412),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_480),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_380),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g573 ( 
.A1(n_482),
.A2(n_125),
.B(n_124),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_480),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_381),
.B(n_8),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_370),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_393),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_385),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_387),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_366),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_397),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_499),
.B(n_8),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_429),
.Y(n_583)
);

OAI21x1_ASAP7_75t_L g584 ( 
.A1(n_389),
.A2(n_128),
.B(n_127),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_499),
.B(n_9),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_396),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_367),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_390),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_402),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_373),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_383),
.B(n_9),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_411),
.B(n_10),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_372),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_440),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_443),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_413),
.Y(n_596)
);

OAI22x1_ASAP7_75t_R g597 ( 
.A1(n_437),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_374),
.B(n_11),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_431),
.Y(n_599)
);

AND2x6_ASAP7_75t_L g600 ( 
.A(n_422),
.B(n_426),
.Y(n_600)
);

OA21x2_ASAP7_75t_L g601 ( 
.A1(n_433),
.A2(n_16),
.B(n_18),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_460),
.A2(n_19),
.B1(n_16),
.B2(n_18),
.Y(n_602)
);

INVx6_ASAP7_75t_L g603 ( 
.A(n_531),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_479),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_496),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_539),
.Y(n_606)
);

BUFx10_ASAP7_75t_L g607 ( 
.A(n_593),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_603),
.Y(n_608)
);

AOI21x1_ASAP7_75t_L g609 ( 
.A1(n_558),
.A2(n_441),
.B(n_435),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_539),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_564),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_539),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_539),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_598),
.B(n_521),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_572),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_562),
.B(n_400),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_562),
.B(n_509),
.Y(n_617)
);

INVxp33_ASAP7_75t_SL g618 ( 
.A(n_593),
.Y(n_618)
);

AND3x2_ASAP7_75t_L g619 ( 
.A(n_552),
.B(n_513),
.C(n_502),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_542),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_542),
.Y(n_621)
);

CKINVDCx6p67_ASAP7_75t_R g622 ( 
.A(n_549),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_542),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_548),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_548),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_L g626 ( 
.A(n_600),
.B(n_371),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_577),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_565),
.B(n_498),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_576),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_600),
.B(n_527),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_567),
.B(n_560),
.Y(n_631)
);

INVxp67_ASAP7_75t_SL g632 ( 
.A(n_541),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_549),
.B(n_421),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_576),
.Y(n_634)
);

INVx5_ASAP7_75t_L g635 ( 
.A(n_551),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_587),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_L g637 ( 
.A(n_600),
.B(n_541),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_580),
.B(n_498),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_603),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_581),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_534),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_576),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_583),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_590),
.B(n_473),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_555),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_594),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_534),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_632),
.B(n_603),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_611),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_615),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_641),
.B(n_536),
.Y(n_651)
);

A2O1A1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_637),
.A2(n_585),
.B(n_575),
.C(n_563),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_627),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_608),
.B(n_590),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_608),
.B(n_543),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_640),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_616),
.B(n_543),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_643),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_644),
.B(n_544),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_646),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_628),
.B(n_544),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_638),
.B(n_550),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_617),
.B(n_550),
.Y(n_663)
);

BUFx5_ASAP7_75t_L g664 ( 
.A(n_641),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_647),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_639),
.B(n_533),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_636),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_629),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_629),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_647),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_631),
.A2(n_535),
.B1(n_602),
.B2(n_545),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_639),
.B(n_570),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_637),
.B(n_536),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_634),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_634),
.B(n_537),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_618),
.B(n_538),
.Y(n_676)
);

AO221x1_ASAP7_75t_L g677 ( 
.A1(n_636),
.A2(n_423),
.B1(n_597),
.B2(n_507),
.C(n_506),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_607),
.B(n_585),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_619),
.B(n_575),
.C(n_563),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_626),
.A2(n_585),
.B1(n_591),
.B2(n_582),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_642),
.B(n_566),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_642),
.B(n_568),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_642),
.B(n_568),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_626),
.B(n_586),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_607),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_622),
.B(n_532),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_609),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_630),
.B(n_561),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_609),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_614),
.B(n_591),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_606),
.Y(n_691)
);

NOR2xp67_ASAP7_75t_L g692 ( 
.A(n_633),
.B(n_578),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_645),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_610),
.B(n_537),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_621),
.B(n_592),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_612),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_613),
.B(n_559),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_620),
.Y(n_698)
);

OAI22xp33_ASAP7_75t_L g699 ( 
.A1(n_620),
.A2(n_505),
.B1(n_449),
.B2(n_477),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_623),
.B(n_578),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_635),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_623),
.B(n_546),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_624),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_625),
.B(n_579),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_673),
.A2(n_513),
.B(n_553),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_673),
.A2(n_573),
.B(n_547),
.Y(n_706)
);

BUFx8_ASAP7_75t_L g707 ( 
.A(n_685),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_648),
.B(n_540),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_652),
.A2(n_584),
.B(n_529),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_659),
.A2(n_601),
.B(n_625),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_657),
.B(n_589),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_661),
.B(n_589),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_655),
.Y(n_713)
);

O2A1O1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_649),
.A2(n_500),
.B(n_516),
.C(n_510),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_662),
.B(n_596),
.Y(n_715)
);

OAI21xp5_ASAP7_75t_L g716 ( 
.A1(n_702),
.A2(n_447),
.B(n_442),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_663),
.B(n_680),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_695),
.A2(n_651),
.B(n_675),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_650),
.B(n_653),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_656),
.B(n_596),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_664),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_671),
.A2(n_473),
.B1(n_514),
.B2(n_404),
.Y(n_722)
);

O2A1O1Ixp5_ASAP7_75t_L g723 ( 
.A1(n_665),
.A2(n_451),
.B(n_454),
.C(n_450),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_658),
.B(n_576),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_660),
.B(n_588),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_670),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_681),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_668),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_676),
.B(n_515),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_672),
.B(n_395),
.Y(n_730)
);

OR2x6_ASAP7_75t_L g731 ( 
.A(n_690),
.B(n_595),
.Y(n_731)
);

NOR3xp33_ASAP7_75t_L g732 ( 
.A(n_678),
.B(n_519),
.C(n_517),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_669),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_687),
.A2(n_464),
.B(n_457),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_689),
.A2(n_469),
.B(n_466),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_666),
.A2(n_476),
.B(n_472),
.Y(n_736)
);

A2O1A1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_679),
.A2(n_485),
.B(n_489),
.C(n_478),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_692),
.B(n_424),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_674),
.A2(n_493),
.B(n_492),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_682),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_664),
.B(n_599),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_686),
.B(n_554),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_654),
.A2(n_448),
.B1(n_462),
.B2(n_446),
.Y(n_743)
);

OAI21xp33_ASAP7_75t_L g744 ( 
.A1(n_683),
.A2(n_501),
.B(n_470),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_684),
.B(n_406),
.Y(n_745)
);

AO21x1_ASAP7_75t_L g746 ( 
.A1(n_688),
.A2(n_511),
.B(n_508),
.Y(n_746)
);

AOI21x1_ASAP7_75t_L g747 ( 
.A1(n_694),
.A2(n_524),
.B(n_484),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_700),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_699),
.A2(n_599),
.B1(n_569),
.B2(n_571),
.Y(n_749)
);

NOR2xp67_ASAP7_75t_L g750 ( 
.A(n_693),
.B(n_604),
.Y(n_750)
);

AND2x6_ASAP7_75t_SL g751 ( 
.A(n_677),
.B(n_605),
.Y(n_751)
);

BUFx12f_ASAP7_75t_L g752 ( 
.A(n_698),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_704),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_691),
.B(n_471),
.Y(n_754)
);

AO21x1_ASAP7_75t_L g755 ( 
.A1(n_697),
.A2(n_523),
.B(n_520),
.Y(n_755)
);

NAND3xp33_ASAP7_75t_L g756 ( 
.A(n_696),
.B(n_569),
.C(n_561),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_703),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_701),
.A2(n_430),
.B1(n_467),
.B2(n_425),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_701),
.A2(n_635),
.B(n_551),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_648),
.B(n_561),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_648),
.B(n_569),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_665),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_685),
.B(n_569),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_673),
.A2(n_382),
.B(n_378),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_673),
.A2(n_392),
.B(n_388),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_648),
.B(n_571),
.Y(n_766)
);

O2A1O1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_652),
.A2(n_518),
.B(n_468),
.C(n_21),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_667),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_648),
.B(n_471),
.Y(n_769)
);

OAI21xp5_ASAP7_75t_L g770 ( 
.A1(n_673),
.A2(n_399),
.B(n_398),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_673),
.A2(n_405),
.B(n_401),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_648),
.B(n_571),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_652),
.A2(n_574),
.B(n_408),
.C(n_410),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_673),
.A2(n_414),
.B(n_407),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_673),
.A2(n_417),
.B(n_416),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_673),
.A2(n_420),
.B(n_418),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_665),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_667),
.B(n_574),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_673),
.A2(n_428),
.B(n_427),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_648),
.B(n_503),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_648),
.B(n_574),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_673),
.A2(n_434),
.B(n_432),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_648),
.B(n_436),
.Y(n_783)
);

OAI21x1_ASAP7_75t_L g784 ( 
.A1(n_687),
.A2(n_504),
.B(n_503),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_680),
.A2(n_439),
.B1(n_445),
.B2(n_438),
.Y(n_785)
);

AND2x6_ASAP7_75t_L g786 ( 
.A(n_673),
.B(n_555),
.Y(n_786)
);

AOI21x1_ASAP7_75t_L g787 ( 
.A1(n_673),
.A2(n_621),
.B(n_556),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_648),
.B(n_452),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_648),
.B(n_504),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_673),
.A2(n_455),
.B(n_453),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_668),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_769),
.B(n_512),
.Y(n_792)
);

AO31x2_ASAP7_75t_L g793 ( 
.A1(n_755),
.A2(n_512),
.A3(n_556),
.B(n_555),
.Y(n_793)
);

OA22x2_ASAP7_75t_L g794 ( 
.A1(n_722),
.A2(n_459),
.B1(n_461),
.B2(n_458),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_731),
.B(n_20),
.Y(n_795)
);

AOI221x1_ASAP7_75t_L g796 ( 
.A1(n_709),
.A2(n_621),
.B1(n_557),
.B2(n_556),
.C(n_555),
.Y(n_796)
);

BUFx12f_ASAP7_75t_L g797 ( 
.A(n_707),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_752),
.Y(n_798)
);

NAND3xp33_ASAP7_75t_L g799 ( 
.A(n_780),
.B(n_465),
.C(n_463),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_768),
.Y(n_800)
);

AO22x2_ASAP7_75t_L g801 ( 
.A1(n_762),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_791),
.Y(n_802)
);

OA21x2_ASAP7_75t_L g803 ( 
.A1(n_710),
.A2(n_483),
.B(n_481),
.Y(n_803)
);

AO21x2_ASAP7_75t_L g804 ( 
.A1(n_716),
.A2(n_557),
.B(n_556),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_707),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_708),
.B(n_748),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_753),
.B(n_488),
.Y(n_807)
);

AOI21xp33_ASAP7_75t_L g808 ( 
.A1(n_729),
.A2(n_491),
.B(n_490),
.Y(n_808)
);

AOI21x1_ASAP7_75t_L g809 ( 
.A1(n_787),
.A2(n_621),
.B(n_557),
.Y(n_809)
);

OAI21xp33_ASAP7_75t_L g810 ( 
.A1(n_770),
.A2(n_495),
.B(n_494),
.Y(n_810)
);

AOI221xp5_ASAP7_75t_SL g811 ( 
.A1(n_719),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.C(n_25),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_763),
.B(n_522),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_734),
.A2(n_735),
.B(n_771),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_783),
.B(n_525),
.Y(n_814)
);

OAI21xp33_ASAP7_75t_L g815 ( 
.A1(n_782),
.A2(n_530),
.B(n_526),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_777),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_727),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_745),
.B(n_23),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_724),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_791),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_778),
.B(n_25),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_712),
.B(n_26),
.Y(n_822)
);

AO31x2_ASAP7_75t_L g823 ( 
.A1(n_746),
.A2(n_29),
.A3(n_27),
.B(n_28),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_773),
.A2(n_137),
.B(n_135),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_715),
.B(n_28),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_740),
.A2(n_140),
.B(n_139),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_731),
.B(n_30),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_741),
.A2(n_146),
.B(n_145),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_788),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_731),
.Y(n_830)
);

AOI21xp33_ASAP7_75t_L g831 ( 
.A1(n_717),
.A2(n_32),
.B(n_33),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_711),
.B(n_750),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_764),
.A2(n_151),
.B(n_149),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_791),
.Y(n_834)
);

NAND2x1_ASAP7_75t_L g835 ( 
.A(n_728),
.B(n_154),
.Y(n_835)
);

OA21x2_ASAP7_75t_L g836 ( 
.A1(n_784),
.A2(n_156),
.B(n_155),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_720),
.B(n_34),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_R g838 ( 
.A(n_747),
.B(n_160),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_767),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_728),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_789),
.B(n_35),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_732),
.B(n_36),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_757),
.B(n_37),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_725),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_765),
.A2(n_163),
.B(n_161),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_737),
.B(n_38),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_L g847 ( 
.A(n_785),
.B(n_39),
.C(n_40),
.Y(n_847)
);

O2A1O1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_714),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_774),
.A2(n_168),
.B(n_166),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_775),
.A2(n_172),
.B(n_170),
.Y(n_850)
);

NOR2xp67_ASAP7_75t_L g851 ( 
.A(n_758),
.B(n_173),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_776),
.A2(n_178),
.B(n_177),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_760),
.B(n_41),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_730),
.B(n_42),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_733),
.Y(n_855)
);

BUFx10_ASAP7_75t_L g856 ( 
.A(n_751),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_761),
.B(n_43),
.Y(n_857)
);

OAI21xp33_ASAP7_75t_L g858 ( 
.A1(n_744),
.A2(n_44),
.B(n_45),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_766),
.B(n_44),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_779),
.A2(n_186),
.B(n_184),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_790),
.A2(n_723),
.B(n_739),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_772),
.B(n_46),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_781),
.B(n_47),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_738),
.A2(n_190),
.B(n_188),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_786),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_736),
.A2(n_193),
.B(n_191),
.Y(n_866)
);

BUFx4f_ASAP7_75t_L g867 ( 
.A(n_786),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_786),
.A2(n_199),
.B(n_195),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_SL g869 ( 
.A(n_743),
.B(n_47),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_754),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_749),
.B(n_48),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_756),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_872)
);

INVx4_ASAP7_75t_L g873 ( 
.A(n_759),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_769),
.B(n_53),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_769),
.B(n_54),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_705),
.A2(n_207),
.B(n_206),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_726),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_769),
.B(n_55),
.Y(n_878)
);

NAND3xp33_ASAP7_75t_L g879 ( 
.A(n_769),
.B(n_55),
.C(n_56),
.Y(n_879)
);

OAI22x1_ASAP7_75t_L g880 ( 
.A1(n_722),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_880)
);

OAI21xp5_ASAP7_75t_L g881 ( 
.A1(n_705),
.A2(n_217),
.B(n_215),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_752),
.Y(n_882)
);

NAND2x1p5_ASAP7_75t_L g883 ( 
.A(n_713),
.B(n_57),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_726),
.Y(n_884)
);

AOI21x1_ASAP7_75t_L g885 ( 
.A1(n_706),
.A2(n_220),
.B(n_218),
.Y(n_885)
);

AND2x2_ASAP7_75t_SL g886 ( 
.A(n_708),
.B(n_58),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_708),
.B(n_59),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_716),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_768),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_705),
.A2(n_224),
.B(n_221),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_769),
.B(n_60),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_769),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_769),
.B(n_64),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_726),
.Y(n_894)
);

NOR2x1_ASAP7_75t_SL g895 ( 
.A(n_721),
.B(n_230),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_718),
.A2(n_233),
.B(n_232),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_769),
.B(n_65),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_791),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_731),
.B(n_66),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_718),
.A2(n_235),
.B(n_234),
.Y(n_900)
);

AOI22x1_ASAP7_75t_L g901 ( 
.A1(n_709),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_769),
.B(n_67),
.Y(n_902)
);

OAI21x1_ASAP7_75t_L g903 ( 
.A1(n_706),
.A2(n_238),
.B(n_237),
.Y(n_903)
);

OAI21x1_ASAP7_75t_L g904 ( 
.A1(n_706),
.A2(n_241),
.B(n_239),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_713),
.B(n_71),
.Y(n_905)
);

INVx4_ASAP7_75t_L g906 ( 
.A(n_752),
.Y(n_906)
);

INVxp67_ASAP7_75t_SL g907 ( 
.A(n_768),
.Y(n_907)
);

OAI21x1_ASAP7_75t_L g908 ( 
.A1(n_706),
.A2(n_243),
.B(n_242),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_718),
.A2(n_248),
.B(n_246),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_769),
.B(n_71),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_718),
.A2(n_250),
.B(n_249),
.Y(n_911)
);

OAI21x1_ASAP7_75t_L g912 ( 
.A1(n_706),
.A2(n_252),
.B(n_251),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_769),
.B(n_72),
.Y(n_913)
);

OAI21x1_ASAP7_75t_L g914 ( 
.A1(n_706),
.A2(n_255),
.B(n_254),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_716),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_915)
);

OR2x6_ASAP7_75t_L g916 ( 
.A(n_906),
.B(n_73),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_802),
.Y(n_917)
);

OA21x2_ASAP7_75t_L g918 ( 
.A1(n_796),
.A2(n_259),
.B(n_257),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_886),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_800),
.Y(n_920)
);

OAI211xp5_ASAP7_75t_L g921 ( 
.A1(n_887),
.A2(n_78),
.B(n_79),
.C(n_80),
.Y(n_921)
);

NAND2x1p5_ASAP7_75t_L g922 ( 
.A(n_798),
.B(n_263),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_813),
.A2(n_78),
.B(n_79),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_889),
.B(n_80),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_806),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_925)
);

BUFx4f_ASAP7_75t_L g926 ( 
.A(n_797),
.Y(n_926)
);

NAND2x1p5_ASAP7_75t_L g927 ( 
.A(n_882),
.B(n_264),
.Y(n_927)
);

BUFx8_ASAP7_75t_L g928 ( 
.A(n_795),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_906),
.Y(n_929)
);

OA21x2_ASAP7_75t_L g930 ( 
.A1(n_876),
.A2(n_302),
.B(n_362),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_869),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_805),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_817),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_830),
.B(n_86),
.Y(n_934)
);

OA21x2_ASAP7_75t_L g935 ( 
.A1(n_881),
.A2(n_303),
.B(n_360),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_856),
.Y(n_936)
);

AOI221xp5_ASAP7_75t_L g937 ( 
.A1(n_880),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.C(n_90),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_907),
.B(n_88),
.Y(n_938)
);

NAND2x1p5_ASAP7_75t_L g939 ( 
.A(n_867),
.B(n_267),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_867),
.B(n_270),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_795),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_817),
.Y(n_942)
);

AOI21x1_ASAP7_75t_L g943 ( 
.A1(n_803),
.A2(n_305),
.B(n_359),
.Y(n_943)
);

BUFx2_ASAP7_75t_SL g944 ( 
.A(n_865),
.Y(n_944)
);

INVx6_ASAP7_75t_L g945 ( 
.A(n_856),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_899),
.B(n_91),
.Y(n_946)
);

OAI21x1_ASAP7_75t_L g947 ( 
.A1(n_903),
.A2(n_307),
.B(n_355),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_816),
.Y(n_948)
);

OAI21x1_ASAP7_75t_SL g949 ( 
.A1(n_895),
.A2(n_92),
.B(n_94),
.Y(n_949)
);

AOI21x1_ASAP7_75t_L g950 ( 
.A1(n_803),
.A2(n_301),
.B(n_354),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_904),
.A2(n_912),
.B(n_908),
.Y(n_951)
);

AOI221xp5_ASAP7_75t_L g952 ( 
.A1(n_915),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.C(n_97),
.Y(n_952)
);

INVx5_ASAP7_75t_L g953 ( 
.A(n_865),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_877),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_899),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_884),
.B(n_96),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_914),
.A2(n_309),
.B(n_353),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_894),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_827),
.B(n_99),
.Y(n_959)
);

OA21x2_ASAP7_75t_L g960 ( 
.A1(n_890),
.A2(n_824),
.B(n_826),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_814),
.A2(n_299),
.B(n_350),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_792),
.B(n_100),
.Y(n_962)
);

AO21x2_ASAP7_75t_L g963 ( 
.A1(n_861),
.A2(n_296),
.B(n_349),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_802),
.Y(n_964)
);

AOI221xp5_ASAP7_75t_L g965 ( 
.A1(n_842),
.A2(n_101),
.B1(n_102),
.B2(n_104),
.C(n_105),
.Y(n_965)
);

AOI21xp33_ASAP7_75t_SL g966 ( 
.A1(n_874),
.A2(n_101),
.B(n_102),
.Y(n_966)
);

NAND3xp33_ASAP7_75t_L g967 ( 
.A(n_892),
.B(n_104),
.C(n_105),
.Y(n_967)
);

INVx5_ASAP7_75t_L g968 ( 
.A(n_802),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_853),
.A2(n_312),
.B(n_344),
.Y(n_969)
);

OAI21x1_ASAP7_75t_L g970 ( 
.A1(n_885),
.A2(n_311),
.B(n_342),
.Y(n_970)
);

BUFx4f_ASAP7_75t_L g971 ( 
.A(n_854),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_840),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_875),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_820),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_840),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_855),
.Y(n_976)
);

OAI221xp5_ASAP7_75t_L g977 ( 
.A1(n_854),
.A2(n_110),
.B1(n_111),
.B2(n_271),
.C(n_272),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_821),
.B(n_364),
.Y(n_978)
);

AO21x2_ASAP7_75t_L g979 ( 
.A1(n_849),
.A2(n_850),
.B(n_804),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_820),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_834),
.B(n_280),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_794),
.A2(n_285),
.B1(n_286),
.B2(n_288),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_883),
.B(n_290),
.Y(n_983)
);

AO21x2_ASAP7_75t_L g984 ( 
.A1(n_868),
.A2(n_291),
.B(n_293),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_905),
.B(n_341),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_896),
.A2(n_295),
.B(n_313),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_822),
.A2(n_314),
.B(n_316),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_857),
.A2(n_317),
.B(n_318),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_832),
.B(n_319),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_843),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_L g991 ( 
.A(n_878),
.B(n_320),
.C(n_322),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_891),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_870),
.B(n_328),
.Y(n_993)
);

INVxp67_ASAP7_75t_SL g994 ( 
.A(n_898),
.Y(n_994)
);

AO22x2_ASAP7_75t_L g995 ( 
.A1(n_893),
.A2(n_329),
.B1(n_330),
.B2(n_331),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_SL g996 ( 
.A1(n_897),
.A2(n_334),
.B(n_336),
.C(n_337),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_SL g997 ( 
.A1(n_902),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.Y(n_997)
);

OR2x6_ASAP7_75t_L g998 ( 
.A(n_851),
.B(n_801),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_900),
.A2(n_911),
.B(n_909),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_838),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_835),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_807),
.B(n_913),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_841),
.Y(n_1003)
);

AOI221xp5_ASAP7_75t_L g1004 ( 
.A1(n_831),
.A2(n_858),
.B1(n_808),
.B2(n_848),
.C(n_910),
.Y(n_1004)
);

AOI22x1_ASAP7_75t_L g1005 ( 
.A1(n_833),
.A2(n_845),
.B1(n_852),
.B2(n_860),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_871),
.Y(n_1006)
);

OAI22x1_ASAP7_75t_L g1007 ( 
.A1(n_879),
.A2(n_901),
.B1(n_818),
.B2(n_847),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_810),
.A2(n_815),
.B1(n_812),
.B2(n_846),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_811),
.B(n_888),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_799),
.A2(n_825),
.B1(n_837),
.B2(n_839),
.Y(n_1010)
);

AOI21x1_ASAP7_75t_L g1011 ( 
.A1(n_862),
.A2(n_863),
.B(n_836),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_828),
.A2(n_844),
.B(n_819),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_866),
.A2(n_859),
.B(n_864),
.C(n_829),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_SL g1014 ( 
.A1(n_872),
.A2(n_895),
.B(n_873),
.C(n_823),
.Y(n_1014)
);

NAND2xp33_ASAP7_75t_SL g1015 ( 
.A(n_823),
.B(n_793),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_823),
.A2(n_886),
.B1(n_887),
.B2(n_869),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_806),
.A2(n_875),
.B1(n_878),
.B2(n_874),
.Y(n_1017)
);

OA21x2_ASAP7_75t_L g1018 ( 
.A1(n_796),
.A2(n_881),
.B(n_876),
.Y(n_1018)
);

OAI221xp5_ASAP7_75t_L g1019 ( 
.A1(n_887),
.A2(n_729),
.B1(n_671),
.B2(n_806),
.C(n_667),
.Y(n_1019)
);

NAND2x1p5_ASAP7_75t_L g1020 ( 
.A(n_798),
.B(n_882),
.Y(n_1020)
);

NAND3xp33_ASAP7_75t_L g1021 ( 
.A(n_887),
.B(n_869),
.C(n_780),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_817),
.Y(n_1022)
);

INVxp33_ASAP7_75t_L g1023 ( 
.A(n_800),
.Y(n_1023)
);

OR2x6_ASAP7_75t_L g1024 ( 
.A(n_906),
.B(n_798),
.Y(n_1024)
);

OAI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_806),
.A2(n_869),
.B1(n_887),
.B2(n_614),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_886),
.B(n_742),
.Y(n_1026)
);

OA21x2_ASAP7_75t_L g1027 ( 
.A1(n_796),
.A2(n_881),
.B(n_876),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_806),
.A2(n_875),
.B1(n_878),
.B2(n_874),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_797),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_SL g1030 ( 
.A(n_798),
.Y(n_1030)
);

INVx6_ASAP7_75t_L g1031 ( 
.A(n_797),
.Y(n_1031)
);

NAND2x1p5_ASAP7_75t_L g1032 ( 
.A(n_798),
.B(n_882),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_805),
.Y(n_1033)
);

AOI21x1_ASAP7_75t_L g1034 ( 
.A1(n_796),
.A2(n_809),
.B(n_803),
.Y(n_1034)
);

BUFx12f_ASAP7_75t_L g1035 ( 
.A(n_1029),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_958),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1026),
.B(n_941),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_933),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_948),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_1019),
.B(n_1025),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_924),
.B(n_955),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_948),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_920),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_1003),
.A2(n_1021),
.B1(n_1016),
.B2(n_962),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_954),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_998),
.A2(n_1016),
.B1(n_971),
.B2(n_919),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_1023),
.B(n_1002),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_946),
.B(n_934),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_942),
.B(n_1022),
.Y(n_1049)
);

INVxp67_ASAP7_75t_L g1050 ( 
.A(n_1006),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_990),
.B(n_1017),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_1033),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_956),
.Y(n_1053)
);

BUFx2_ASAP7_75t_SL g1054 ( 
.A(n_1030),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_972),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_975),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_926),
.Y(n_1057)
);

AOI21xp33_ASAP7_75t_L g1058 ( 
.A1(n_1028),
.A2(n_1007),
.B(n_1004),
.Y(n_1058)
);

NOR2x1_ASAP7_75t_SL g1059 ( 
.A(n_944),
.B(n_953),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_938),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_923),
.A2(n_1013),
.B(n_1009),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_934),
.B(n_959),
.Y(n_1062)
);

NOR2x1_ASAP7_75t_L g1063 ( 
.A(n_980),
.B(n_964),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_931),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_976),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_932),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_931),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_981),
.Y(n_1068)
);

INVxp67_ASAP7_75t_L g1069 ( 
.A(n_994),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_925),
.Y(n_1070)
);

AOI21x1_ASAP7_75t_L g1071 ( 
.A1(n_1034),
.A2(n_1011),
.B(n_950),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_928),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_937),
.A2(n_952),
.B1(n_967),
.B2(n_965),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_916),
.B(n_1000),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_917),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_936),
.B(n_945),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1010),
.A2(n_960),
.B(n_1012),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_951),
.A2(n_999),
.B(n_1005),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1008),
.B(n_978),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_974),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_926),
.Y(n_1081)
);

OA21x2_ASAP7_75t_L g1082 ( 
.A1(n_943),
.A2(n_950),
.B(n_1005),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_1030),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_945),
.B(n_983),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_973),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_993),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_964),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_997),
.A2(n_977),
.B1(n_1024),
.B2(n_929),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_968),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_985),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_1024),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_SL g1092 ( 
.A1(n_997),
.A2(n_995),
.B1(n_921),
.B2(n_935),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_1032),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_1020),
.B(n_927),
.Y(n_1094)
);

OAI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_966),
.A2(n_992),
.B1(n_987),
.B2(n_922),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_1031),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_966),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_939),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1031),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_995),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_982),
.B(n_940),
.Y(n_1101)
);

AOI211xp5_ASAP7_75t_L g1102 ( 
.A1(n_1014),
.A2(n_996),
.B(n_992),
.C(n_991),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_949),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_989),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1015),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_963),
.B(n_984),
.Y(n_1106)
);

BUFx2_ASAP7_75t_SL g1107 ( 
.A(n_1001),
.Y(n_1107)
);

INVxp67_ASAP7_75t_L g1108 ( 
.A(n_961),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1018),
.A2(n_1027),
.B(n_988),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_1001),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_918),
.B(n_930),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_979),
.Y(n_1112)
);

OAI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_930),
.A2(n_935),
.B1(n_918),
.B2(n_969),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_943),
.A2(n_986),
.B1(n_947),
.B2(n_957),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1036),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1068),
.B(n_970),
.Y(n_1116)
);

OAI31xp33_ASAP7_75t_SL g1117 ( 
.A1(n_1095),
.A2(n_1040),
.A3(n_1051),
.B(n_1061),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_1052),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1086),
.A2(n_1044),
.B1(n_1073),
.B2(n_1040),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1039),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1042),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1098),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_1043),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_1043),
.Y(n_1124)
);

BUFx2_ASAP7_75t_SL g1125 ( 
.A(n_1052),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1037),
.B(n_1062),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_1086),
.B(n_1051),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_1064),
.B(n_1067),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1045),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1048),
.B(n_1041),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1049),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1049),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1047),
.B(n_1060),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1050),
.B(n_1084),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1038),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_1091),
.Y(n_1136)
);

BUFx12f_ASAP7_75t_L g1137 ( 
.A(n_1081),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_1105),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_1093),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_1050),
.B(n_1053),
.Y(n_1140)
);

AO21x2_ASAP7_75t_L g1141 ( 
.A1(n_1113),
.A2(n_1071),
.B(n_1109),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1100),
.B(n_1058),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1055),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1112),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1056),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1058),
.B(n_1061),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_1112),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1074),
.B(n_1090),
.Y(n_1148)
);

NOR2x1p5_ASAP7_75t_L g1149 ( 
.A(n_1081),
.B(n_1099),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1076),
.B(n_1065),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1046),
.B(n_1054),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1088),
.B(n_1097),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1104),
.B(n_1085),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1099),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1079),
.B(n_1070),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_SL g1156 ( 
.A(n_1066),
.B(n_1096),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1094),
.B(n_1096),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1083),
.B(n_1089),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1083),
.B(n_1080),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1073),
.B(n_1069),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_1066),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1075),
.Y(n_1162)
);

AND2x4_ASAP7_75t_SL g1163 ( 
.A(n_1098),
.B(n_1072),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_1057),
.Y(n_1164)
);

AND2x4_ASAP7_75t_SL g1165 ( 
.A(n_1098),
.B(n_1072),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1077),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1092),
.B(n_1103),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1087),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1101),
.B(n_1111),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_1138),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1120),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1121),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1140),
.B(n_1153),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1129),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1129),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1127),
.B(n_1095),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1169),
.B(n_1106),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1116),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1127),
.B(n_1110),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_1123),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1136),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1128),
.B(n_1063),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_1135),
.Y(n_1183)
);

AND2x2_ASAP7_75t_SL g1184 ( 
.A(n_1117),
.B(n_1082),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1115),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1128),
.B(n_1107),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1119),
.A2(n_1113),
.B1(n_1108),
.B2(n_1035),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1167),
.B(n_1082),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1138),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1133),
.B(n_1059),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1167),
.B(n_1078),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1131),
.B(n_1102),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1132),
.B(n_1102),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1143),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1145),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1146),
.B(n_1108),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1116),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1139),
.Y(n_1198)
);

INVxp67_ASAP7_75t_SL g1199 ( 
.A(n_1144),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1183),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1192),
.B(n_1155),
.Y(n_1201)
);

OR2x2_ASAP7_75t_L g1202 ( 
.A(n_1196),
.B(n_1144),
.Y(n_1202)
);

OR2x2_ASAP7_75t_L g1203 ( 
.A(n_1196),
.B(n_1147),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1192),
.B(n_1142),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1171),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1172),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1189),
.B(n_1147),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1188),
.B(n_1166),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1174),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1170),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1177),
.B(n_1191),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1193),
.B(n_1142),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1193),
.B(n_1160),
.Y(n_1213)
);

INVxp67_ASAP7_75t_SL g1214 ( 
.A(n_1199),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1177),
.B(n_1141),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1191),
.B(n_1141),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1185),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1194),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1178),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1195),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1175),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1176),
.B(n_1182),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1211),
.B(n_1197),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1200),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1205),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1210),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1206),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1217),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1218),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1220),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1219),
.Y(n_1231)
);

NAND2x1p5_ASAP7_75t_L g1232 ( 
.A(n_1207),
.B(n_1184),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_1202),
.B(n_1173),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1213),
.B(n_1222),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1207),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1209),
.Y(n_1236)
);

INVxp67_ASAP7_75t_L g1237 ( 
.A(n_1202),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1209),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1219),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1221),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1236),
.Y(n_1241)
);

NAND2x1_ASAP7_75t_L g1242 ( 
.A(n_1231),
.B(n_1180),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_1233),
.B(n_1203),
.Y(n_1243)
);

OAI321xp33_ASAP7_75t_L g1244 ( 
.A1(n_1232),
.A2(n_1187),
.A3(n_1152),
.B1(n_1212),
.B2(n_1204),
.C(n_1201),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1238),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1235),
.B(n_1214),
.Y(n_1246)
);

OAI21xp33_ASAP7_75t_L g1247 ( 
.A1(n_1232),
.A2(n_1184),
.B(n_1216),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1240),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1225),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1226),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1232),
.A2(n_1187),
.B(n_1114),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1227),
.Y(n_1252)
);

AOI21xp33_ASAP7_75t_L g1253 ( 
.A1(n_1224),
.A2(n_1179),
.B(n_1186),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1228),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1234),
.A2(n_1181),
.B(n_1124),
.C(n_1151),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1247),
.A2(n_1237),
.B1(n_1233),
.B2(n_1203),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1241),
.Y(n_1257)
);

OAI21xp33_ASAP7_75t_L g1258 ( 
.A1(n_1246),
.A2(n_1216),
.B(n_1208),
.Y(n_1258)
);

OAI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1244),
.A2(n_1190),
.B1(n_1215),
.B2(n_1198),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1250),
.B(n_1223),
.Y(n_1260)
);

NAND2xp33_ASAP7_75t_SL g1261 ( 
.A(n_1242),
.B(n_1118),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1245),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1248),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1261),
.B(n_1118),
.Y(n_1264)
);

NOR3xp33_ASAP7_75t_L g1265 ( 
.A(n_1259),
.B(n_1255),
.C(n_1253),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1257),
.B(n_1262),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1263),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1258),
.B(n_1161),
.Y(n_1268)
);

OAI21xp33_ASAP7_75t_SL g1269 ( 
.A1(n_1268),
.A2(n_1260),
.B(n_1243),
.Y(n_1269)
);

NOR3xp33_ASAP7_75t_L g1270 ( 
.A(n_1265),
.B(n_1259),
.C(n_1253),
.Y(n_1270)
);

NAND4xp25_ASAP7_75t_L g1271 ( 
.A(n_1264),
.B(n_1156),
.C(n_1251),
.D(n_1256),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1267),
.Y(n_1272)
);

NAND5xp2_ASAP7_75t_L g1273 ( 
.A(n_1266),
.B(n_1251),
.C(n_1254),
.D(n_1249),
.E(n_1252),
.Y(n_1273)
);

OAI211xp5_ASAP7_75t_L g1274 ( 
.A1(n_1265),
.A2(n_1246),
.B(n_1154),
.C(n_1239),
.Y(n_1274)
);

NOR3xp33_ASAP7_75t_L g1275 ( 
.A(n_1270),
.B(n_1158),
.C(n_1159),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1274),
.B(n_1231),
.Y(n_1276)
);

NOR3xp33_ASAP7_75t_L g1277 ( 
.A(n_1273),
.B(n_1164),
.C(n_1154),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1275),
.B(n_1272),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1277),
.B(n_1269),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1278),
.Y(n_1280)
);

OAI221xp5_ASAP7_75t_L g1281 ( 
.A1(n_1280),
.A2(n_1271),
.B1(n_1279),
.B2(n_1276),
.C(n_1125),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1281),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_SL g1283 ( 
.A1(n_1281),
.A2(n_1137),
.B1(n_1164),
.B2(n_1149),
.Y(n_1283)
);

AOI211xp5_ASAP7_75t_L g1284 ( 
.A1(n_1283),
.A2(n_1137),
.B(n_1148),
.C(n_1198),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1282),
.A2(n_1229),
.B1(n_1230),
.B2(n_1165),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_1285),
.A2(n_1134),
.B(n_1223),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1284),
.A2(n_1165),
.B(n_1163),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1287),
.A2(n_1130),
.B(n_1239),
.Y(n_1288)
);

OA22x2_ASAP7_75t_L g1289 ( 
.A1(n_1286),
.A2(n_1163),
.B1(n_1150),
.B2(n_1239),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1289),
.B(n_1288),
.Y(n_1290)
);

AO21x2_ASAP7_75t_L g1291 ( 
.A1(n_1290),
.A2(n_1157),
.B(n_1126),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1291),
.A2(n_1122),
.B1(n_1168),
.B2(n_1162),
.Y(n_1292)
);


endmodule