module real_jpeg_25586_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_242;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_167;
wire n_128;
wire n_179;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_1),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_1),
.B(n_125),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_111),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_1),
.A2(n_28),
.B(n_43),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_1),
.B(n_89),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_1),
.A2(n_25),
.B1(n_227),
.B2(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_1),
.A2(n_64),
.B(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_2),
.A2(n_64),
.B1(n_65),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_87),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_2),
.A2(n_87),
.B1(n_110),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_87),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_5),
.A2(n_71),
.B1(n_73),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_5),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_123),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_123),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_123),
.Y(n_227)
);

INVx8_ASAP7_75t_SL g63 ( 
.A(n_6),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_7),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_8),
.A2(n_40),
.B1(n_47),
.B2(n_48),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_8),
.A2(n_40),
.B1(n_64),
.B2(n_65),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_9),
.A2(n_50),
.B1(n_64),
.B2(n_65),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_10),
.A2(n_71),
.B1(n_73),
.B2(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_10),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_10),
.A2(n_64),
.B1(n_65),
.B2(n_78),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_78),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_78),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_11),
.A2(n_69),
.B1(n_73),
.B2(n_76),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_11),
.A2(n_64),
.B1(n_65),
.B2(n_76),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_76),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_76),
.Y(n_217)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_13),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_15),
.Y(n_120)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_15),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_150),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_149),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_127),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_20),
.B(n_127),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_92),
.C(n_102),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_21),
.A2(n_22),
.B1(n_92),
.B2(n_93),
.Y(n_167)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_56),
.B1(n_57),
.B2(n_91),
.Y(n_22)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_24),
.B(n_41),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_35),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_25),
.A2(n_118),
.B(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_25),
.A2(n_96),
.B(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_25),
.A2(n_118),
.B1(n_217),
.B2(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_25),
.A2(n_35),
.B(n_130),
.Y(n_251)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_26),
.B(n_39),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_26),
.A2(n_33),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_26),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_28),
.B1(n_43),
.B2(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_27),
.B(n_232),
.Y(n_231)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_38),
.B(n_111),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B(n_51),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_42),
.A2(n_46),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_42),
.B(n_53),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_42),
.A2(n_100),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_42),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_42),
.B(n_111),
.Y(n_225)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_SL g201 ( 
.A1(n_45),
.A2(n_48),
.B(n_111),
.C(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_48),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_47),
.B(n_84),
.Y(n_250)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI32xp33_ASAP7_75t_L g249 ( 
.A1(n_48),
.A2(n_64),
.A3(n_83),
.B1(n_243),
.B2(n_250),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_54),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_54),
.A2(n_134),
.B(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_54),
.A2(n_200),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_54),
.A2(n_208),
.B1(n_209),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_79),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_58),
.B(n_79),
.C(n_91),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_72),
.B2(n_77),
.Y(n_58)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_59),
.A2(n_77),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_68),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_60),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_62),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g108 ( 
.A1(n_61),
.A2(n_65),
.A3(n_74),
.B1(n_109),
.B2(n_112),
.Y(n_108)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_64),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_65),
.B1(n_83),
.B2(n_84),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_65),
.B(n_111),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_73),
.A2(n_109),
.B(n_111),
.Y(n_162)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_86),
.B(n_88),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_80),
.A2(n_82),
.B1(n_182),
.B2(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_81),
.B(n_90),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_81),
.A2(n_89),
.B1(n_105),
.B2(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_81),
.A2(n_89),
.B1(n_164),
.B2(n_181),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_86),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_82),
.A2(n_145),
.B(n_146),
.Y(n_144)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_99),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_99),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_95),
.A2(n_116),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_100),
.A2(n_101),
.B(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_100),
.A2(n_266),
.B(n_267),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_102),
.A2(n_103),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.C(n_121),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_121),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_108),
.A2(n_113),
.B1(n_114),
.B2(n_177),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_108),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_122),
.A2(n_124),
.B1(n_125),
.B2(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_125),
.B(n_142),
.Y(n_141)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_127),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_136),
.CI(n_148),
.CON(n_127),
.SN(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_131),
.B1(n_132),
.B2(n_135),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_129),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_147),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_189),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_169),
.B(n_188),
.Y(n_152)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_153),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_166),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_154),
.B(n_166),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.C(n_165),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_156),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_158),
.B(n_165),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_163),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_163),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_160),
.B(n_208),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_170),
.B(n_173),
.Y(n_278)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_178),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_174),
.B(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_176),
.A2(n_178),
.B1(n_179),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_176),
.Y(n_275)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.C(n_184),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_180),
.B(n_260),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_183),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_277),
.C(n_278),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_271),
.B(n_276),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_255),
.B(n_270),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_236),
.B(n_254),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_213),
.B(n_235),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_203),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_195),
.B(n_203),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_197),
.B1(n_201),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_201),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_211),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_210),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_210),
.C(n_211),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_207),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_212),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_223),
.B(n_234),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_221),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_215),
.B(n_221),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_219),
.Y(n_230)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_228),
.B(n_233),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_225),
.B(n_226),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_237),
.B(n_238),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_248),
.B1(n_252),
.B2(n_253),
.Y(n_238)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.Y(n_239)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_244),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_247),
.C(n_252),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_251),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_256),
.B(n_257),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_262),
.B2(n_263),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_265),
.C(n_268),
.Y(n_272)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_268),
.B2(n_269),
.Y(n_263)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_264),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_272),
.B(n_273),
.Y(n_276)
);


endmodule