module fake_jpeg_10032_n_35 (n_3, n_2, n_1, n_0, n_4, n_5, n_35);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_35;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_5),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_7),
.B(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

NOR3xp33_ASAP7_75t_SL g18 ( 
.A(n_15),
.B(n_16),
.C(n_8),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_0),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_16),
.A2(n_8),
.B1(n_6),
.B2(n_9),
.Y(n_17)
);

OAI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_9),
.B1(n_15),
.B2(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_20),
.B(n_6),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_22),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_12),
.B1(n_13),
.B2(n_10),
.Y(n_23)
);

OAI21xp33_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_24),
.B(n_1),
.Y(n_27)
);

AND2x6_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_27),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g28 ( 
.A(n_25),
.B(n_21),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_23),
.C(n_19),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_31),
.C(n_29),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_1),
.C(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_2),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_2),
.C(n_3),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_3),
.Y(n_35)
);


endmodule