module fake_netlist_6_617_n_1693 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1693);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1693;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_153),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_117),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_140),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_17),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_2),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_132),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_31),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_120),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_52),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_29),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_24),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_88),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_61),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_124),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_90),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_60),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_12),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_104),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_13),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_23),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_89),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_127),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_131),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_67),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_92),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

INVxp33_ASAP7_75t_SL g191 ( 
.A(n_62),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_71),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_75),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_142),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_84),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_39),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_151),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_82),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_58),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_107),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_68),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_64),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_114),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_13),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_17),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_94),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_34),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_121),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_126),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_10),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_109),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_3),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_20),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_125),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_35),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_111),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_18),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_47),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_23),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_21),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_48),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_63),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_45),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_44),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_81),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_18),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_74),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_7),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_72),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_41),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_105),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_44),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_134),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_26),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_16),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_148),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_0),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_141),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_98),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_155),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_99),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_122),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_5),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_24),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_19),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_139),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_101),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_34),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_96),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_145),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_39),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_95),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_97),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_130),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_7),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_138),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_33),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_46),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_118),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_49),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_137),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_6),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_16),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_40),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_26),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_115),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_76),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_78),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_93),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_29),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_106),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_0),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_15),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_53),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_133),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_91),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_10),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_85),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_87),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_35),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_65),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_66),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_3),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_4),
.Y(n_284)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_51),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_21),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_12),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_116),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_36),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_146),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_43),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_5),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_110),
.Y(n_293)
);

BUFx2_ASAP7_75t_R g294 ( 
.A(n_56),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_154),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_32),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_28),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_30),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_11),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_2),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_77),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_73),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_9),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_54),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_129),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_103),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_69),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_28),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_80),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_25),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_197),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_158),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_180),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_241),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_303),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_229),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_258),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_176),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_301),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_303),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_201),
.Y(n_324)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_162),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_213),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_183),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_183),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_158),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_196),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_170),
.Y(n_331)
);

INVxp33_ASAP7_75t_SL g332 ( 
.A(n_162),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_196),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_205),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_203),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_205),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_206),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_220),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_220),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_281),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_302),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_209),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_285),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_198),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_299),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_285),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_238),
.Y(n_347)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_163),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_178),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_211),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_221),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_285),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_222),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_225),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_299),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_227),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_231),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_310),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_182),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_233),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_236),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_285),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_210),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_239),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_285),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_242),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_246),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_217),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_247),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_178),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_219),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_249),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_230),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_234),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_243),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_245),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_253),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_251),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_257),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_265),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_308),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_312),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_344),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_351),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_364),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_312),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_313),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_313),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_317),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_344),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_321),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_317),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_344),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_318),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_318),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_344),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_323),
.B(n_188),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_323),
.Y(n_398)
);

BUFx12f_ASAP7_75t_L g399 ( 
.A(n_311),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_358),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_200),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_358),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_359),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_319),
.B(n_191),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_352),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_359),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_366),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_363),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_343),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_352),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_362),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_362),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_314),
.B(n_200),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_365),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_365),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_363),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_368),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_343),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_314),
.B(n_188),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_367),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_368),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_371),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_369),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_343),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_314),
.B(n_259),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_329),
.B(n_259),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_329),
.B(n_199),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_320),
.B(n_278),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_326),
.A2(n_263),
.B1(n_272),
.B2(n_277),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_346),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_329),
.B(n_278),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_371),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_340),
.B(n_175),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_349),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_373),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_349),
.B(n_156),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_349),
.B(n_199),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_373),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_R g439 ( 
.A(n_324),
.B(n_254),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_341),
.B(n_223),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_346),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_346),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_327),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_345),
.B(n_156),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_327),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_315),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_434),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_304),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_399),
.B(n_215),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_405),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_384),
.Y(n_451)
);

INVx6_ASAP7_75t_L g452 ( 
.A(n_397),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_405),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_409),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_405),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_433),
.B(n_335),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_409),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_410),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_410),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_409),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_409),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_L g462 ( 
.A(n_401),
.B(n_198),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_409),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_394),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_394),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_410),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_404),
.A2(n_316),
.B1(n_377),
.B2(n_354),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_411),
.Y(n_468)
);

AND3x1_ASAP7_75t_L g469 ( 
.A(n_404),
.B(n_215),
.C(n_345),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_433),
.B(n_337),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_411),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_409),
.Y(n_473)
);

OR2x6_ASAP7_75t_L g474 ( 
.A(n_399),
.B(n_446),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_409),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_411),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_409),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_414),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_414),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_384),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_440),
.B(n_342),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_414),
.Y(n_482)
);

OAI21xp33_ASAP7_75t_SL g483 ( 
.A1(n_428),
.A2(n_174),
.B(n_161),
.Y(n_483)
);

AO21x2_ASAP7_75t_L g484 ( 
.A1(n_436),
.A2(n_167),
.B(n_159),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_440),
.B(n_350),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_434),
.B(n_353),
.Y(n_486)
);

BUFx10_ASAP7_75t_L g487 ( 
.A(n_428),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_441),
.Y(n_488)
);

INVxp33_ASAP7_75t_L g489 ( 
.A(n_429),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_415),
.Y(n_490)
);

NAND3xp33_ASAP7_75t_L g491 ( 
.A(n_444),
.B(n_357),
.C(n_356),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

BUFx10_ASAP7_75t_L g493 ( 
.A(n_419),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_415),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_400),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_441),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_397),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_436),
.B(n_315),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_415),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_402),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_401),
.B(n_360),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_402),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_418),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_385),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_419),
.B(n_361),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_403),
.Y(n_506)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_441),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_418),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_418),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_396),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_439),
.B(n_347),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_427),
.Y(n_512)
);

INVx8_ASAP7_75t_L g513 ( 
.A(n_399),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_424),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_424),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_419),
.B(n_372),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_439),
.B(n_347),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_397),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_441),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_382),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_419),
.B(n_326),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_444),
.B(n_325),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_424),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_382),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_397),
.B(n_304),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_397),
.A2(n_332),
.B1(n_348),
.B2(n_192),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_446),
.B(n_157),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_403),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_446),
.B(n_157),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_386),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_441),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_427),
.B(n_160),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_427),
.B(n_160),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_385),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_430),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_437),
.B(n_164),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_413),
.A2(n_174),
.B(n_161),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_442),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_437),
.A2(n_322),
.B1(n_173),
.B2(n_194),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_406),
.Y(n_540)
);

BUFx4f_ASAP7_75t_L g541 ( 
.A(n_443),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_406),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_437),
.Y(n_543)
);

AND2x2_ASAP7_75t_SL g544 ( 
.A(n_413),
.B(n_192),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_425),
.B(n_307),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_391),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_430),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_430),
.Y(n_548)
);

BUFx4f_ASAP7_75t_L g549 ( 
.A(n_443),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_408),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_408),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_425),
.B(n_307),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_412),
.Y(n_553)
);

CKINVDCx11_ASAP7_75t_R g554 ( 
.A(n_391),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_416),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_426),
.B(n_256),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_426),
.B(n_164),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_431),
.A2(n_207),
.B1(n_264),
.B2(n_248),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_442),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_431),
.A2(n_195),
.B1(n_202),
.B2(n_250),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_386),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_387),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_429),
.B(n_166),
.Y(n_563)
);

AOI21x1_ASAP7_75t_L g564 ( 
.A1(n_387),
.A2(n_202),
.B(n_195),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_442),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_416),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_388),
.Y(n_567)
);

INVxp33_ASAP7_75t_L g568 ( 
.A(n_417),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_442),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_412),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_407),
.B(n_166),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_396),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_412),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_417),
.Y(n_574)
);

BUFx8_ASAP7_75t_SL g575 ( 
.A(n_407),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_388),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_412),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_389),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_442),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_389),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_396),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_392),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_420),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_396),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_392),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_396),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_L g587 ( 
.A(n_443),
.B(n_198),
.Y(n_587)
);

BUFx6f_ASAP7_75t_SL g588 ( 
.A(n_421),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_420),
.B(n_168),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_443),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_423),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_421),
.Y(n_592)
);

INVxp33_ASAP7_75t_L g593 ( 
.A(n_422),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_568),
.B(n_423),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_450),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_497),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_L g597 ( 
.A(n_505),
.B(n_285),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_501),
.B(n_395),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_512),
.B(n_395),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_522),
.B(n_204),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_481),
.B(n_168),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_450),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_447),
.B(n_355),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_497),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_456),
.B(n_171),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_593),
.B(n_355),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_453),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_518),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_447),
.B(n_331),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_453),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_512),
.B(n_398),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_544),
.B(n_398),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_518),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_471),
.B(n_171),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_544),
.A2(n_260),
.B1(n_194),
.B2(n_193),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_543),
.B(n_487),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_566),
.B(n_445),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g618 ( 
.A(n_513),
.B(n_294),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_566),
.B(n_445),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_543),
.B(n_376),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_574),
.B(n_445),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_487),
.B(n_422),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_485),
.B(n_173),
.Y(n_623)
);

INVxp67_ASAP7_75t_SL g624 ( 
.A(n_488),
.Y(n_624)
);

NOR2x1p5_ASAP7_75t_L g625 ( 
.A(n_498),
.B(n_163),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_448),
.B(n_432),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_452),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_455),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_448),
.B(n_432),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_455),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_487),
.B(n_179),
.Y(n_631)
);

OAI22xp33_ASAP7_75t_L g632 ( 
.A1(n_498),
.A2(n_279),
.B1(n_306),
.B2(n_250),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_574),
.B(n_445),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_458),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_467),
.B(n_179),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_546),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_470),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_452),
.Y(n_638)
);

OR2x6_ASAP7_75t_L g639 ( 
.A(n_513),
.B(n_374),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_452),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_510),
.B(n_198),
.Y(n_641)
);

A2O1A1Ixp33_ASAP7_75t_L g642 ( 
.A1(n_537),
.A2(n_306),
.B(n_279),
.C(n_269),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_452),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_458),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_486),
.B(n_181),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_470),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_L g647 ( 
.A(n_516),
.B(n_285),
.Y(n_647)
);

NOR2x1p5_ASAP7_75t_L g648 ( 
.A(n_491),
.B(n_165),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_510),
.B(n_572),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_526),
.B(n_435),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_563),
.B(n_181),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_492),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_459),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_556),
.B(n_185),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_495),
.B(n_445),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_500),
.B(n_502),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_448),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_SL g658 ( 
.A(n_588),
.B(n_286),
.Y(n_658)
);

OAI221xp5_ASAP7_75t_L g659 ( 
.A1(n_483),
.A2(n_435),
.B1(n_438),
.B2(n_172),
.C(n_240),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_459),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_521),
.B(n_185),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_493),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_510),
.B(n_198),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_466),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_466),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_493),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_506),
.B(n_528),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_540),
.B(n_443),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_542),
.B(n_550),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_468),
.Y(n_670)
);

CKINVDCx11_ASAP7_75t_R g671 ( 
.A(n_554),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_551),
.B(n_443),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_468),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_510),
.B(n_285),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_472),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_557),
.B(n_186),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_555),
.B(n_443),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_472),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_592),
.B(n_443),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_520),
.B(n_438),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_532),
.B(n_186),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_479),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_520),
.B(n_374),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_484),
.A2(n_560),
.B1(n_489),
.B2(n_462),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_493),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_464),
.B(n_252),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_465),
.B(n_252),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_539),
.B(n_187),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_524),
.B(n_269),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_533),
.B(n_187),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_524),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_530),
.B(n_383),
.Y(n_692)
);

INVxp33_ASAP7_75t_SL g693 ( 
.A(n_451),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_536),
.B(n_193),
.Y(n_694)
);

NAND2xp33_ASAP7_75t_L g695 ( 
.A(n_510),
.B(n_267),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_561),
.B(n_383),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_583),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_562),
.B(n_383),
.Y(n_698)
);

INVxp33_ASAP7_75t_SL g699 ( 
.A(n_451),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_511),
.B(n_375),
.Y(n_700)
);

AOI221xp5_ASAP7_75t_L g701 ( 
.A1(n_469),
.A2(n_284),
.B1(n_283),
.B2(n_165),
.C(n_287),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_572),
.B(n_177),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_525),
.A2(n_393),
.B(n_390),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_527),
.B(n_267),
.Y(n_704)
);

NOR3xp33_ASAP7_75t_L g705 ( 
.A(n_571),
.B(n_375),
.C(n_381),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_567),
.B(n_390),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_529),
.B(n_268),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_588),
.A2(n_276),
.B1(n_268),
.B2(n_271),
.Y(n_708)
);

BUFx6f_ASAP7_75t_SL g709 ( 
.A(n_474),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_545),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_517),
.B(n_271),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_576),
.B(n_390),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_576),
.B(n_393),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_479),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_572),
.Y(n_715)
);

A2O1A1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_578),
.A2(n_218),
.B(n_184),
.C(n_189),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_552),
.B(n_378),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_578),
.B(n_393),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_580),
.B(n_274),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_558),
.B(n_378),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_482),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_572),
.B(n_584),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_589),
.Y(n_723)
);

AO221x1_ASAP7_75t_L g724 ( 
.A1(n_572),
.A2(n_305),
.B1(n_290),
.B2(n_266),
.C(n_261),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_513),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_580),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_581),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_582),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_582),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_482),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_484),
.A2(n_214),
.B1(n_309),
.B2(n_190),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_585),
.B(n_274),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_490),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_490),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_494),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_488),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_531),
.B(n_569),
.Y(n_737)
);

OAI22xp33_ASAP7_75t_L g738 ( 
.A1(n_449),
.A2(n_216),
.B1(n_208),
.B2(n_288),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_588),
.B(n_275),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_531),
.B(n_293),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_494),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_581),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_513),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_581),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_584),
.B(n_295),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_584),
.B(n_275),
.Y(n_746)
);

BUFx6f_ASAP7_75t_SL g747 ( 
.A(n_474),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_499),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_484),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_591),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_531),
.B(n_276),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_591),
.B(n_379),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_569),
.B(n_282),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_584),
.B(n_282),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_569),
.B(n_212),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_584),
.B(n_224),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_488),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_496),
.B(n_538),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_595),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_627),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_601),
.A2(n_559),
.B1(n_538),
.B2(n_496),
.Y(n_761)
);

AND3x2_ASAP7_75t_SL g762 ( 
.A(n_600),
.B(n_554),
.C(n_297),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_600),
.B(n_480),
.Y(n_763)
);

AND2x6_ASAP7_75t_L g764 ( 
.A(n_727),
.B(n_457),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_636),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_601),
.A2(n_559),
.B1(n_538),
.B2(n_496),
.Y(n_766)
);

NAND2x1p5_ASAP7_75t_L g767 ( 
.A(n_662),
.B(n_559),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_598),
.B(n_565),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_727),
.B(n_565),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_605),
.B(n_480),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_742),
.B(n_565),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_622),
.B(n_504),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_626),
.B(n_449),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_620),
.B(n_504),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_742),
.B(n_476),
.Y(n_775)
);

AND2x6_ASAP7_75t_SL g776 ( 
.A(n_651),
.B(n_474),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_SL g777 ( 
.A(n_605),
.B(n_534),
.C(n_287),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_671),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_637),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_626),
.B(n_449),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_629),
.B(n_449),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_606),
.B(n_534),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_614),
.B(n_575),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_602),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_602),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_646),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_607),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_627),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_744),
.B(n_476),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_607),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_614),
.B(n_575),
.Y(n_791)
);

NOR3xp33_ASAP7_75t_SL g792 ( 
.A(n_701),
.B(n_284),
.C(n_169),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_609),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_680),
.Y(n_794)
);

NAND2xp33_ASAP7_75t_SL g795 ( 
.A(n_725),
.B(n_169),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_638),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_629),
.B(n_474),
.Y(n_797)
);

OR2x6_ASAP7_75t_L g798 ( 
.A(n_639),
.B(n_379),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_658),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_638),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_680),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_691),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_616),
.B(n_586),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_610),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_752),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_744),
.B(n_478),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_604),
.Y(n_807)
);

AND2x6_ASAP7_75t_L g808 ( 
.A(n_662),
.B(n_457),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_717),
.B(n_478),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_662),
.B(n_586),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_662),
.B(n_586),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_750),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_731),
.A2(n_462),
.B1(n_586),
.B2(n_579),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_666),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_710),
.A2(n_586),
.B1(n_475),
.B2(n_460),
.Y(n_815)
);

BUFx4f_ASAP7_75t_L g816 ( 
.A(n_639),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_631),
.B(n_457),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_612),
.A2(n_477),
.B(n_460),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_731),
.A2(n_579),
.B1(n_499),
.B2(n_535),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_693),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_726),
.B(n_503),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_594),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_603),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_697),
.Y(n_824)
);

BUFx12f_ASAP7_75t_L g825 ( 
.A(n_625),
.Y(n_825)
);

AOI221xp5_ASAP7_75t_SL g826 ( 
.A1(n_632),
.A2(n_380),
.B1(n_381),
.B2(n_333),
.C(n_334),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_610),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_654),
.A2(n_645),
.B1(n_608),
.B2(n_613),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_631),
.B(n_460),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_728),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_729),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_628),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_650),
.B(n_503),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_749),
.B(n_508),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_700),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_604),
.B(n_508),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_640),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_639),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_684),
.B(n_509),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_736),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_757),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_628),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_684),
.B(n_509),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_652),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_596),
.Y(n_845)
);

BUFx4f_ASAP7_75t_L g846 ( 
.A(n_743),
.Y(n_846)
);

OR2x6_ASAP7_75t_L g847 ( 
.A(n_723),
.B(n_380),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_624),
.B(n_514),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_640),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_699),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_651),
.A2(n_535),
.B1(n_514),
.B2(n_515),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_720),
.B(n_270),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_630),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_654),
.B(n_515),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_704),
.A2(n_547),
.B1(n_548),
.B2(n_523),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_630),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_657),
.B(n_463),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_719),
.Y(n_858)
);

NOR2x1_ASAP7_75t_L g859 ( 
.A(n_648),
.B(n_463),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_643),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_683),
.B(n_523),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_666),
.Y(n_862)
);

INVx5_ASAP7_75t_L g863 ( 
.A(n_666),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_634),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_683),
.B(n_547),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_599),
.B(n_548),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_611),
.B(n_463),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_656),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_667),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_739),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_666),
.B(n_454),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_634),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_644),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_617),
.B(n_473),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_619),
.B(n_473),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_644),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_643),
.B(n_473),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_653),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_621),
.B(n_475),
.Y(n_879)
);

NOR3xp33_ASAP7_75t_L g880 ( 
.A(n_635),
.B(n_228),
.C(n_232),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_653),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_660),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_660),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_715),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_664),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_645),
.B(n_475),
.Y(n_886)
);

NAND2xp33_ASAP7_75t_SL g887 ( 
.A(n_709),
.B(n_270),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_SL g888 ( 
.A1(n_618),
.A2(n_707),
.B1(n_704),
.B2(n_711),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_685),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_669),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_665),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_633),
.B(n_477),
.Y(n_892)
);

O2A1O1Ixp5_ASAP7_75t_L g893 ( 
.A1(n_642),
.A2(n_564),
.B(n_541),
.C(n_549),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_665),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_685),
.B(n_454),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_670),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_739),
.Y(n_897)
);

AOI221xp5_ASAP7_75t_L g898 ( 
.A1(n_707),
.A2(n_273),
.B1(n_280),
.B2(n_283),
.C(n_300),
.Y(n_898)
);

OR2x4_ASAP7_75t_L g899 ( 
.A(n_711),
.B(n_661),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_685),
.B(n_454),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_689),
.B(n_477),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_670),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_685),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_615),
.A2(n_280),
.B1(n_298),
.B2(n_297),
.Y(n_904)
);

BUFx10_ASAP7_75t_L g905 ( 
.A(n_661),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_673),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_673),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_675),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_675),
.B(n_553),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_678),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_678),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_682),
.B(n_553),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_682),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_755),
.B(n_454),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_755),
.B(n_454),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_676),
.B(n_681),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_714),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_659),
.A2(n_570),
.B1(n_577),
.B2(n_573),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_714),
.Y(n_919)
);

INVxp67_ASAP7_75t_L g920 ( 
.A(n_719),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_721),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_758),
.Y(n_922)
);

BUFx4f_ASAP7_75t_L g923 ( 
.A(n_721),
.Y(n_923)
);

BUFx5_ASAP7_75t_L g924 ( 
.A(n_715),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_597),
.A2(n_461),
.B1(n_590),
.B2(n_577),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_647),
.A2(n_461),
.B1(n_590),
.B2(n_573),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_681),
.B(n_328),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_737),
.A2(n_549),
.B(n_541),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_730),
.Y(n_929)
);

AO21x1_ASAP7_75t_L g930 ( 
.A1(n_702),
.A2(n_564),
.B(n_587),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_730),
.B(n_570),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_676),
.B(n_461),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_733),
.B(n_461),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_690),
.A2(n_461),
.B1(n_590),
.B2(n_587),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_690),
.A2(n_549),
.B1(n_541),
.B2(n_226),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_694),
.A2(n_235),
.B1(n_237),
.B2(n_244),
.Y(n_936)
);

INVx4_ASAP7_75t_L g937 ( 
.A(n_709),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_733),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_802),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_858),
.B(n_732),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_759),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_858),
.B(n_732),
.Y(n_942)
);

OR2x6_ASAP7_75t_SL g943 ( 
.A(n_778),
.B(n_273),
.Y(n_943)
);

NOR3xp33_ASAP7_75t_L g944 ( 
.A(n_888),
.B(n_688),
.C(n_694),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_888),
.B(n_708),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_920),
.B(n_623),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_914),
.A2(n_722),
.B(n_649),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_920),
.B(n_751),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_915),
.A2(n_649),
.B(n_722),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_782),
.B(n_753),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_824),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_769),
.A2(n_740),
.B(n_754),
.Y(n_952)
);

AOI22x1_ASAP7_75t_L g953 ( 
.A1(n_928),
.A2(n_927),
.B1(n_785),
.B2(n_787),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_769),
.A2(n_746),
.B(n_754),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_784),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_774),
.B(n_738),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_890),
.B(n_746),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_771),
.A2(n_655),
.B(n_698),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_765),
.Y(n_959)
);

AOI221x1_ASAP7_75t_L g960 ( 
.A1(n_880),
.A2(n_777),
.B1(n_817),
.B2(n_829),
.C(n_886),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_763),
.B(n_747),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_771),
.A2(n_706),
.B(n_712),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_775),
.A2(n_713),
.B(n_696),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_916),
.A2(n_756),
.B(n_686),
.C(n_687),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_770),
.A2(n_679),
.B(n_668),
.C(n_672),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_777),
.A2(n_716),
.B(n_705),
.C(n_695),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_890),
.B(n_734),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_899),
.B(n_747),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_868),
.B(n_734),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_790),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_804),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_827),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_775),
.A2(n_806),
.B(n_789),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_789),
.A2(n_692),
.B(n_718),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_806),
.A2(n_677),
.B(n_745),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_869),
.B(n_735),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_899),
.B(n_702),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_835),
.B(n_748),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_863),
.A2(n_745),
.B(n_703),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_793),
.B(n_334),
.Y(n_980)
);

NOR2x1_ASAP7_75t_L g981 ( 
.A(n_820),
.B(n_674),
.Y(n_981)
);

OAI21xp33_ASAP7_75t_L g982 ( 
.A1(n_898),
.A2(n_298),
.B(n_296),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_768),
.B(n_741),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_863),
.A2(n_674),
.B(n_641),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_839),
.A2(n_748),
.B1(n_741),
.B2(n_735),
.Y(n_985)
);

BUFx4f_ASAP7_75t_L g986 ( 
.A(n_825),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_863),
.A2(n_663),
.B(n_641),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_863),
.A2(n_663),
.B(n_519),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_862),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_R g990 ( 
.A(n_799),
.B(n_296),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_R g991 ( 
.A(n_850),
.B(n_292),
.Y(n_991)
);

NAND2x1p5_ASAP7_75t_L g992 ( 
.A(n_814),
.B(n_507),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_862),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_839),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_793),
.B(n_255),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_768),
.B(n_724),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_843),
.A2(n_291),
.B1(n_262),
.B2(n_339),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_832),
.Y(n_998)
);

INVx4_ASAP7_75t_L g999 ( 
.A(n_862),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_903),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_905),
.B(n_519),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_805),
.B(n_1),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_SL g1003 ( 
.A1(n_783),
.A2(n_339),
.B1(n_338),
.B2(n_336),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_905),
.B(n_519),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_870),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_828),
.A2(n_519),
.B1(n_507),
.B2(n_338),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_903),
.Y(n_1007)
);

OAI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_897),
.A2(n_336),
.B1(n_333),
.B2(n_330),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_830),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_772),
.B(n_1),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_903),
.Y(n_1011)
);

O2A1O1Ixp5_ASAP7_75t_L g1012 ( 
.A1(n_932),
.A2(n_330),
.B(n_328),
.C(n_149),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_814),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_822),
.B(n_4),
.Y(n_1014)
);

BUFx12f_ASAP7_75t_L g1015 ( 
.A(n_937),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_880),
.A2(n_519),
.B(n_507),
.C(n_9),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_852),
.A2(n_6),
.B(n_8),
.C(n_11),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_800),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_928),
.A2(n_507),
.B(n_144),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_884),
.A2(n_507),
.B(n_135),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_904),
.A2(n_8),
.B(n_14),
.C(n_15),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_794),
.B(n_128),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_823),
.B(n_14),
.Y(n_1023)
);

O2A1O1Ixp5_ASAP7_75t_L g1024 ( 
.A1(n_893),
.A2(n_112),
.B(n_102),
.C(n_100),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_831),
.B(n_19),
.Y(n_1025)
);

OAI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_792),
.A2(n_20),
.B(n_22),
.Y(n_1026)
);

OA22x2_ASAP7_75t_L g1027 ( 
.A1(n_847),
.A2(n_22),
.B1(n_25),
.B2(n_27),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_776),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_842),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_812),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_884),
.A2(n_83),
.B(n_79),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_856),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_801),
.B(n_59),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_843),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_889),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_864),
.Y(n_1036)
);

NAND2x1p5_ASAP7_75t_L g1037 ( 
.A(n_889),
.B(n_70),
.Y(n_1037)
);

NAND2x1_ASAP7_75t_L g1038 ( 
.A(n_808),
.B(n_57),
.Y(n_1038)
);

BUFx10_ASAP7_75t_L g1039 ( 
.A(n_791),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_937),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_867),
.A2(n_55),
.B(n_50),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_847),
.B(n_32),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_800),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_847),
.Y(n_1044)
);

BUFx12f_ASAP7_75t_L g1045 ( 
.A(n_797),
.Y(n_1045)
);

O2A1O1Ixp5_ASAP7_75t_L g1046 ( 
.A1(n_893),
.A2(n_33),
.B(n_36),
.C(n_37),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_809),
.B(n_37),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_797),
.B(n_38),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_867),
.A2(n_43),
.B(n_40),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_SL g1050 ( 
.A(n_816),
.B(n_38),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_800),
.B(n_41),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_844),
.B(n_42),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_807),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_779),
.A2(n_786),
.B(n_833),
.C(n_809),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_845),
.B(n_42),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_833),
.A2(n_813),
.B1(n_854),
.B2(n_792),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_807),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_874),
.A2(n_875),
.B(n_879),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_859),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_773),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_854),
.B(n_866),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_SL g1062 ( 
.A(n_887),
.B(n_904),
.C(n_795),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_773),
.B(n_780),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_807),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_780),
.B(n_781),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_901),
.A2(n_848),
.B(n_836),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_803),
.A2(n_865),
.B(n_861),
.C(n_841),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_838),
.B(n_922),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_922),
.B(n_798),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_781),
.B(n_798),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_853),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_901),
.A2(n_848),
.B(n_836),
.Y(n_1072)
);

NAND2x1_ASAP7_75t_SL g1073 ( 
.A(n_760),
.B(n_788),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_816),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_861),
.A2(n_865),
.B(n_818),
.C(n_840),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_818),
.A2(n_923),
.B(n_761),
.C(n_766),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_846),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_973),
.A2(n_923),
.B(n_866),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_940),
.B(n_922),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_942),
.B(n_936),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_939),
.Y(n_1081)
);

BUFx10_ASAP7_75t_L g1082 ( 
.A(n_968),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_948),
.B(n_760),
.Y(n_1083)
);

AOI21x1_ASAP7_75t_L g1084 ( 
.A1(n_954),
.A2(n_900),
.B(n_871),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1014),
.B(n_798),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_957),
.B(n_796),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1066),
.A2(n_895),
.B(n_811),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_SL g1088 ( 
.A1(n_1076),
.A2(n_934),
.B(n_767),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_953),
.A2(n_1058),
.B(n_949),
.Y(n_1089)
);

OAI22x1_ASAP7_75t_L g1090 ( 
.A1(n_945),
.A2(n_762),
.B1(n_810),
.B2(n_815),
.Y(n_1090)
);

NOR2xp67_ASAP7_75t_L g1091 ( 
.A(n_1013),
.B(n_860),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_1053),
.Y(n_1092)
);

OAI22x1_ASAP7_75t_L g1093 ( 
.A1(n_1010),
.A2(n_762),
.B1(n_938),
.B2(n_917),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_1005),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_947),
.A2(n_879),
.B(n_892),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1072),
.A2(n_874),
.B(n_875),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_1030),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1061),
.B(n_788),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1056),
.A2(n_952),
.B(n_958),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1056),
.A2(n_962),
.B(n_963),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_976),
.B(n_796),
.Y(n_1101)
);

AOI221x1_ASAP7_75t_L g1102 ( 
.A1(n_944),
.A2(n_892),
.B1(n_834),
.B2(n_821),
.C(n_913),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_951),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_1063),
.B(n_1065),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_1063),
.B(n_877),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_967),
.B(n_821),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_977),
.A2(n_935),
.B(n_860),
.C(n_849),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_951),
.Y(n_1108)
);

AOI221xp5_ASAP7_75t_SL g1109 ( 
.A1(n_1026),
.A2(n_911),
.B1(n_907),
.B2(n_896),
.C(n_894),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_946),
.B(n_857),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_974),
.A2(n_834),
.B(n_933),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_1044),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_975),
.A2(n_933),
.B(n_924),
.Y(n_1113)
);

OA21x2_ASAP7_75t_L g1114 ( 
.A1(n_1024),
.A2(n_826),
.B(n_930),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_1065),
.B(n_877),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1054),
.A2(n_767),
.B1(n_855),
.B2(n_851),
.Y(n_1116)
);

AO31x2_ASAP7_75t_L g1117 ( 
.A1(n_960),
.A2(n_876),
.A3(n_882),
.B(n_881),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_985),
.A2(n_931),
.B(n_912),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_985),
.A2(n_931),
.B(n_912),
.Y(n_1119)
);

INVx5_ASAP7_75t_L g1120 ( 
.A(n_1000),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_965),
.A2(n_924),
.B(n_909),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_978),
.B(n_929),
.Y(n_1122)
);

NOR4xp25_ASAP7_75t_L g1123 ( 
.A(n_1021),
.B(n_878),
.C(n_873),
.D(n_918),
.Y(n_1123)
);

NOR2xp67_ASAP7_75t_L g1124 ( 
.A(n_1013),
.B(n_849),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_980),
.B(n_1060),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_966),
.A2(n_837),
.B(n_857),
.C(n_919),
.Y(n_1126)
);

AOI221xp5_ASAP7_75t_L g1127 ( 
.A1(n_982),
.A2(n_902),
.B1(n_921),
.B2(n_908),
.C(n_906),
.Y(n_1127)
);

AOI21x1_ASAP7_75t_SL g1128 ( 
.A1(n_996),
.A2(n_909),
.B(n_808),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1009),
.A2(n_819),
.B1(n_910),
.B2(n_885),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_961),
.B(n_837),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_1070),
.B(n_1040),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_979),
.A2(n_924),
.B(n_764),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1019),
.A2(n_891),
.B(n_883),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_1074),
.Y(n_1134)
);

AOI22x1_ASAP7_75t_L g1135 ( 
.A1(n_984),
.A2(n_872),
.B1(n_764),
.B2(n_808),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_1075),
.A2(n_925),
.A3(n_926),
.B(n_764),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_983),
.A2(n_924),
.B(n_808),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_956),
.A2(n_764),
.B1(n_808),
.B2(n_924),
.Y(n_1138)
);

NOR2xp67_ASAP7_75t_L g1139 ( 
.A(n_1035),
.B(n_764),
.Y(n_1139)
);

CKINVDCx6p67_ASAP7_75t_R g1140 ( 
.A(n_1015),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1071),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1067),
.A2(n_924),
.B(n_987),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_941),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_964),
.A2(n_1046),
.B(n_1012),
.Y(n_1144)
);

NOR4xp25_ASAP7_75t_L g1145 ( 
.A(n_1017),
.B(n_1026),
.C(n_1034),
.D(n_982),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_1016),
.A2(n_1006),
.A3(n_1034),
.B(n_997),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_1048),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_950),
.B(n_1047),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1020),
.A2(n_988),
.B(n_1038),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1041),
.A2(n_1049),
.B(n_1025),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1069),
.B(n_969),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1031),
.A2(n_1035),
.B(n_1022),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1068),
.B(n_997),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1052),
.A2(n_1062),
.B1(n_1027),
.B2(n_1033),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_955),
.Y(n_1155)
);

INVx3_ASAP7_75t_SL g1156 ( 
.A(n_1028),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1055),
.A2(n_995),
.B(n_981),
.C(n_1033),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1001),
.A2(n_1004),
.B(n_1059),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1070),
.B(n_1050),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1073),
.A2(n_1037),
.B(n_970),
.Y(n_1160)
);

OA21x2_ASAP7_75t_L g1161 ( 
.A1(n_971),
.A2(n_1029),
.B(n_972),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_998),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1037),
.A2(n_1036),
.B(n_1032),
.Y(n_1163)
);

O2A1O1Ixp5_ASAP7_75t_SL g1164 ( 
.A1(n_1051),
.A2(n_994),
.B(n_1011),
.C(n_989),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1042),
.B(n_1048),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1045),
.Y(n_1166)
);

OAI22x1_ASAP7_75t_L g1167 ( 
.A1(n_1023),
.A2(n_1002),
.B1(n_1077),
.B2(n_1050),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_SL g1168 ( 
.A(n_986),
.B(n_999),
.Y(n_1168)
);

AO31x2_ASAP7_75t_L g1169 ( 
.A1(n_994),
.A2(n_1008),
.A3(n_1003),
.B(n_992),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1003),
.A2(n_1039),
.B1(n_1064),
.B2(n_989),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_992),
.A2(n_1064),
.B(n_1011),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_993),
.A2(n_1007),
.B(n_1000),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1007),
.A2(n_1057),
.B(n_1053),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_986),
.Y(n_1174)
);

AO32x2_ASAP7_75t_L g1175 ( 
.A1(n_1039),
.A2(n_1053),
.A3(n_1057),
.B1(n_1018),
.B2(n_1043),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1057),
.A2(n_1018),
.B(n_1043),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1018),
.B(n_1043),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_991),
.B(n_990),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_943),
.A2(n_960),
.A3(n_1076),
.B(n_1056),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_SL g1180 ( 
.A(n_944),
.B(n_888),
.C(n_600),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_959),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_953),
.A2(n_1058),
.B(n_949),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_944),
.A2(n_916),
.B(n_600),
.C(n_601),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_944),
.A2(n_916),
.B(n_600),
.C(n_601),
.Y(n_1184)
);

AOI21x1_ASAP7_75t_L g1185 ( 
.A1(n_954),
.A2(n_915),
.B(n_914),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_951),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_940),
.B(n_890),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_940),
.B(n_890),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_940),
.B(n_890),
.Y(n_1189)
);

AO32x2_ASAP7_75t_L g1190 ( 
.A1(n_1034),
.A2(n_1056),
.A3(n_997),
.B1(n_985),
.B2(n_994),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_939),
.Y(n_1191)
);

BUFx10_ASAP7_75t_L g1192 ( 
.A(n_968),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_973),
.A2(n_742),
.B(n_727),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_940),
.B(n_890),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1005),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_940),
.B(n_890),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_953),
.A2(n_1058),
.B(n_949),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_973),
.A2(n_742),
.B(n_727),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_940),
.B(n_600),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1000),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_944),
.A2(n_888),
.B(n_916),
.C(n_601),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_953),
.A2(n_1058),
.B(n_949),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_960),
.A2(n_1076),
.A3(n_1056),
.B(n_930),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_973),
.A2(n_742),
.B(n_727),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1005),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_973),
.A2(n_742),
.B(n_727),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_953),
.A2(n_1058),
.B(n_949),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_951),
.B(n_888),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1104),
.B(n_1105),
.Y(n_1209)
);

INVxp67_ASAP7_75t_SL g1210 ( 
.A(n_1098),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1132),
.A2(n_1113),
.B(n_1137),
.Y(n_1211)
);

OA21x2_ASAP7_75t_L g1212 ( 
.A1(n_1100),
.A2(n_1102),
.B(n_1099),
.Y(n_1212)
);

INVxp67_ASAP7_75t_L g1213 ( 
.A(n_1186),
.Y(n_1213)
);

NAND2x1p5_ASAP7_75t_L g1214 ( 
.A(n_1120),
.B(n_1159),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1187),
.B(n_1188),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1089),
.A2(n_1197),
.B(n_1182),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1180),
.A2(n_1199),
.B1(n_1154),
.B2(n_1208),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1183),
.A2(n_1184),
.B(n_1201),
.C(n_1157),
.Y(n_1218)
);

AO21x2_ASAP7_75t_L g1219 ( 
.A1(n_1100),
.A2(n_1099),
.B(n_1144),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1202),
.A2(n_1207),
.B(n_1133),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_1096),
.A2(n_1121),
.A3(n_1078),
.B(n_1116),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1081),
.Y(n_1222)
);

INVx1_ASAP7_75t_SL g1223 ( 
.A(n_1103),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1154),
.A2(n_1167),
.B1(n_1093),
.B2(n_1080),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1108),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1125),
.B(n_1165),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1149),
.A2(n_1142),
.B(n_1111),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1150),
.A2(n_1148),
.B(n_1153),
.C(n_1144),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1095),
.A2(n_1206),
.B(n_1204),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1193),
.A2(n_1198),
.B(n_1128),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1189),
.B(n_1194),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1150),
.A2(n_1164),
.B(n_1088),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1181),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1087),
.A2(n_1152),
.B(n_1106),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1097),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1085),
.B(n_1147),
.Y(n_1236)
);

AOI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1084),
.A2(n_1185),
.B(n_1090),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1145),
.A2(n_1196),
.B(n_1079),
.C(n_1151),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1086),
.B(n_1145),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1118),
.A2(n_1119),
.B(n_1135),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1123),
.A2(n_1126),
.B(n_1107),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1120),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1131),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_SL g1244 ( 
.A1(n_1158),
.A2(n_1176),
.B(n_1083),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1163),
.A2(n_1160),
.B(n_1171),
.Y(n_1245)
);

INVxp67_ASAP7_75t_SL g1246 ( 
.A(n_1122),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1114),
.A2(n_1161),
.B(n_1129),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1114),
.A2(n_1161),
.B(n_1129),
.Y(n_1248)
);

OR2x6_ASAP7_75t_L g1249 ( 
.A(n_1130),
.B(n_1139),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1138),
.A2(n_1172),
.B(n_1173),
.Y(n_1250)
);

INVx8_ASAP7_75t_L g1251 ( 
.A(n_1200),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1139),
.A2(n_1123),
.B(n_1101),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1110),
.A2(n_1112),
.B(n_1141),
.C(n_1191),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1109),
.A2(n_1127),
.B(n_1155),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1143),
.Y(n_1255)
);

O2A1O1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1147),
.A2(n_1162),
.B(n_1168),
.C(n_1177),
.Y(n_1256)
);

O2A1O1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1168),
.A2(n_1178),
.B(n_1092),
.C(n_1156),
.Y(n_1257)
);

OAI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1170),
.A2(n_1205),
.B1(n_1195),
.B2(n_1094),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1092),
.A2(n_1166),
.B(n_1190),
.C(n_1115),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1134),
.B(n_1170),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1179),
.B(n_1082),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1174),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1117),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1082),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1192),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1179),
.B(n_1109),
.Y(n_1266)
);

INVx2_ASAP7_75t_SL g1267 ( 
.A(n_1192),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_SL g1268 ( 
.A1(n_1190),
.A2(n_1179),
.B1(n_1146),
.B2(n_1203),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1200),
.B(n_1091),
.Y(n_1269)
);

INVx5_ASAP7_75t_L g1270 ( 
.A(n_1175),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1091),
.A2(n_1124),
.B(n_1136),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1140),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1190),
.A2(n_1203),
.B(n_1146),
.Y(n_1273)
);

INVx1_ASAP7_75t_SL g1274 ( 
.A(n_1117),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1169),
.B(n_1203),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1169),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1146),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1136),
.A2(n_1132),
.B(n_1113),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1169),
.A2(n_1100),
.B(n_1099),
.Y(n_1279)
);

NOR2xp67_ASAP7_75t_L g1280 ( 
.A(n_1097),
.B(n_793),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1132),
.A2(n_1113),
.B(n_1137),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1104),
.B(n_1105),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1193),
.A2(n_1204),
.B(n_1198),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1180),
.A2(n_944),
.B1(n_888),
.B2(n_945),
.Y(n_1284)
);

AOI32xp33_ASAP7_75t_L g1285 ( 
.A1(n_1199),
.A2(n_600),
.A3(n_489),
.B1(n_888),
.B2(n_1050),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1132),
.A2(n_1113),
.B(n_1137),
.Y(n_1286)
);

OAI222xp33_ASAP7_75t_L g1287 ( 
.A1(n_1154),
.A2(n_888),
.B1(n_1034),
.B2(n_945),
.C1(n_1021),
.C2(n_1183),
.Y(n_1287)
);

NOR2xp67_ASAP7_75t_L g1288 ( 
.A(n_1097),
.B(n_793),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1201),
.A2(n_1184),
.B(n_1183),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1199),
.B(n_321),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_1103),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1132),
.A2(n_1113),
.B(n_1137),
.Y(n_1292)
);

OA21x2_ASAP7_75t_L g1293 ( 
.A1(n_1100),
.A2(n_1102),
.B(n_1099),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1199),
.A2(n_888),
.B1(n_600),
.B2(n_770),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1181),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1106),
.B(n_1201),
.Y(n_1296)
);

O2A1O1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1180),
.A2(n_1201),
.B(n_916),
.C(n_1184),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_SL g1298 ( 
.A1(n_1199),
.A2(n_1050),
.B1(n_600),
.B2(n_618),
.Y(n_1298)
);

INVx3_ASAP7_75t_SL g1299 ( 
.A(n_1094),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1181),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1097),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1098),
.Y(n_1302)
);

AOI221xp5_ASAP7_75t_L g1303 ( 
.A1(n_1199),
.A2(n_600),
.B1(n_1180),
.B2(n_770),
.C(n_1145),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1201),
.A2(n_1184),
.B(n_1183),
.Y(n_1304)
);

AO32x2_ASAP7_75t_L g1305 ( 
.A1(n_1154),
.A2(n_1034),
.A3(n_1056),
.B1(n_997),
.B2(n_994),
.Y(n_1305)
);

NAND2x1p5_ASAP7_75t_L g1306 ( 
.A(n_1120),
.B(n_863),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1102),
.A2(n_1201),
.A3(n_960),
.B(n_1096),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_SL g1308 ( 
.A1(n_1158),
.A2(n_1184),
.B(n_1183),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1201),
.A2(n_1184),
.B(n_1183),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1180),
.A2(n_944),
.B1(n_888),
.B2(n_945),
.Y(n_1310)
);

OA21x2_ASAP7_75t_L g1311 ( 
.A1(n_1100),
.A2(n_1102),
.B(n_1099),
.Y(n_1311)
);

AOI221xp5_ASAP7_75t_L g1312 ( 
.A1(n_1199),
.A2(n_600),
.B1(n_1180),
.B2(n_770),
.C(n_1145),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1132),
.A2(n_1113),
.B(n_1137),
.Y(n_1313)
);

OAI221xp5_ASAP7_75t_L g1314 ( 
.A1(n_1201),
.A2(n_888),
.B1(n_600),
.B2(n_944),
.C(n_1180),
.Y(n_1314)
);

INVx4_ASAP7_75t_L g1315 ( 
.A(n_1120),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1180),
.A2(n_770),
.B1(n_600),
.B2(n_888),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1199),
.A2(n_888),
.B1(n_600),
.B2(n_770),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_SL g1318 ( 
.A1(n_1158),
.A2(n_1184),
.B(n_1183),
.Y(n_1318)
);

OAI222xp33_ASAP7_75t_L g1319 ( 
.A1(n_1154),
.A2(n_888),
.B1(n_1034),
.B2(n_945),
.C1(n_1021),
.C2(n_1183),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1180),
.A2(n_944),
.B1(n_888),
.B2(n_945),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_SL g1321 ( 
.A1(n_1201),
.A2(n_916),
.B(n_1180),
.C(n_1157),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1132),
.A2(n_1113),
.B(n_1137),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1104),
.B(n_1105),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1193),
.A2(n_1204),
.B(n_1198),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1236),
.B(n_1226),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1234),
.A2(n_1219),
.B(n_1232),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1215),
.B(n_1231),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1298),
.A2(n_1316),
.B1(n_1317),
.B2(n_1294),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1233),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1223),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1298),
.A2(n_1294),
.B1(n_1317),
.B2(n_1217),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1285),
.A2(n_1284),
.B1(n_1310),
.B2(n_1320),
.Y(n_1332)
);

O2A1O1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1287),
.A2(n_1319),
.B(n_1314),
.C(n_1218),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1303),
.B(n_1312),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1303),
.B(n_1312),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1210),
.B(n_1302),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1210),
.B(n_1302),
.Y(n_1337)
);

O2A1O1Ixp5_ASAP7_75t_L g1338 ( 
.A1(n_1287),
.A2(n_1319),
.B(n_1289),
.C(n_1304),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1314),
.A2(n_1224),
.B1(n_1290),
.B2(n_1280),
.Y(n_1339)
);

O2A1O1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1321),
.A2(n_1289),
.B(n_1309),
.C(n_1304),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1291),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1297),
.A2(n_1309),
.B(n_1228),
.C(n_1232),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1238),
.B(n_1291),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_SL g1344 ( 
.A1(n_1257),
.A2(n_1297),
.B(n_1296),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1241),
.A2(n_1240),
.B(n_1248),
.Y(n_1345)
);

AOI21x1_ASAP7_75t_SL g1346 ( 
.A1(n_1239),
.A2(n_1266),
.B(n_1296),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1238),
.B(n_1213),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1225),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1288),
.A2(n_1260),
.B1(n_1214),
.B2(n_1258),
.Y(n_1349)
);

A2O1A1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1241),
.A2(n_1253),
.B(n_1256),
.C(n_1257),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1253),
.A2(n_1256),
.B(n_1259),
.C(n_1252),
.Y(n_1351)
);

O2A1O1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1308),
.A2(n_1318),
.B(n_1259),
.C(n_1213),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1234),
.A2(n_1219),
.B(n_1283),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1283),
.A2(n_1324),
.B(n_1212),
.Y(n_1354)
);

O2A1O1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1252),
.A2(n_1214),
.B(n_1254),
.C(n_1244),
.Y(n_1355)
);

BUFx4f_ASAP7_75t_SL g1356 ( 
.A(n_1299),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1235),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1262),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1265),
.A2(n_1300),
.B1(n_1295),
.B2(n_1243),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1251),
.Y(n_1360)
);

AND2x2_ASAP7_75t_SL g1361 ( 
.A(n_1212),
.B(n_1293),
.Y(n_1361)
);

O2A1O1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1254),
.A2(n_1277),
.B(n_1255),
.C(n_1276),
.Y(n_1362)
);

AOI21x1_ASAP7_75t_SL g1363 ( 
.A1(n_1266),
.A2(n_1275),
.B(n_1269),
.Y(n_1363)
);

AOI21x1_ASAP7_75t_SL g1364 ( 
.A1(n_1269),
.A2(n_1305),
.B(n_1323),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1209),
.B(n_1282),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1301),
.Y(n_1366)
);

OR2x2_ASAP7_75t_SL g1367 ( 
.A(n_1242),
.B(n_1311),
.Y(n_1367)
);

AOI21x1_ASAP7_75t_SL g1368 ( 
.A1(n_1305),
.A2(n_1323),
.B(n_1282),
.Y(n_1368)
);

O2A1O1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1273),
.A2(n_1249),
.B(n_1279),
.C(n_1311),
.Y(n_1369)
);

O2A1O1Ixp5_ASAP7_75t_L g1370 ( 
.A1(n_1237),
.A2(n_1273),
.B(n_1324),
.C(n_1263),
.Y(n_1370)
);

A2O1A1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1271),
.A2(n_1268),
.B(n_1305),
.C(n_1270),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1279),
.A2(n_1293),
.B(n_1274),
.C(n_1272),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1251),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1270),
.A2(n_1268),
.B1(n_1315),
.B2(n_1242),
.Y(n_1374)
);

AOI21x1_ASAP7_75t_SL g1375 ( 
.A1(n_1307),
.A2(n_1270),
.B(n_1221),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_1251),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1274),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1247),
.A2(n_1278),
.B(n_1230),
.Y(n_1378)
);

AOI21x1_ASAP7_75t_SL g1379 ( 
.A1(n_1307),
.A2(n_1221),
.B(n_1250),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1307),
.B(n_1315),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1227),
.A2(n_1229),
.B(n_1322),
.Y(n_1381)
);

O2A1O1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1306),
.A2(n_1245),
.B(n_1281),
.C(n_1211),
.Y(n_1382)
);

AOI221xp5_ASAP7_75t_L g1383 ( 
.A1(n_1286),
.A2(n_1292),
.B1(n_1313),
.B2(n_1220),
.C(n_1216),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1298),
.A2(n_1316),
.B1(n_1317),
.B2(n_1294),
.Y(n_1384)
);

NOR2xp67_ASAP7_75t_L g1385 ( 
.A(n_1267),
.B(n_1264),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1232),
.A2(n_1241),
.B(n_1240),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1314),
.A2(n_1157),
.B(n_1183),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1298),
.A2(n_1316),
.B1(n_1317),
.B2(n_1294),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1242),
.Y(n_1389)
);

OA21x2_ASAP7_75t_L g1390 ( 
.A1(n_1232),
.A2(n_1241),
.B(n_1240),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1215),
.B(n_1231),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1236),
.B(n_1246),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1236),
.B(n_1226),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1234),
.A2(n_1100),
.B(n_1193),
.Y(n_1394)
);

O2A1O1Ixp5_ASAP7_75t_L g1395 ( 
.A1(n_1294),
.A2(n_1317),
.B(n_1232),
.C(n_1304),
.Y(n_1395)
);

AOI21x1_ASAP7_75t_SL g1396 ( 
.A1(n_1239),
.A2(n_1266),
.B(n_1261),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1236),
.B(n_1226),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1236),
.B(n_1246),
.Y(n_1398)
);

O2A1O1Ixp5_ASAP7_75t_L g1399 ( 
.A1(n_1294),
.A2(n_1317),
.B(n_1319),
.C(n_1287),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1222),
.Y(n_1400)
);

O2A1O1Ixp5_ASAP7_75t_L g1401 ( 
.A1(n_1294),
.A2(n_1317),
.B(n_1319),
.C(n_1287),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1354),
.A2(n_1326),
.B(n_1353),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1361),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1354),
.A2(n_1326),
.B(n_1353),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1399),
.A2(n_1401),
.B(n_1338),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1380),
.B(n_1371),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1347),
.B(n_1343),
.Y(n_1407)
);

AOI211xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1328),
.A2(n_1388),
.B(n_1384),
.C(n_1331),
.Y(n_1408)
);

OA21x2_ASAP7_75t_L g1409 ( 
.A1(n_1370),
.A2(n_1395),
.B(n_1394),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1336),
.B(n_1337),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1395),
.A2(n_1333),
.B(n_1387),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1377),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1378),
.Y(n_1413)
);

NAND4xp25_ASAP7_75t_L g1414 ( 
.A(n_1340),
.B(n_1333),
.C(n_1335),
.D(n_1334),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1394),
.A2(n_1340),
.B(n_1342),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1367),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1400),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1366),
.B(n_1348),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1345),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1362),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_1356),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1362),
.Y(n_1422)
);

AO21x2_ASAP7_75t_L g1423 ( 
.A1(n_1381),
.A2(n_1351),
.B(n_1372),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1369),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1392),
.B(n_1398),
.Y(n_1425)
);

OR2x6_ASAP7_75t_L g1426 ( 
.A(n_1369),
.B(n_1344),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1386),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1329),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1383),
.A2(n_1350),
.B(n_1374),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1386),
.B(n_1390),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1390),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1372),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1325),
.B(n_1393),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1355),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1382),
.Y(n_1435)
);

BUFx8_ASAP7_75t_SL g1436 ( 
.A(n_1357),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1382),
.Y(n_1437)
);

AO21x2_ASAP7_75t_L g1438 ( 
.A1(n_1352),
.A2(n_1332),
.B(n_1379),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1341),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1330),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1352),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1327),
.B(n_1391),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1412),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1430),
.B(n_1397),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1430),
.B(n_1375),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1417),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1413),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1413),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1427),
.B(n_1402),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1427),
.B(n_1368),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1412),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1439),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1414),
.A2(n_1339),
.B1(n_1349),
.B2(n_1365),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1416),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1406),
.B(n_1396),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1406),
.B(n_1396),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1413),
.Y(n_1457)
);

OAI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1408),
.A2(n_1359),
.B1(n_1358),
.B2(n_1385),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1402),
.B(n_1368),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1402),
.B(n_1404),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1411),
.A2(n_1389),
.B1(n_1360),
.B2(n_1376),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1431),
.B(n_1409),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1409),
.B(n_1364),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1411),
.A2(n_1389),
.B1(n_1373),
.B2(n_1346),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1402),
.B(n_1363),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1445),
.B(n_1403),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1453),
.A2(n_1415),
.B1(n_1407),
.B2(n_1426),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1446),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1446),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1445),
.B(n_1403),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1445),
.B(n_1403),
.Y(n_1471)
);

OAI31xp33_ASAP7_75t_SL g1472 ( 
.A1(n_1458),
.A2(n_1405),
.A3(n_1408),
.B(n_1441),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1443),
.B(n_1432),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1447),
.Y(n_1474)
);

OAI221xp5_ASAP7_75t_SL g1475 ( 
.A1(n_1453),
.A2(n_1415),
.B1(n_1407),
.B2(n_1426),
.C(n_1432),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1458),
.A2(n_1405),
.B1(n_1426),
.B2(n_1438),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1444),
.B(n_1403),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1464),
.A2(n_1438),
.B1(n_1441),
.B2(n_1434),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1460),
.A2(n_1449),
.B(n_1462),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1449),
.B(n_1463),
.Y(n_1480)
);

OAI31xp33_ASAP7_75t_SL g1481 ( 
.A1(n_1455),
.A2(n_1456),
.A3(n_1450),
.B(n_1424),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1449),
.B(n_1423),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_R g1483 ( 
.A(n_1464),
.B(n_1421),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1455),
.A2(n_1438),
.B1(n_1429),
.B2(n_1423),
.Y(n_1484)
);

AOI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1460),
.A2(n_1419),
.B(n_1437),
.Y(n_1485)
);

AO21x2_ASAP7_75t_L g1486 ( 
.A1(n_1460),
.A2(n_1423),
.B(n_1435),
.Y(n_1486)
);

INVxp67_ASAP7_75t_R g1487 ( 
.A(n_1465),
.Y(n_1487)
);

NAND3xp33_ASAP7_75t_L g1488 ( 
.A(n_1461),
.B(n_1409),
.C(n_1422),
.Y(n_1488)
);

OAI31xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1455),
.A2(n_1422),
.A3(n_1420),
.B(n_1425),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1452),
.Y(n_1490)
);

AO21x2_ASAP7_75t_L g1491 ( 
.A1(n_1460),
.A2(n_1423),
.B(n_1435),
.Y(n_1491)
);

AOI221xp5_ASAP7_75t_L g1492 ( 
.A1(n_1456),
.A2(n_1420),
.B1(n_1410),
.B2(n_1442),
.C(n_1440),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1479),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1479),
.Y(n_1494)
);

AO21x2_ASAP7_75t_L g1495 ( 
.A1(n_1486),
.A2(n_1491),
.B(n_1488),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1479),
.B(n_1462),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_SL g1497 ( 
.A(n_1483),
.B(n_1461),
.C(n_1452),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1469),
.Y(n_1498)
);

INVxp67_ASAP7_75t_L g1499 ( 
.A(n_1473),
.Y(n_1499)
);

OA21x2_ASAP7_75t_L g1500 ( 
.A1(n_1484),
.A2(n_1465),
.B(n_1459),
.Y(n_1500)
);

AOI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1485),
.A2(n_1457),
.B(n_1448),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1469),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1468),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1479),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1479),
.B(n_1459),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1473),
.B(n_1443),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1479),
.B(n_1459),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1485),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1466),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1490),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1480),
.B(n_1463),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1490),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1468),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1482),
.B(n_1451),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1474),
.Y(n_1515)
);

BUFx5_ASAP7_75t_L g1516 ( 
.A(n_1482),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1503),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1503),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1509),
.B(n_1487),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1495),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1513),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1513),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1506),
.B(n_1482),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1499),
.B(n_1492),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1509),
.B(n_1480),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1509),
.B(n_1487),
.Y(n_1526)
);

INVx1_ASAP7_75t_SL g1527 ( 
.A(n_1510),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1499),
.B(n_1492),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1512),
.B(n_1489),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1512),
.B(n_1489),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1511),
.B(n_1487),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1512),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1498),
.Y(n_1533)
);

INVxp67_ASAP7_75t_SL g1534 ( 
.A(n_1512),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1510),
.B(n_1436),
.Y(n_1535)
);

INVx2_ASAP7_75t_SL g1536 ( 
.A(n_1498),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1498),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1506),
.B(n_1481),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1497),
.A2(n_1467),
.B1(n_1476),
.B2(n_1483),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1495),
.B(n_1480),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1501),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1506),
.B(n_1486),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1495),
.B(n_1466),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1511),
.B(n_1466),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1511),
.B(n_1516),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1500),
.Y(n_1546)
);

OAI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1497),
.A2(n_1467),
.B(n_1476),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1502),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1511),
.B(n_1470),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1516),
.B(n_1470),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1516),
.B(n_1470),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1516),
.B(n_1471),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1514),
.B(n_1418),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1501),
.Y(n_1554)
);

A2O1A1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1505),
.A2(n_1481),
.B(n_1472),
.C(n_1475),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1502),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1514),
.B(n_1433),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1514),
.B(n_1456),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1558),
.B(n_1500),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1527),
.Y(n_1560)
);

BUFx2_ASAP7_75t_R g1561 ( 
.A(n_1529),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1533),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1532),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1519),
.B(n_1505),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1519),
.B(n_1505),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1526),
.B(n_1505),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1526),
.B(n_1507),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1553),
.B(n_1471),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1533),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1537),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1537),
.Y(n_1571)
);

INVxp67_ASAP7_75t_SL g1572 ( 
.A(n_1530),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1548),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1548),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1534),
.B(n_1471),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1556),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1556),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1524),
.B(n_1500),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1539),
.B(n_1472),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1532),
.B(n_1477),
.Y(n_1580)
);

NOR2xp67_ASAP7_75t_SL g1581 ( 
.A(n_1547),
.B(n_1488),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1531),
.B(n_1507),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1517),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1517),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1536),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1535),
.B(n_1433),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1536),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1525),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1525),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1531),
.B(n_1507),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1528),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1557),
.B(n_1477),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1538),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1588),
.B(n_1544),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1569),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1588),
.B(n_1544),
.Y(n_1596)
);

INVxp67_ASAP7_75t_SL g1597 ( 
.A(n_1563),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1575),
.B(n_1580),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1589),
.B(n_1549),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1579),
.B(n_1555),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1578),
.B(n_1593),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1569),
.Y(n_1602)
);

NOR2x1_ASAP7_75t_L g1603 ( 
.A(n_1560),
.B(n_1518),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1591),
.B(n_1549),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1589),
.B(n_1585),
.Y(n_1605)
);

INVx3_ASAP7_75t_SL g1606 ( 
.A(n_1578),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1564),
.B(n_1525),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1570),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1568),
.B(n_1523),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1561),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1582),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1585),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1572),
.B(n_1525),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1581),
.B(n_1583),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1564),
.B(n_1550),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1565),
.B(n_1550),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1586),
.B(n_1551),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1570),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1597),
.B(n_1581),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1603),
.B(n_1584),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1600),
.B(n_1592),
.Y(n_1621)
);

OAI32xp33_ASAP7_75t_L g1622 ( 
.A1(n_1614),
.A2(n_1546),
.A3(n_1610),
.B1(n_1601),
.B2(n_1559),
.Y(n_1622)
);

AOI211xp5_ASAP7_75t_L g1623 ( 
.A1(n_1606),
.A2(n_1475),
.B(n_1559),
.C(n_1543),
.Y(n_1623)
);

O2A1O1Ixp33_ASAP7_75t_L g1624 ( 
.A1(n_1606),
.A2(n_1520),
.B(n_1587),
.C(n_1504),
.Y(n_1624)
);

AOI221xp5_ASAP7_75t_L g1625 ( 
.A1(n_1606),
.A2(n_1543),
.B1(n_1495),
.B2(n_1540),
.C(n_1520),
.Y(n_1625)
);

AOI221x1_ASAP7_75t_L g1626 ( 
.A1(n_1605),
.A2(n_1587),
.B1(n_1521),
.B2(n_1522),
.C(n_1518),
.Y(n_1626)
);

AOI21xp33_ASAP7_75t_L g1627 ( 
.A1(n_1601),
.A2(n_1495),
.B(n_1562),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1612),
.B(n_1582),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1613),
.B(n_1590),
.Y(n_1629)
);

INVxp67_ASAP7_75t_SL g1630 ( 
.A(n_1604),
.Y(n_1630)
);

AO21x1_ASAP7_75t_L g1631 ( 
.A1(n_1605),
.A2(n_1573),
.B(n_1571),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1595),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1617),
.A2(n_1495),
.B(n_1520),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1594),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1595),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1605),
.Y(n_1636)
);

CKINVDCx14_ASAP7_75t_R g1637 ( 
.A(n_1594),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1634),
.B(n_1637),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1636),
.B(n_1596),
.Y(n_1639)
);

BUFx12f_ASAP7_75t_L g1640 ( 
.A(n_1630),
.Y(n_1640)
);

INVxp67_ASAP7_75t_L g1641 ( 
.A(n_1619),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1621),
.B(n_1598),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1629),
.A2(n_1611),
.B1(n_1609),
.B2(n_1598),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1636),
.Y(n_1644)
);

NOR2x1_ASAP7_75t_L g1645 ( 
.A(n_1620),
.B(n_1602),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1628),
.B(n_1596),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1631),
.B(n_1609),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1626),
.B(n_1599),
.Y(n_1648)
);

OAI211xp5_ASAP7_75t_L g1649 ( 
.A1(n_1647),
.A2(n_1622),
.B(n_1623),
.C(n_1624),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1639),
.Y(n_1650)
);

OAI221xp5_ASAP7_75t_L g1651 ( 
.A1(n_1648),
.A2(n_1625),
.B1(n_1627),
.B2(n_1633),
.C(n_1611),
.Y(n_1651)
);

AOI211xp5_ASAP7_75t_L g1652 ( 
.A1(n_1642),
.A2(n_1635),
.B(n_1632),
.C(n_1608),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1640),
.Y(n_1653)
);

AOI21xp33_ASAP7_75t_L g1654 ( 
.A1(n_1638),
.A2(n_1608),
.B(n_1602),
.Y(n_1654)
);

AOI221xp5_ASAP7_75t_SL g1655 ( 
.A1(n_1641),
.A2(n_1618),
.B1(n_1599),
.B2(n_1607),
.C(n_1576),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1644),
.Y(n_1656)
);

AOI221xp5_ASAP7_75t_L g1657 ( 
.A1(n_1643),
.A2(n_1618),
.B1(n_1543),
.B2(n_1520),
.C(n_1540),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1646),
.A2(n_1645),
.B1(n_1607),
.B2(n_1616),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1648),
.A2(n_1577),
.B(n_1573),
.Y(n_1659)
);

A2O1A1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1649),
.A2(n_1504),
.B(n_1543),
.C(n_1521),
.Y(n_1660)
);

OAI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1658),
.A2(n_1574),
.B1(n_1571),
.B2(n_1478),
.C(n_1504),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1656),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1653),
.A2(n_1616),
.B1(n_1615),
.B2(n_1540),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1650),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1660),
.B(n_1655),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1664),
.Y(n_1666)
);

INVxp67_ASAP7_75t_SL g1667 ( 
.A(n_1662),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1663),
.B(n_1652),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1661),
.Y(n_1669)
);

INVxp33_ASAP7_75t_L g1670 ( 
.A(n_1663),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_R g1671 ( 
.A(n_1666),
.B(n_1654),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1670),
.B(n_1659),
.Y(n_1672)
);

NAND2xp33_ASAP7_75t_SL g1673 ( 
.A(n_1668),
.B(n_1615),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1667),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1665),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1674),
.Y(n_1676)
);

NOR4xp75_ASAP7_75t_L g1677 ( 
.A(n_1672),
.B(n_1651),
.C(n_1673),
.D(n_1671),
.Y(n_1677)
);

OAI211xp5_ASAP7_75t_SL g1678 ( 
.A1(n_1675),
.A2(n_1669),
.B(n_1657),
.C(n_1574),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1677),
.Y(n_1679)
);

OAI322xp33_ASAP7_75t_L g1680 ( 
.A1(n_1679),
.A2(n_1676),
.A3(n_1678),
.B1(n_1542),
.B2(n_1522),
.C1(n_1493),
.C2(n_1494),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1680),
.A2(n_1540),
.B1(n_1567),
.B2(n_1566),
.Y(n_1681)
);

OA22x2_ASAP7_75t_L g1682 ( 
.A1(n_1681),
.A2(n_1567),
.B1(n_1565),
.B2(n_1566),
.Y(n_1682)
);

AOI22x1_ASAP7_75t_L g1683 ( 
.A1(n_1682),
.A2(n_1590),
.B1(n_1554),
.B2(n_1541),
.Y(n_1683)
);

AOI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1683),
.A2(n_1545),
.B1(n_1541),
.B2(n_1554),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1683),
.A2(n_1545),
.B1(n_1541),
.B2(n_1554),
.Y(n_1685)
);

XNOR2xp5_ASAP7_75t_L g1686 ( 
.A(n_1684),
.B(n_1428),
.Y(n_1686)
);

AOI22x1_ASAP7_75t_L g1687 ( 
.A1(n_1685),
.A2(n_1542),
.B1(n_1551),
.B2(n_1552),
.Y(n_1687)
);

OAI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1686),
.A2(n_1552),
.B(n_1523),
.Y(n_1688)
);

AOI222xp33_ASAP7_75t_L g1689 ( 
.A1(n_1687),
.A2(n_1493),
.B1(n_1494),
.B2(n_1507),
.C1(n_1496),
.C2(n_1515),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1688),
.Y(n_1690)
);

AOI322xp5_ASAP7_75t_L g1691 ( 
.A1(n_1689),
.A2(n_1493),
.A3(n_1494),
.B1(n_1496),
.B2(n_1508),
.C1(n_1478),
.C2(n_1454),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1690),
.A2(n_1691),
.B1(n_1493),
.B2(n_1494),
.Y(n_1692)
);

AOI211xp5_ASAP7_75t_L g1693 ( 
.A1(n_1692),
.A2(n_1428),
.B(n_1508),
.C(n_1439),
.Y(n_1693)
);


endmodule