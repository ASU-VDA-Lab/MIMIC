module fake_jpeg_9302_n_141 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_13),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_37),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_3),
.Y(n_52)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_23),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_26),
.B1(n_27),
.B2(n_23),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_26),
.B1(n_23),
.B2(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_28),
.B1(n_16),
.B2(n_20),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_32),
.A2(n_36),
.B1(n_29),
.B2(n_20),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_67),
.Y(n_73)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

AO22x2_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_38),
.B1(n_30),
.B2(n_31),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_50),
.B1(n_43),
.B2(n_44),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_29),
.B1(n_16),
.B2(n_36),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_38),
.B1(n_30),
.B2(n_15),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_47),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_13),
.B1(n_22),
.B2(n_19),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_50),
.A2(n_15),
.B1(n_22),
.B2(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_30),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_17),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_43),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_51),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_82),
.B1(n_57),
.B2(n_72),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_77),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_52),
.C(n_31),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

AO21x1_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_83),
.B(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_45),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_3),
.Y(n_98)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_98),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_80),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_94),
.B1(n_72),
.B2(n_82),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_57),
.B1(n_56),
.B2(n_59),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_96),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_97),
.B(n_54),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_105),
.B1(n_98),
.B2(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_78),
.C(n_74),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_107),
.C(n_108),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_79),
.B1(n_81),
.B2(n_59),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_76),
.C(n_31),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_35),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_31),
.C(n_35),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_92),
.C(n_89),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_87),
.B1(n_94),
.B2(n_93),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_110),
.A2(n_109),
.B1(n_106),
.B2(n_95),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_115),
.Y(n_122)
);

XNOR2x1_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_92),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_114),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_SL g115 ( 
.A(n_107),
.B(n_21),
.C(n_6),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_70),
.B1(n_95),
.B2(n_55),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_119),
.B(n_124),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_84),
.B1(n_65),
.B2(n_46),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_123),
.A2(n_119),
.B(n_84),
.C(n_122),
.Y(n_129)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_117),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_126),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_117),
.C(n_112),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_113),
.B1(n_118),
.B2(n_115),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_129),
.B(n_35),
.C(n_6),
.Y(n_132)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_123),
.B(n_5),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_133),
.B1(n_129),
.B2(n_9),
.Y(n_135)
);

AOI31xp67_ASAP7_75t_SL g136 ( 
.A1(n_132),
.A2(n_10),
.A3(n_11),
.B(n_12),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_7),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_136),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_138),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_137),
.B(n_130),
.Y(n_140)
);

A2O1A1O1Ixp25_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_5),
.B(n_10),
.C(n_12),
.D(n_136),
.Y(n_141)
);


endmodule