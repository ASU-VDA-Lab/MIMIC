module fake_aes_2931_n_1423 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_137, n_277, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_241, n_95, n_238, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_210, n_184, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1423);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_241;
input n_95;
input n_238;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_210;
input n_184;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1423;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_311;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1209;
wire n_1399;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_315;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1204;
wire n_1094;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_1275;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_1410;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g310 ( .A(n_24), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_306), .Y(n_311) );
INVxp33_ASAP7_75t_L g312 ( .A(n_142), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_266), .Y(n_313) );
CKINVDCx16_ASAP7_75t_R g314 ( .A(n_203), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_134), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_309), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_191), .Y(n_317) );
INVx1_ASAP7_75t_SL g318 ( .A(n_44), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_12), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_250), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_123), .Y(n_321) );
CKINVDCx16_ASAP7_75t_R g322 ( .A(n_16), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_211), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_118), .Y(n_324) );
CKINVDCx14_ASAP7_75t_R g325 ( .A(n_132), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_26), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_269), .Y(n_327) );
INVxp33_ASAP7_75t_L g328 ( .A(n_110), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_258), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_73), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_174), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_200), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_244), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_46), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g335 ( .A(n_235), .Y(n_335) );
XNOR2xp5_ASAP7_75t_L g336 ( .A(n_14), .B(n_71), .Y(n_336) );
INVxp67_ASAP7_75t_SL g337 ( .A(n_229), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_238), .Y(n_338) );
INVxp67_ASAP7_75t_L g339 ( .A(n_95), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_181), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_242), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_165), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_97), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_225), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_278), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_13), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_62), .Y(n_347) );
INVxp33_ASAP7_75t_SL g348 ( .A(n_136), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_171), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_30), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_130), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_227), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_216), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_277), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_236), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_143), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_221), .Y(n_357) );
CKINVDCx16_ASAP7_75t_R g358 ( .A(n_100), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_257), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_103), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_220), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_98), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_63), .Y(n_363) );
INVxp67_ASAP7_75t_SL g364 ( .A(n_276), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_148), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_74), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_232), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_27), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_215), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_82), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_187), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_146), .Y(n_372) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_153), .Y(n_373) );
INVxp33_ASAP7_75t_SL g374 ( .A(n_89), .Y(n_374) );
INVxp33_ASAP7_75t_L g375 ( .A(n_296), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_268), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_264), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_27), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_297), .Y(n_379) );
NOR2xp67_ASAP7_75t_L g380 ( .A(n_152), .B(n_1), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_265), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_111), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_80), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_169), .Y(n_384) );
BUFx5_ASAP7_75t_L g385 ( .A(n_49), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_53), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_199), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_254), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_68), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_19), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_156), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_209), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_12), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_18), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_57), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_303), .Y(n_396) );
INVxp67_ASAP7_75t_SL g397 ( .A(n_50), .Y(n_397) );
INVx2_ASAP7_75t_SL g398 ( .A(n_15), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_263), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_124), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_139), .Y(n_401) );
CKINVDCx16_ASAP7_75t_R g402 ( .A(n_73), .Y(n_402) );
INVxp67_ASAP7_75t_L g403 ( .A(n_275), .Y(n_403) );
INVxp33_ASAP7_75t_L g404 ( .A(n_289), .Y(n_404) );
BUFx3_ASAP7_75t_L g405 ( .A(n_157), .Y(n_405) );
INVxp33_ASAP7_75t_L g406 ( .A(n_70), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_39), .Y(n_407) );
CKINVDCx16_ASAP7_75t_R g408 ( .A(n_32), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_128), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_149), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_137), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_202), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_24), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_219), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_92), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_271), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_55), .Y(n_417) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_167), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_300), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_104), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_57), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_29), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_164), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_288), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_114), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_180), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_150), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_284), .Y(n_428) );
BUFx2_ASAP7_75t_L g429 ( .A(n_231), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_48), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_281), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_75), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_106), .Y(n_433) );
CKINVDCx16_ASAP7_75t_R g434 ( .A(n_293), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_183), .Y(n_435) );
BUFx3_ASAP7_75t_L g436 ( .A(n_64), .Y(n_436) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_1), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_129), .Y(n_438) );
INVxp33_ASAP7_75t_SL g439 ( .A(n_54), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_10), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_120), .Y(n_441) );
INVxp33_ASAP7_75t_SL g442 ( .A(n_96), .Y(n_442) );
INVxp67_ASAP7_75t_SL g443 ( .A(n_255), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_198), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_305), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_194), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_144), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_50), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_260), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_112), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_102), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_154), .Y(n_452) );
CKINVDCx16_ASAP7_75t_R g453 ( .A(n_179), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_90), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_173), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_5), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_47), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_140), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_273), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_240), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_272), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_245), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_42), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_349), .Y(n_464) );
INVx2_ASAP7_75t_SL g465 ( .A(n_321), .Y(n_465) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_349), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_385), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_406), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_314), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_349), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_385), .Y(n_471) );
BUFx2_ASAP7_75t_L g472 ( .A(n_389), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_322), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_385), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_398), .B(n_0), .Y(n_475) );
NAND2xp33_ASAP7_75t_SL g476 ( .A(n_406), .B(n_0), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_358), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_312), .B(n_2), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_385), .Y(n_479) );
INVx4_ASAP7_75t_L g480 ( .A(n_429), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_349), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_434), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_385), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_418), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_385), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_385), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_312), .B(n_2), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_366), .B(n_3), .Y(n_488) );
AOI22xp33_ASAP7_75t_SL g489 ( .A1(n_319), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_366), .Y(n_490) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_418), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_402), .Y(n_492) );
BUFx2_ASAP7_75t_L g493 ( .A(n_389), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_328), .B(n_4), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_418), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_413), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_408), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_413), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_461), .B(n_6), .Y(n_499) );
AND2x6_ASAP7_75t_L g500 ( .A(n_488), .B(n_405), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_488), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_480), .B(n_465), .Y(n_502) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_466), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_480), .B(n_328), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_488), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_480), .B(n_375), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_488), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_468), .B(n_390), .Y(n_508) );
OR2x2_ASAP7_75t_SL g509 ( .A(n_468), .B(n_453), .Y(n_509) );
BUFx2_ASAP7_75t_L g510 ( .A(n_469), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_472), .B(n_436), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_488), .Y(n_512) );
NAND3x1_ASAP7_75t_L g513 ( .A(n_478), .B(n_346), .C(n_310), .Y(n_513) );
NOR2xp33_ASAP7_75t_SL g514 ( .A(n_478), .B(n_332), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_480), .B(n_375), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_465), .A2(n_439), .B1(n_335), .B2(n_381), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_478), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_472), .B(n_318), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_477), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_485), .Y(n_520) );
INVx2_ASAP7_75t_SL g521 ( .A(n_487), .Y(n_521) );
AND2x6_ASAP7_75t_L g522 ( .A(n_487), .B(n_405), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_487), .Y(n_523) );
BUFx2_ASAP7_75t_L g524 ( .A(n_482), .Y(n_524) );
CKINVDCx16_ASAP7_75t_R g525 ( .A(n_473), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_485), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_494), .Y(n_527) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_466), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_493), .B(n_404), .Y(n_529) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_466), .Y(n_530) );
AND2x6_ASAP7_75t_L g531 ( .A(n_494), .B(n_313), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_493), .B(n_404), .Y(n_532) );
OR2x6_ASAP7_75t_L g533 ( .A(n_494), .B(n_422), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_475), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_492), .Y(n_535) );
INVx4_ASAP7_75t_L g536 ( .A(n_485), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_499), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_497), .Y(n_538) );
INVx3_ASAP7_75t_L g539 ( .A(n_485), .Y(n_539) );
NOR2xp33_ASAP7_75t_SL g540 ( .A(n_499), .B(n_332), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_465), .B(n_325), .Y(n_541) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_466), .Y(n_542) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_466), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_490), .B(n_325), .Y(n_544) );
BUFx3_ASAP7_75t_L g545 ( .A(n_467), .Y(n_545) );
AO22x2_ASAP7_75t_L g546 ( .A1(n_475), .A2(n_437), .B1(n_397), .B2(n_422), .Y(n_546) );
NOR2xp33_ASAP7_75t_R g547 ( .A(n_514), .B(n_335), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_539), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_539), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_534), .B(n_348), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_515), .B(n_348), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_539), .Y(n_552) );
INVx3_ASAP7_75t_L g553 ( .A(n_500), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_515), .B(n_374), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_537), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_529), .B(n_334), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_521), .Y(n_557) );
BUFx2_ASAP7_75t_L g558 ( .A(n_518), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_541), .B(n_374), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_504), .B(n_442), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_521), .Y(n_561) );
AND2x6_ASAP7_75t_L g562 ( .A(n_501), .B(n_311), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_533), .B(n_381), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_513), .A2(n_476), .B1(n_439), .B2(n_384), .Y(n_564) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_505), .A2(n_471), .B(n_467), .Y(n_565) );
NOR2x1p5_ASAP7_75t_L g566 ( .A(n_518), .B(n_368), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_506), .B(n_442), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_546), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_502), .B(n_490), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_507), .Y(n_570) );
AOI21xp33_ASAP7_75t_L g571 ( .A1(n_502), .A2(n_364), .B(n_337), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_512), .A2(n_474), .B(n_471), .Y(n_572) );
A2O1A1Ixp33_ASAP7_75t_L g573 ( .A1(n_517), .A2(n_474), .B(n_483), .C(n_479), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_546), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_546), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_523), .B(n_496), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_532), .B(n_529), .Y(n_577) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_500), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_533), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_508), .B(n_386), .Y(n_580) );
A2O1A1Ixp33_ASAP7_75t_L g581 ( .A1(n_527), .A2(n_479), .B(n_486), .C(n_483), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_533), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_541), .B(n_486), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_511), .B(n_315), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_511), .B(n_496), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_533), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_511), .B(n_498), .Y(n_587) );
BUFx2_ASAP7_75t_L g588 ( .A(n_510), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_508), .B(n_320), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_520), .Y(n_590) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_500), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_531), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_531), .B(n_498), .Y(n_593) );
INVx5_ASAP7_75t_L g594 ( .A(n_500), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_531), .Y(n_595) );
INVxp67_ASAP7_75t_L g596 ( .A(n_531), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_531), .B(n_384), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_520), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_509), .A2(n_388), .B1(n_409), .B2(n_387), .Y(n_599) );
INVx2_ASAP7_75t_SL g600 ( .A(n_522), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_544), .B(n_339), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_526), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_540), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_513), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_526), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_500), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_535), .Y(n_607) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_500), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_536), .B(n_331), .Y(n_609) );
BUFx2_ASAP7_75t_L g610 ( .A(n_524), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_522), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_536), .B(n_338), .Y(n_612) );
BUFx4f_ASAP7_75t_SL g613 ( .A(n_538), .Y(n_613) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_522), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_536), .B(n_403), .Y(n_615) );
INVxp67_ASAP7_75t_L g616 ( .A(n_522), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_522), .B(n_344), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_545), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_519), .B(n_345), .Y(n_619) );
INVx5_ASAP7_75t_L g620 ( .A(n_503), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_545), .B(n_355), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_503), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_516), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g624 ( .A(n_503), .B(n_347), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g625 ( .A(n_538), .Y(n_625) );
INVx3_ASAP7_75t_L g626 ( .A(n_503), .Y(n_626) );
BUFx2_ASAP7_75t_L g627 ( .A(n_525), .Y(n_627) );
NOR3xp33_ASAP7_75t_SL g628 ( .A(n_528), .B(n_456), .C(n_407), .Y(n_628) );
NOR3xp33_ASAP7_75t_SL g629 ( .A(n_528), .B(n_336), .C(n_356), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_528), .B(n_360), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_528), .B(n_489), .Y(n_631) );
INVx5_ASAP7_75t_L g632 ( .A(n_530), .Y(n_632) );
AND2x4_ASAP7_75t_L g633 ( .A(n_543), .B(n_387), .Y(n_633) );
BUFx3_ASAP7_75t_L g634 ( .A(n_530), .Y(n_634) );
INVx2_ASAP7_75t_SL g635 ( .A(n_530), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_530), .Y(n_636) );
NOR2x1p5_ASAP7_75t_L g637 ( .A(n_542), .B(n_319), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_542), .B(n_316), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_577), .B(n_388), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_557), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_555), .B(n_409), .Y(n_641) );
NAND2x1p5_ASAP7_75t_L g642 ( .A(n_594), .B(n_436), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_580), .B(n_425), .Y(n_643) );
INVx4_ASAP7_75t_L g644 ( .A(n_594), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_548), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_558), .B(n_489), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_549), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_569), .B(n_425), .Y(n_648) );
OR2x6_ASAP7_75t_L g649 ( .A(n_563), .B(n_440), .Y(n_649) );
AOI21xp33_ASAP7_75t_L g650 ( .A1(n_631), .A2(n_443), .B(n_373), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_569), .B(n_433), .Y(n_651) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_578), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_568), .A2(n_462), .B1(n_433), .B2(n_330), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_572), .A2(n_323), .B(n_317), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_578), .B(n_462), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_607), .Y(n_656) );
BUFx3_ASAP7_75t_L g657 ( .A(n_588), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_633), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_552), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_572), .A2(n_327), .B(n_324), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_610), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_574), .A2(n_326), .B1(n_350), .B2(n_330), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_623), .A2(n_575), .B1(n_604), .B2(n_582), .Y(n_663) );
BUFx2_ASAP7_75t_SL g664 ( .A(n_563), .Y(n_664) );
INVx3_ASAP7_75t_L g665 ( .A(n_578), .Y(n_665) );
INVx3_ASAP7_75t_L g666 ( .A(n_578), .Y(n_666) );
BUFx2_ASAP7_75t_L g667 ( .A(n_547), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_583), .B(n_363), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_556), .B(n_326), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_570), .Y(n_670) );
INVx3_ASAP7_75t_L g671 ( .A(n_591), .Y(n_671) );
INVx3_ASAP7_75t_L g672 ( .A(n_591), .Y(n_672) );
BUFx12f_ASAP7_75t_L g673 ( .A(n_625), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_579), .A2(n_393), .B1(n_350), .B2(n_378), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_591), .B(n_370), .Y(n_675) );
AOI21xp33_ASAP7_75t_L g676 ( .A1(n_551), .A2(n_340), .B(n_329), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g677 ( .A1(n_576), .A2(n_581), .B(n_573), .C(n_585), .Y(n_677) );
INVx4_ASAP7_75t_L g678 ( .A(n_594), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_590), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_561), .Y(n_680) );
BUFx12f_ASAP7_75t_L g681 ( .A(n_627), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_576), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_550), .B(n_394), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_598), .Y(n_684) );
BUFx6f_ASAP7_75t_L g685 ( .A(n_591), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_594), .B(n_379), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_593), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_585), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_597), .B(n_393), .Y(n_689) );
BUFx3_ASAP7_75t_L g690 ( .A(n_613), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_565), .A2(n_342), .B(n_341), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_602), .Y(n_692) );
CKINVDCx5p33_ASAP7_75t_R g693 ( .A(n_547), .Y(n_693) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_614), .Y(n_694) );
INVx4_ASAP7_75t_L g695 ( .A(n_614), .Y(n_695) );
INVx3_ASAP7_75t_SL g696 ( .A(n_633), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_587), .Y(n_697) );
O2A1O1Ixp33_ASAP7_75t_L g698 ( .A1(n_587), .A2(n_417), .B(n_421), .C(n_395), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_589), .B(n_559), .Y(n_699) );
NAND2x1_ASAP7_75t_SL g700 ( .A(n_597), .B(n_380), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_605), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_586), .A2(n_432), .B1(n_448), .B2(n_430), .Y(n_702) );
INVx8_ASAP7_75t_L g703 ( .A(n_614), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_566), .B(n_457), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_624), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_592), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_564), .A2(n_554), .B1(n_603), .B2(n_567), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_599), .B(n_463), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_624), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_562), .A2(n_440), .B1(n_351), .B2(n_354), .Y(n_710) );
INVx3_ASAP7_75t_L g711 ( .A(n_614), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_595), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_565), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_L g714 ( .A1(n_601), .A2(n_357), .B(n_359), .C(n_343), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_562), .B(n_361), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_618), .Y(n_716) );
NAND2xp5_ASAP7_75t_SL g717 ( .A(n_553), .B(n_383), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_560), .A2(n_365), .B(n_362), .Y(n_718) );
CKINVDCx5p33_ASAP7_75t_R g719 ( .A(n_613), .Y(n_719) );
INVx5_ASAP7_75t_L g720 ( .A(n_553), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_596), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_606), .Y(n_722) );
O2A1O1Ixp33_ASAP7_75t_L g723 ( .A1(n_571), .A2(n_369), .B(n_371), .C(n_367), .Y(n_723) );
INVx2_ASAP7_75t_SL g724 ( .A(n_637), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_615), .A2(n_377), .B(n_376), .Y(n_725) );
INVx1_ASAP7_75t_SL g726 ( .A(n_562), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_562), .B(n_382), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_584), .B(n_396), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_603), .B(n_401), .Y(n_729) );
INVx1_ASAP7_75t_SL g730 ( .A(n_562), .Y(n_730) );
O2A1O1Ixp33_ASAP7_75t_SL g731 ( .A1(n_611), .A2(n_392), .B(n_399), .C(n_391), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_596), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g733 ( .A1(n_601), .A2(n_410), .B(n_400), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_638), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_629), .B(n_6), .Y(n_735) );
OR2x6_ASAP7_75t_L g736 ( .A(n_600), .B(n_608), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_615), .A2(n_414), .B(n_412), .Y(n_737) );
INVx4_ASAP7_75t_L g738 ( .A(n_608), .Y(n_738) );
BUFx3_ASAP7_75t_L g739 ( .A(n_620), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_629), .B(n_7), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_616), .A2(n_419), .B1(n_420), .B2(n_415), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_638), .Y(n_742) );
INVx3_ASAP7_75t_L g743 ( .A(n_620), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_630), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_609), .A2(n_424), .B(n_423), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_621), .Y(n_746) );
A2O1A1Ixp33_ASAP7_75t_L g747 ( .A1(n_616), .A2(n_428), .B(n_431), .C(n_426), .Y(n_747) );
BUFx12f_ASAP7_75t_L g748 ( .A(n_620), .Y(n_748) );
AOI21xp5_ASAP7_75t_L g749 ( .A1(n_612), .A2(n_438), .B(n_435), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_628), .A2(n_444), .B1(n_446), .B2(n_441), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_634), .Y(n_751) );
BUFx6f_ASAP7_75t_L g752 ( .A(n_620), .Y(n_752) );
INVx3_ASAP7_75t_L g753 ( .A(n_632), .Y(n_753) );
INVx2_ASAP7_75t_SL g754 ( .A(n_619), .Y(n_754) );
O2A1O1Ixp33_ASAP7_75t_L g755 ( .A1(n_628), .A2(n_449), .B(n_450), .C(n_447), .Y(n_755) );
O2A1O1Ixp33_ASAP7_75t_SL g756 ( .A1(n_617), .A2(n_454), .B(n_455), .C(n_452), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_635), .B(n_458), .Y(n_757) );
O2A1O1Ixp33_ASAP7_75t_L g758 ( .A1(n_636), .A2(n_333), .B(n_352), .C(n_313), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_626), .B(n_411), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_622), .A2(n_352), .B(n_333), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_632), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_632), .B(n_7), .Y(n_762) );
AO21x2_ASAP7_75t_L g763 ( .A1(n_632), .A2(n_372), .B(n_353), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_626), .B(n_353), .Y(n_764) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_558), .Y(n_765) );
BUFx6f_ASAP7_75t_L g766 ( .A(n_578), .Y(n_766) );
BUFx2_ASAP7_75t_L g767 ( .A(n_588), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_613), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_548), .Y(n_769) );
OR2x2_ASAP7_75t_L g770 ( .A(n_607), .B(n_8), .Y(n_770) );
O2A1O1Ixp33_ASAP7_75t_L g771 ( .A1(n_568), .A2(n_416), .B(n_451), .C(n_372), .Y(n_771) );
BUFx12f_ASAP7_75t_L g772 ( .A(n_625), .Y(n_772) );
BUFx6f_ASAP7_75t_L g773 ( .A(n_578), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_577), .B(n_427), .Y(n_774) );
INVx1_ASAP7_75t_SL g775 ( .A(n_656), .Y(n_775) );
OA21x2_ASAP7_75t_L g776 ( .A1(n_691), .A2(n_451), .B(n_416), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_670), .Y(n_777) );
OA21x2_ASAP7_75t_L g778 ( .A1(n_691), .A2(n_460), .B(n_459), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_648), .B(n_445), .Y(n_779) );
NOR2xp67_ASAP7_75t_L g780 ( .A(n_661), .B(n_8), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_640), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_648), .B(n_9), .Y(n_782) );
OAI21xp5_ASAP7_75t_L g783 ( .A1(n_654), .A2(n_460), .B(n_459), .Y(n_783) );
AO31x2_ASAP7_75t_L g784 ( .A1(n_713), .A2(n_464), .A3(n_481), .B(n_470), .Y(n_784) );
INVx1_ASAP7_75t_SL g785 ( .A(n_767), .Y(n_785) );
OAI21x1_ASAP7_75t_L g786 ( .A1(n_760), .A2(n_470), .B(n_464), .Y(n_786) );
BUFx2_ASAP7_75t_SL g787 ( .A(n_657), .Y(n_787) );
NAND3xp33_ASAP7_75t_L g788 ( .A(n_755), .B(n_418), .C(n_464), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_679), .Y(n_789) );
INVx3_ASAP7_75t_L g790 ( .A(n_748), .Y(n_790) );
OR2x2_ASAP7_75t_L g791 ( .A(n_653), .B(n_9), .Y(n_791) );
INVxp67_ASAP7_75t_L g792 ( .A(n_765), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_680), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g794 ( .A1(n_725), .A2(n_543), .B(n_542), .Y(n_794) );
AOI22x1_ASAP7_75t_L g795 ( .A1(n_654), .A2(n_495), .B1(n_484), .B2(n_481), .Y(n_795) );
OAI21x1_ASAP7_75t_L g796 ( .A1(n_642), .A2(n_495), .B(n_484), .Y(n_796) );
NAND2x1p5_ASAP7_75t_L g797 ( .A(n_752), .B(n_484), .Y(n_797) );
CKINVDCx8_ASAP7_75t_R g798 ( .A(n_664), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_688), .A2(n_495), .B1(n_491), .B2(n_466), .Y(n_799) );
NAND3xp33_ASAP7_75t_L g800 ( .A(n_755), .B(n_491), .C(n_466), .Y(n_800) );
BUFx2_ASAP7_75t_L g801 ( .A(n_765), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_684), .Y(n_802) );
OR2x2_ASAP7_75t_L g803 ( .A(n_653), .B(n_10), .Y(n_803) );
AND2x4_ASAP7_75t_L g804 ( .A(n_682), .B(n_11), .Y(n_804) );
OR3x4_ASAP7_75t_SL g805 ( .A(n_768), .B(n_11), .C(n_13), .Y(n_805) );
INVx4_ASAP7_75t_L g806 ( .A(n_752), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_658), .Y(n_807) );
OAI21x1_ASAP7_75t_SL g808 ( .A1(n_677), .A2(n_14), .B(n_15), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_692), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_639), .B(n_16), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_701), .Y(n_811) );
NAND2x1p5_ASAP7_75t_L g812 ( .A(n_752), .B(n_491), .Y(n_812) );
OR2x2_ASAP7_75t_L g813 ( .A(n_662), .B(n_17), .Y(n_813) );
OAI21xp5_ASAP7_75t_L g814 ( .A1(n_660), .A2(n_491), .B(n_78), .Y(n_814) );
AOI21x1_ASAP7_75t_L g815 ( .A1(n_764), .A2(n_491), .B(n_542), .Y(n_815) );
BUFx2_ASAP7_75t_L g816 ( .A(n_681), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_651), .B(n_17), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_658), .Y(n_818) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_649), .Y(n_819) );
OAI21x1_ASAP7_75t_L g820 ( .A1(n_771), .A2(n_491), .B(n_543), .Y(n_820) );
OAI21x1_ASAP7_75t_L g821 ( .A1(n_771), .A2(n_491), .B(n_543), .Y(n_821) );
AOI211xp5_ASAP7_75t_L g822 ( .A1(n_643), .A2(n_18), .B(n_19), .C(n_20), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_646), .B(n_20), .Y(n_823) );
AND2x2_ASAP7_75t_L g824 ( .A(n_651), .B(n_21), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_697), .A2(n_21), .B1(n_22), .B2(n_23), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_649), .A2(n_22), .B1(n_23), .B2(n_25), .Y(n_826) );
INVx8_ASAP7_75t_L g827 ( .A(n_703), .Y(n_827) );
OA21x2_ASAP7_75t_L g828 ( .A1(n_660), .A2(n_79), .B(n_77), .Y(n_828) );
INVx3_ASAP7_75t_SL g829 ( .A(n_719), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_707), .B(n_25), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_716), .Y(n_831) );
OR2x2_ASAP7_75t_L g832 ( .A(n_662), .B(n_26), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_722), .Y(n_833) );
A2O1A1Ixp33_ASAP7_75t_L g834 ( .A1(n_677), .A2(n_28), .B(n_29), .C(n_30), .Y(n_834) );
OAI21x1_ASAP7_75t_L g835 ( .A1(n_642), .A2(n_83), .B(n_81), .Y(n_835) );
BUFx2_ASAP7_75t_L g836 ( .A(n_649), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_694), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_668), .Y(n_838) );
AO21x2_ASAP7_75t_L g839 ( .A1(n_763), .A2(n_85), .B(n_84), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_694), .Y(n_840) );
O2A1O1Ixp33_ASAP7_75t_SL g841 ( .A1(n_750), .A2(n_163), .B(n_307), .C(n_304), .Y(n_841) );
A2O1A1Ixp33_ASAP7_75t_L g842 ( .A1(n_723), .A2(n_28), .B(n_31), .C(n_32), .Y(n_842) );
OAI21x1_ASAP7_75t_L g843 ( .A1(n_764), .A2(n_87), .B(n_86), .Y(n_843) );
OAI21x1_ASAP7_75t_L g844 ( .A1(n_706), .A2(n_91), .B(n_88), .Y(n_844) );
INVx4_ASAP7_75t_L g845 ( .A(n_696), .Y(n_845) );
CKINVDCx5p33_ASAP7_75t_R g846 ( .A(n_673), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_694), .Y(n_847) );
A2O1A1Ixp33_ASAP7_75t_L g848 ( .A1(n_723), .A2(n_31), .B(n_33), .C(n_34), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_650), .A2(n_33), .B1(n_34), .B2(n_35), .Y(n_849) );
AO21x2_ASAP7_75t_L g850 ( .A1(n_763), .A2(n_94), .B(n_93), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_652), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_669), .B(n_35), .Y(n_852) );
AOI22x1_ASAP7_75t_L g853 ( .A1(n_725), .A2(n_175), .B1(n_302), .B2(n_301), .Y(n_853) );
NAND2x1p5_ASAP7_75t_L g854 ( .A(n_726), .B(n_36), .Y(n_854) );
BUFx2_ASAP7_75t_L g855 ( .A(n_696), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_668), .Y(n_856) );
OA21x2_ASAP7_75t_L g857 ( .A1(n_737), .A2(n_101), .B(n_99), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_652), .Y(n_858) );
AOI21xp33_ASAP7_75t_L g859 ( .A1(n_641), .A2(n_36), .B(n_37), .Y(n_859) );
OAI21x1_ASAP7_75t_L g860 ( .A1(n_758), .A2(n_107), .B(n_105), .Y(n_860) );
OAI21xp5_ASAP7_75t_L g861 ( .A1(n_737), .A2(n_109), .B(n_108), .Y(n_861) );
OAI21x1_ASAP7_75t_L g862 ( .A1(n_712), .A2(n_115), .B(n_113), .Y(n_862) );
OAI21x1_ASAP7_75t_L g863 ( .A1(n_705), .A2(n_117), .B(n_116), .Y(n_863) );
AO21x2_ASAP7_75t_L g864 ( .A1(n_731), .A2(n_121), .B(n_119), .Y(n_864) );
OAI21x1_ASAP7_75t_L g865 ( .A1(n_709), .A2(n_125), .B(n_122), .Y(n_865) );
AOI21xp33_ASAP7_75t_L g866 ( .A1(n_774), .A2(n_37), .B(n_38), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_730), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_867) );
AND2x4_ASAP7_75t_L g868 ( .A(n_746), .B(n_40), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_689), .B(n_41), .Y(n_869) );
NAND2x1p5_ASAP7_75t_L g870 ( .A(n_739), .B(n_41), .Y(n_870) );
OAI21xp5_ASAP7_75t_L g871 ( .A1(n_718), .A2(n_188), .B(n_299), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_683), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_652), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_683), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_708), .B(n_42), .Y(n_875) );
AND2x4_ASAP7_75t_L g876 ( .A(n_754), .B(n_43), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_663), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_770), .Y(n_878) );
OAI21x1_ASAP7_75t_L g879 ( .A1(n_757), .A2(n_189), .B(n_298), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_757), .Y(n_880) );
OAI21x1_ASAP7_75t_L g881 ( .A1(n_744), .A2(n_186), .B(n_295), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_650), .A2(n_45), .B1(n_46), .B2(n_47), .Y(n_882) );
OAI21x1_ASAP7_75t_L g883 ( .A1(n_743), .A2(n_192), .B(n_294), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_702), .Y(n_884) );
OAI21x1_ASAP7_75t_L g885 ( .A1(n_743), .A2(n_190), .B(n_292), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_733), .B(n_48), .Y(n_886) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_736), .Y(n_887) );
AOI21xp5_ASAP7_75t_L g888 ( .A1(n_718), .A2(n_185), .B(n_291), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_710), .A2(n_49), .B1(n_51), .B2(n_52), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_702), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_685), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_674), .B(n_51), .Y(n_892) );
AOI21xp5_ASAP7_75t_L g893 ( .A1(n_745), .A2(n_193), .B(n_290), .Y(n_893) );
AO21x2_ASAP7_75t_L g894 ( .A1(n_715), .A2(n_184), .B(n_287), .Y(n_894) );
CKINVDCx11_ASAP7_75t_R g895 ( .A(n_772), .Y(n_895) );
AOI21xp5_ASAP7_75t_L g896 ( .A1(n_745), .A2(n_182), .B(n_286), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_704), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_733), .B(n_52), .Y(n_898) );
OAI21x1_ASAP7_75t_L g899 ( .A1(n_758), .A2(n_195), .B(n_285), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_685), .Y(n_900) );
OAI21x1_ASAP7_75t_L g901 ( .A1(n_753), .A2(n_178), .B(n_283), .Y(n_901) );
NOR2x1_ASAP7_75t_R g902 ( .A(n_693), .B(n_53), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_714), .B(n_54), .Y(n_903) );
OAI21x1_ASAP7_75t_L g904 ( .A1(n_753), .A2(n_196), .B(n_282), .Y(n_904) );
NAND2xp5_ASAP7_75t_SL g905 ( .A(n_685), .B(n_126), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_676), .A2(n_55), .B1(n_56), .B2(n_58), .Y(n_906) );
CKINVDCx14_ASAP7_75t_R g907 ( .A(n_667), .Y(n_907) );
OAI21xp5_ASAP7_75t_L g908 ( .A1(n_687), .A2(n_197), .B(n_280), .Y(n_908) );
INVx2_ASAP7_75t_L g909 ( .A(n_766), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_735), .Y(n_910) );
NAND2x1p5_ASAP7_75t_L g911 ( .A(n_695), .B(n_56), .Y(n_911) );
INVx4_ASAP7_75t_SL g912 ( .A(n_766), .Y(n_912) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_736), .Y(n_913) );
AOI21x1_ASAP7_75t_L g914 ( .A1(n_715), .A2(n_177), .B(n_279), .Y(n_914) );
AOI22xp33_ASAP7_75t_SL g915 ( .A1(n_740), .A2(n_58), .B1(n_59), .B2(n_60), .Y(n_915) );
OAI22xp33_ASAP7_75t_L g916 ( .A1(n_724), .A2(n_59), .B1(n_60), .B2(n_61), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_645), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_698), .B(n_61), .Y(n_918) );
BUFx2_ASAP7_75t_L g919 ( .A(n_690), .Y(n_919) );
OAI21xp5_ASAP7_75t_L g920 ( .A1(n_742), .A2(n_204), .B(n_274), .Y(n_920) );
INVxp67_ASAP7_75t_L g921 ( .A(n_655), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_699), .B(n_62), .Y(n_922) );
CKINVDCx11_ASAP7_75t_R g923 ( .A(n_895), .Y(n_923) );
AOI21xp5_ASAP7_75t_L g924 ( .A1(n_794), .A2(n_749), .B(n_676), .Y(n_924) );
OAI22xp5_ASAP7_75t_SL g925 ( .A1(n_907), .A2(n_750), .B1(n_729), .B2(n_728), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_804), .A2(n_727), .B1(n_741), .B2(n_747), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_910), .A2(n_741), .B1(n_734), .B2(n_727), .Y(n_927) );
OAI22xp33_ASAP7_75t_L g928 ( .A1(n_791), .A2(n_736), .B1(n_738), .B2(n_766), .Y(n_928) );
CKINVDCx5p33_ASAP7_75t_R g929 ( .A(n_895), .Y(n_929) );
AOI21xp5_ASAP7_75t_L g930 ( .A1(n_838), .A2(n_749), .B(n_756), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g931 ( .A1(n_804), .A2(n_698), .B1(n_738), .B2(n_695), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_884), .A2(n_762), .B1(n_721), .B2(n_732), .Y(n_932) );
OA21x2_ASAP7_75t_L g933 ( .A1(n_820), .A2(n_700), .B(n_769), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_781), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_890), .B(n_647), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_856), .A2(n_659), .B1(n_720), .B2(n_761), .Y(n_936) );
CKINVDCx11_ASAP7_75t_R g937 ( .A(n_829), .Y(n_937) );
CKINVDCx5p33_ASAP7_75t_R g938 ( .A(n_846), .Y(n_938) );
NAND2xp33_ASAP7_75t_R g939 ( .A(n_846), .B(n_665), .Y(n_939) );
OAI221xp5_ASAP7_75t_L g940 ( .A1(n_872), .A2(n_717), .B1(n_759), .B2(n_675), .C(n_686), .Y(n_940) );
A2O1A1Ixp33_ASAP7_75t_L g941 ( .A1(n_817), .A2(n_666), .B(n_671), .C(n_672), .Y(n_941) );
OR2x2_ASAP7_75t_L g942 ( .A(n_775), .B(n_63), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g943 ( .A1(n_803), .A2(n_773), .B1(n_703), .B2(n_720), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_874), .A2(n_720), .B1(n_666), .B2(n_671), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_793), .Y(n_945) );
OAI221xp5_ASAP7_75t_L g946 ( .A1(n_897), .A2(n_720), .B1(n_644), .B2(n_678), .C(n_751), .Y(n_946) );
NOR2xp33_ASAP7_75t_L g947 ( .A(n_785), .B(n_644), .Y(n_947) );
OAI22xp33_ASAP7_75t_SL g948 ( .A1(n_813), .A2(n_678), .B1(n_672), .B2(n_665), .Y(n_948) );
OAI211xp5_ASAP7_75t_L g949 ( .A1(n_822), .A2(n_711), .B(n_703), .C(n_773), .Y(n_949) );
A2O1A1Ixp33_ASAP7_75t_L g950 ( .A1(n_817), .A2(n_880), .B(n_804), .C(n_834), .Y(n_950) );
OR2x2_ASAP7_75t_L g951 ( .A(n_801), .B(n_64), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_792), .B(n_65), .Y(n_952) );
INVx3_ASAP7_75t_L g953 ( .A(n_827), .Y(n_953) );
OAI221xp5_ASAP7_75t_L g954 ( .A1(n_792), .A2(n_711), .B1(n_773), .B2(n_67), .C(n_68), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_831), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_875), .B(n_65), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g957 ( .A1(n_819), .A2(n_66), .B1(n_67), .B2(n_69), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g958 ( .A1(n_819), .A2(n_66), .B1(n_69), .B2(n_70), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_823), .B(n_71), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_876), .Y(n_960) );
AOI21xp5_ASAP7_75t_L g961 ( .A1(n_814), .A2(n_210), .B(n_270), .Y(n_961) );
OAI22xp33_ASAP7_75t_L g962 ( .A1(n_832), .A2(n_72), .B1(n_74), .B2(n_75), .Y(n_962) );
AOI21xp5_ASAP7_75t_L g963 ( .A1(n_782), .A2(n_212), .B(n_267), .Y(n_963) );
INVx2_ASAP7_75t_L g964 ( .A(n_777), .Y(n_964) );
INVx1_ASAP7_75t_SL g965 ( .A(n_787), .Y(n_965) );
NOR2xp33_ASAP7_75t_L g966 ( .A(n_836), .B(n_72), .Y(n_966) );
NOR2xp33_ASAP7_75t_L g967 ( .A(n_845), .B(n_76), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_876), .Y(n_968) );
AOI322xp5_ASAP7_75t_L g969 ( .A1(n_892), .A2(n_76), .A3(n_127), .B1(n_131), .B2(n_133), .C1(n_135), .C2(n_138), .Y(n_969) );
INVx2_ASAP7_75t_L g970 ( .A(n_777), .Y(n_970) );
AOI221xp5_ASAP7_75t_L g971 ( .A1(n_878), .A2(n_852), .B1(n_859), .B2(n_918), .C(n_869), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_898), .B(n_876), .Y(n_972) );
INVx2_ASAP7_75t_SL g973 ( .A(n_790), .Y(n_973) );
AO21x2_ASAP7_75t_L g974 ( .A1(n_820), .A2(n_141), .B(n_145), .Y(n_974) );
INVx3_ASAP7_75t_L g975 ( .A(n_827), .Y(n_975) );
AO21x2_ASAP7_75t_L g976 ( .A1(n_821), .A2(n_147), .B(n_151), .Y(n_976) );
CKINVDCx5p33_ASAP7_75t_R g977 ( .A(n_816), .Y(n_977) );
OAI21x1_ASAP7_75t_L g978 ( .A1(n_815), .A2(n_155), .B(n_158), .Y(n_978) );
NOR2xp33_ASAP7_75t_L g979 ( .A(n_845), .B(n_159), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_868), .A2(n_160), .B1(n_161), .B2(n_162), .Y(n_980) );
INVx2_ASAP7_75t_L g981 ( .A(n_789), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_824), .B(n_166), .Y(n_982) );
OAI211xp5_ASAP7_75t_L g983 ( .A1(n_915), .A2(n_168), .B(n_170), .C(n_172), .Y(n_983) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_868), .A2(n_176), .B1(n_201), .B2(n_205), .Y(n_984) );
NAND4xp25_ASAP7_75t_L g985 ( .A(n_915), .B(n_206), .C(n_207), .D(n_208), .Y(n_985) );
OAI21xp33_ASAP7_75t_L g986 ( .A1(n_810), .A2(n_213), .B(n_214), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_830), .A2(n_217), .B1(n_218), .B2(n_222), .Y(n_987) );
AOI21xp5_ASAP7_75t_L g988 ( .A1(n_776), .A2(n_223), .B(n_224), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_903), .A2(n_226), .B1(n_228), .B2(n_230), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_870), .Y(n_990) );
AND2x4_ASAP7_75t_L g991 ( .A(n_806), .B(n_233), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_886), .A2(n_234), .B1(n_237), .B2(n_239), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_868), .A2(n_241), .B1(n_243), .B2(n_246), .Y(n_993) );
NAND3xp33_ASAP7_75t_L g994 ( .A(n_834), .B(n_842), .C(n_848), .Y(n_994) );
HB1xp67_ASAP7_75t_L g995 ( .A(n_789), .Y(n_995) );
NOR2x1p5_ASAP7_75t_L g996 ( .A(n_790), .B(n_247), .Y(n_996) );
OAI22xp5_ASAP7_75t_L g997 ( .A1(n_870), .A2(n_248), .B1(n_249), .B2(n_251), .Y(n_997) );
BUFx2_ASAP7_75t_L g998 ( .A(n_855), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_807), .B(n_252), .Y(n_999) );
AOI221xp5_ASAP7_75t_L g1000 ( .A1(n_866), .A2(n_253), .B1(n_256), .B2(n_259), .C(n_261), .Y(n_1000) );
OAI221xp5_ASAP7_75t_L g1001 ( .A1(n_921), .A2(n_262), .B1(n_308), .B2(n_798), .C(n_779), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_922), .A2(n_921), .B1(n_907), .B2(n_826), .Y(n_1002) );
OAI22xp33_ASAP7_75t_L g1003 ( .A1(n_854), .A2(n_911), .B1(n_780), .B2(n_916), .Y(n_1003) );
HB1xp67_ASAP7_75t_L g1004 ( .A(n_802), .Y(n_1004) );
AND2x4_ASAP7_75t_L g1005 ( .A(n_806), .B(n_887), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_818), .B(n_917), .Y(n_1006) );
OAI22xp33_ASAP7_75t_L g1007 ( .A1(n_854), .A2(n_911), .B1(n_916), .B2(n_877), .Y(n_1007) );
AND2x2_ASAP7_75t_SL g1008 ( .A(n_887), .B(n_913), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_913), .A2(n_808), .B1(n_889), .B2(n_906), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_906), .A2(n_788), .B1(n_800), .B2(n_919), .Y(n_1010) );
OAI221xp5_ASAP7_75t_SL g1011 ( .A1(n_842), .A2(n_848), .B1(n_849), .B2(n_882), .C(n_825), .Y(n_1011) );
AOI221xp5_ASAP7_75t_L g1012 ( .A1(n_783), .A2(n_882), .B1(n_849), .B2(n_825), .C(n_867), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_802), .B(n_811), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_809), .B(n_811), .Y(n_1014) );
BUFx12f_ASAP7_75t_L g1015 ( .A(n_829), .Y(n_1015) );
OAI22xp5_ASAP7_75t_L g1016 ( .A1(n_809), .A2(n_833), .B1(n_861), .B2(n_871), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_833), .B(n_776), .Y(n_1017) );
NAND2xp5_ASAP7_75t_SL g1018 ( .A(n_912), .B(n_920), .Y(n_1018) );
OAI22xp33_ASAP7_75t_L g1019 ( .A1(n_805), .A2(n_908), .B1(n_857), .B2(n_828), .Y(n_1019) );
OAI22xp33_ASAP7_75t_L g1020 ( .A1(n_805), .A2(n_857), .B1(n_828), .B2(n_776), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_778), .B(n_902), .Y(n_1021) );
OAI211xp5_ASAP7_75t_SL g1022 ( .A1(n_888), .A2(n_799), .B(n_893), .C(n_896), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_778), .B(n_784), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_778), .A2(n_853), .B1(n_795), .B2(n_857), .Y(n_1024) );
AND2x4_ASAP7_75t_L g1025 ( .A(n_912), .B(n_840), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_784), .Y(n_1026) );
OA21x2_ASAP7_75t_L g1027 ( .A1(n_860), .A2(n_899), .B(n_879), .Y(n_1027) );
O2A1O1Ixp33_ASAP7_75t_L g1028 ( .A1(n_841), .A2(n_905), .B(n_839), .C(n_850), .Y(n_1028) );
OAI22xp5_ASAP7_75t_L g1029 ( .A1(n_799), .A2(n_797), .B1(n_847), .B2(n_840), .Y(n_1029) );
OR2x2_ASAP7_75t_L g1030 ( .A(n_797), .B(n_784), .Y(n_1030) );
INVx2_ASAP7_75t_L g1031 ( .A(n_784), .Y(n_1031) );
OA21x2_ASAP7_75t_L g1032 ( .A1(n_860), .A2(n_899), .B(n_843), .Y(n_1032) );
CKINVDCx5p33_ASAP7_75t_R g1033 ( .A(n_912), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_839), .A2(n_850), .B1(n_894), .B2(n_828), .Y(n_1034) );
OAI22xp5_ASAP7_75t_L g1035 ( .A1(n_837), .A2(n_847), .B1(n_873), .B2(n_858), .Y(n_1035) );
INVx2_ASAP7_75t_L g1036 ( .A(n_786), .Y(n_1036) );
OAI21xp5_ASAP7_75t_L g1037 ( .A1(n_796), .A2(n_873), .B(n_891), .Y(n_1037) );
AOI221xp5_ASAP7_75t_L g1038 ( .A1(n_841), .A2(n_905), .B1(n_894), .B2(n_864), .C(n_837), .Y(n_1038) );
NAND3xp33_ASAP7_75t_L g1039 ( .A(n_851), .B(n_909), .C(n_900), .Y(n_1039) );
NAND2xp5_ASAP7_75t_SL g1040 ( .A(n_851), .B(n_909), .Y(n_1040) );
BUFx2_ASAP7_75t_SL g1041 ( .A(n_858), .Y(n_1041) );
AO21x2_ASAP7_75t_L g1042 ( .A1(n_864), .A2(n_914), .B(n_881), .Y(n_1042) );
OR2x2_ASAP7_75t_L g1043 ( .A(n_812), .B(n_900), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_891), .A2(n_835), .B1(n_812), .B2(n_844), .Y(n_1044) );
INVx2_ASAP7_75t_SL g1045 ( .A(n_883), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_885), .B(n_901), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_862), .A2(n_863), .B1(n_865), .B2(n_904), .Y(n_1047) );
BUFx8_ASAP7_75t_SL g1048 ( .A(n_816), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_801), .B(n_537), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_804), .A2(n_651), .B1(n_648), .B2(n_563), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_801), .B(n_537), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_884), .A2(n_890), .B1(n_838), .B2(n_856), .Y(n_1052) );
BUFx3_ASAP7_75t_L g1053 ( .A(n_790), .Y(n_1053) );
BUFx6f_ASAP7_75t_L g1054 ( .A(n_827), .Y(n_1054) );
AOI21xp5_ASAP7_75t_L g1055 ( .A1(n_794), .A2(n_691), .B(n_713), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_1013), .B(n_995), .Y(n_1056) );
AND2x4_ASAP7_75t_L g1057 ( .A(n_990), .B(n_1005), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_995), .B(n_1004), .Y(n_1058) );
HB1xp67_ASAP7_75t_L g1059 ( .A(n_1004), .Y(n_1059) );
INVx3_ASAP7_75t_L g1060 ( .A(n_1054), .Y(n_1060) );
INVx3_ASAP7_75t_L g1061 ( .A(n_1054), .Y(n_1061) );
INVx2_ASAP7_75t_L g1062 ( .A(n_1014), .Y(n_1062) );
INVx2_ASAP7_75t_L g1063 ( .A(n_964), .Y(n_1063) );
OR2x2_ASAP7_75t_L g1064 ( .A(n_1052), .B(n_972), .Y(n_1064) );
AND2x4_ASAP7_75t_L g1065 ( .A(n_1025), .B(n_1037), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_970), .B(n_981), .Y(n_1066) );
INVx2_ASAP7_75t_L g1067 ( .A(n_1017), .Y(n_1067) );
AOI221xp5_ASAP7_75t_L g1068 ( .A1(n_962), .A2(n_971), .B1(n_1050), .B2(n_1011), .C(n_1049), .Y(n_1068) );
BUFx3_ASAP7_75t_L g1069 ( .A(n_1054), .Y(n_1069) );
NAND3xp33_ASAP7_75t_L g1070 ( .A(n_1021), .B(n_969), .C(n_967), .Y(n_1070) );
INVx2_ASAP7_75t_L g1071 ( .A(n_1026), .Y(n_1071) );
OAI21xp5_ASAP7_75t_L g1072 ( .A1(n_950), .A2(n_930), .B(n_1012), .Y(n_1072) );
INVxp67_ASAP7_75t_L g1073 ( .A(n_1051), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1052), .B(n_934), .Y(n_1074) );
INVx2_ASAP7_75t_L g1075 ( .A(n_1031), .Y(n_1075) );
OR2x6_ASAP7_75t_L g1076 ( .A(n_1041), .B(n_991), .Y(n_1076) );
AO21x2_ASAP7_75t_L g1077 ( .A1(n_1020), .A2(n_1019), .B(n_1055), .Y(n_1077) );
OR2x2_ASAP7_75t_L g1078 ( .A(n_935), .B(n_1006), .Y(n_1078) );
BUFx3_ASAP7_75t_L g1079 ( .A(n_1054), .Y(n_1079) );
INVx3_ASAP7_75t_L g1080 ( .A(n_1025), .Y(n_1080) );
AOI22xp5_ASAP7_75t_L g1081 ( .A1(n_962), .A2(n_926), .B1(n_925), .B2(n_1002), .Y(n_1081) );
AO21x2_ASAP7_75t_L g1082 ( .A1(n_1020), .A2(n_1019), .B(n_1028), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_945), .B(n_955), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1023), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g1085 ( .A(n_965), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_960), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_968), .B(n_956), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1030), .Y(n_1088) );
INVx3_ASAP7_75t_L g1089 ( .A(n_991), .Y(n_1089) );
AND2x4_ASAP7_75t_L g1090 ( .A(n_1005), .B(n_996), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1008), .B(n_952), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_927), .B(n_953), .Y(n_1092) );
INVx2_ASAP7_75t_L g1093 ( .A(n_1036), .Y(n_1093) );
INVx2_ASAP7_75t_L g1094 ( .A(n_974), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_933), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1096 ( .A(n_951), .B(n_998), .Y(n_1096) );
OR2x2_ASAP7_75t_L g1097 ( .A(n_959), .B(n_994), .Y(n_1097) );
BUFx6f_ASAP7_75t_SL g1098 ( .A(n_1053), .Y(n_1098) );
INVx3_ASAP7_75t_L g1099 ( .A(n_1033), .Y(n_1099) );
NOR2xp33_ASAP7_75t_L g1100 ( .A(n_977), .B(n_947), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_933), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1008), .B(n_932), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_1007), .A2(n_1009), .B1(n_985), .B2(n_928), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_975), .B(n_966), .Y(n_1104) );
NOR2xp33_ASAP7_75t_L g1105 ( .A(n_973), .B(n_975), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_974), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_976), .Y(n_1107) );
OAI221xp5_ASAP7_75t_SL g1108 ( .A1(n_1003), .A2(n_1007), .B1(n_942), .B2(n_954), .C(n_928), .Y(n_1108) );
INVx2_ASAP7_75t_L g1109 ( .A(n_976), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1039), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1040), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_932), .B(n_999), .Y(n_1112) );
AND2x4_ASAP7_75t_L g1113 ( .A(n_1046), .B(n_1043), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1003), .B(n_931), .Y(n_1114) );
INVx5_ASAP7_75t_L g1115 ( .A(n_1015), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1035), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_993), .B(n_936), .Y(n_1117) );
INVx2_ASAP7_75t_SL g1118 ( .A(n_979), .Y(n_1118) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1045), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1120 ( .A(n_1011), .B(n_943), .Y(n_1120) );
BUFx2_ASAP7_75t_L g1121 ( .A(n_943), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1027), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1027), .Y(n_1123) );
INVx3_ASAP7_75t_L g1124 ( .A(n_978), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_993), .B(n_936), .Y(n_1125) );
BUFx2_ASAP7_75t_L g1126 ( .A(n_1029), .Y(n_1126) );
AND2x4_ASAP7_75t_L g1127 ( .A(n_941), .B(n_1018), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_924), .B(n_957), .Y(n_1128) );
BUFx3_ASAP7_75t_L g1129 ( .A(n_1048), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_958), .B(n_982), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_944), .B(n_989), .Y(n_1131) );
INVx3_ASAP7_75t_L g1132 ( .A(n_1032), .Y(n_1132) );
BUFx3_ASAP7_75t_L g1133 ( .A(n_937), .Y(n_1133) );
INVx2_ASAP7_75t_SL g1134 ( .A(n_997), .Y(n_1134) );
AND2x4_ASAP7_75t_L g1135 ( .A(n_944), .B(n_988), .Y(n_1135) );
OR2x2_ASAP7_75t_L g1136 ( .A(n_1016), .B(n_949), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_1001), .A2(n_948), .B1(n_1010), .B2(n_940), .Y(n_1137) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_987), .B(n_984), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1042), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_989), .B(n_992), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_992), .B(n_987), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1028), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_980), .B(n_1034), .Y(n_1143) );
INVxp67_ASAP7_75t_SL g1144 ( .A(n_939), .Y(n_1144) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_983), .B(n_986), .Y(n_1145) );
AND2x4_ASAP7_75t_L g1146 ( .A(n_1044), .B(n_1047), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1024), .Y(n_1147) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_946), .B(n_1024), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1038), .Y(n_1149) );
INVx2_ASAP7_75t_L g1150 ( .A(n_1022), .Y(n_1150) );
INVxp67_ASAP7_75t_SL g1151 ( .A(n_961), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_938), .B(n_1000), .Y(n_1152) );
INVx3_ASAP7_75t_L g1153 ( .A(n_923), .Y(n_1153) );
BUFx3_ASAP7_75t_L g1154 ( .A(n_929), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_963), .B(n_1022), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1049), .B(n_646), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1084), .B(n_1088), .Y(n_1157) );
INVx1_ASAP7_75t_SL g1158 ( .A(n_1076), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_1074), .B(n_1084), .Y(n_1159) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_1078), .B(n_1074), .Y(n_1160) );
BUFx3_ASAP7_75t_L g1161 ( .A(n_1076), .Y(n_1161) );
HB1xp67_ASAP7_75t_L g1162 ( .A(n_1058), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1088), .B(n_1058), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_1056), .B(n_1064), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1056), .B(n_1113), .Y(n_1165) );
HB1xp67_ASAP7_75t_L g1166 ( .A(n_1059), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1064), .B(n_1112), .Y(n_1167) );
AND2x6_ASAP7_75t_L g1168 ( .A(n_1089), .B(n_1117), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1169 ( .A(n_1067), .B(n_1113), .Y(n_1169) );
NOR2xp33_ASAP7_75t_SL g1170 ( .A(n_1076), .B(n_1108), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1113), .B(n_1067), .Y(n_1171) );
NOR2xp33_ASAP7_75t_L g1172 ( .A(n_1073), .B(n_1156), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1113), .B(n_1066), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1066), .B(n_1120), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1120), .B(n_1062), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1071), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1062), .B(n_1071), .Y(n_1177) );
INVx1_ASAP7_75t_SL g1178 ( .A(n_1076), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1112), .B(n_1086), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1075), .Y(n_1180) );
HB1xp67_ASAP7_75t_L g1181 ( .A(n_1085), .Y(n_1181) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1122), .Y(n_1182) );
NAND2xp5_ASAP7_75t_SL g1183 ( .A(n_1090), .B(n_1118), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1063), .B(n_1086), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1122), .Y(n_1185) );
INVx2_ASAP7_75t_L g1186 ( .A(n_1123), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1150), .B(n_1128), .Y(n_1187) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_1068), .A2(n_1081), .B1(n_1102), .B2(n_1103), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1123), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1150), .B(n_1128), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1102), .B(n_1147), .Y(n_1191) );
AOI21xp33_ASAP7_75t_L g1192 ( .A1(n_1134), .A2(n_1137), .B(n_1070), .Y(n_1192) );
INVx2_ASAP7_75t_L g1193 ( .A(n_1132), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1147), .B(n_1087), .Y(n_1194) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1132), .Y(n_1195) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1132), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1093), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1087), .B(n_1149), .Y(n_1198) );
NAND4xp25_ASAP7_75t_L g1199 ( .A(n_1081), .B(n_1097), .C(n_1152), .D(n_1114), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1078), .B(n_1097), .Y(n_1200) );
AOI221xp5_ASAP7_75t_L g1201 ( .A1(n_1072), .A2(n_1104), .B1(n_1092), .B2(n_1083), .C(n_1149), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1096), .B(n_1057), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1143), .B(n_1116), .Y(n_1203) );
INVx4_ASAP7_75t_L g1204 ( .A(n_1089), .Y(n_1204) );
OR2x2_ASAP7_75t_L g1205 ( .A(n_1096), .B(n_1126), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1116), .B(n_1117), .Y(n_1206) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_1125), .A2(n_1141), .B1(n_1140), .B2(n_1131), .Y(n_1207) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1125), .B(n_1089), .Y(n_1208) );
NAND2xp5_ASAP7_75t_L g1209 ( .A(n_1057), .B(n_1091), .Y(n_1209) );
CKINVDCx5p33_ASAP7_75t_R g1210 ( .A(n_1129), .Y(n_1210) );
INVx3_ASAP7_75t_L g1211 ( .A(n_1146), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1057), .B(n_1091), .Y(n_1212) );
NAND4xp25_ASAP7_75t_L g1213 ( .A(n_1153), .B(n_1133), .C(n_1090), .D(n_1129), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1143), .B(n_1065), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1095), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1095), .Y(n_1216) );
HB1xp67_ASAP7_75t_L g1217 ( .A(n_1090), .Y(n_1217) );
INVx2_ASAP7_75t_L g1218 ( .A(n_1139), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1065), .B(n_1146), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1101), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1101), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1118), .B(n_1130), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1130), .B(n_1144), .Y(n_1223) );
OR2x2_ASAP7_75t_SL g1224 ( .A(n_1136), .B(n_1148), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1065), .B(n_1146), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1139), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1065), .B(n_1146), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1077), .B(n_1082), .Y(n_1228) );
AND2x4_ASAP7_75t_L g1229 ( .A(n_1127), .B(n_1119), .Y(n_1229) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1119), .Y(n_1230) );
OR2x2_ASAP7_75t_L g1231 ( .A(n_1126), .B(n_1121), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1111), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1173), .B(n_1080), .Y(n_1233) );
HB1xp67_ASAP7_75t_L g1234 ( .A(n_1166), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1162), .B(n_1121), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1200), .Y(n_1236) );
NOR2xp33_ASAP7_75t_L g1237 ( .A(n_1199), .B(n_1134), .Y(n_1237) );
OAI21xp5_ASAP7_75t_L g1238 ( .A1(n_1192), .A2(n_1199), .B(n_1188), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1173), .B(n_1165), .Y(n_1239) );
AND2x4_ASAP7_75t_L g1240 ( .A(n_1229), .B(n_1127), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1200), .Y(n_1241) );
INVx2_ASAP7_75t_L g1242 ( .A(n_1182), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1157), .Y(n_1243) );
AND2x4_ASAP7_75t_L g1244 ( .A(n_1229), .B(n_1127), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1157), .Y(n_1245) );
AOI22xp33_ASAP7_75t_L g1246 ( .A1(n_1192), .A2(n_1141), .B1(n_1140), .B2(n_1138), .Y(n_1246) );
NAND2xp5_ASAP7_75t_SL g1247 ( .A(n_1170), .B(n_1127), .Y(n_1247) );
NOR2xp33_ASAP7_75t_L g1248 ( .A(n_1222), .B(n_1099), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1214), .B(n_1077), .Y(n_1249) );
OR2x2_ASAP7_75t_L g1250 ( .A(n_1164), .B(n_1153), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1198), .B(n_1080), .Y(n_1251) );
OR2x2_ASAP7_75t_L g1252 ( .A(n_1164), .B(n_1080), .Y(n_1252) );
NOR2xp33_ASAP7_75t_L g1253 ( .A(n_1223), .B(n_1099), .Y(n_1253) );
INVx3_ASAP7_75t_L g1254 ( .A(n_1204), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1165), .B(n_1079), .Y(n_1255) );
INVx4_ASAP7_75t_L g1256 ( .A(n_1161), .Y(n_1256) );
OR2x2_ASAP7_75t_L g1257 ( .A(n_1169), .B(n_1069), .Y(n_1257) );
HB1xp67_ASAP7_75t_L g1258 ( .A(n_1230), .Y(n_1258) );
NAND2xp5_ASAP7_75t_L g1259 ( .A(n_1194), .B(n_1111), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1163), .B(n_1069), .Y(n_1260) );
OR2x2_ASAP7_75t_L g1261 ( .A(n_1169), .B(n_1079), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1262 ( .A(n_1160), .B(n_1100), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1181), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1194), .B(n_1207), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1163), .B(n_1060), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1184), .Y(n_1266) );
NOR2xp33_ASAP7_75t_R g1267 ( .A(n_1170), .B(n_1115), .Y(n_1267) );
AND2x4_ASAP7_75t_SL g1268 ( .A(n_1217), .B(n_1099), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1184), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1171), .B(n_1060), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1201), .B(n_1110), .Y(n_1271) );
NOR2x1_ASAP7_75t_L g1272 ( .A(n_1213), .B(n_1161), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1171), .B(n_1060), .Y(n_1273) );
NAND3xp33_ASAP7_75t_L g1274 ( .A(n_1172), .B(n_1105), .C(n_1142), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1185), .Y(n_1275) );
CKINVDCx16_ASAP7_75t_R g1276 ( .A(n_1224), .Y(n_1276) );
OR2x2_ASAP7_75t_L g1277 ( .A(n_1205), .B(n_1061), .Y(n_1277) );
INVx1_ASAP7_75t_SL g1278 ( .A(n_1210), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1174), .B(n_1110), .Y(n_1279) );
NAND4xp25_ASAP7_75t_SL g1280 ( .A(n_1158), .B(n_1115), .C(n_1098), .D(n_1136), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1185), .Y(n_1281) );
NAND3xp33_ASAP7_75t_SL g1282 ( .A(n_1158), .B(n_1115), .C(n_1098), .Y(n_1282) );
HB1xp67_ASAP7_75t_L g1283 ( .A(n_1230), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1189), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1214), .B(n_1155), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1189), .Y(n_1286) );
OR2x2_ASAP7_75t_L g1287 ( .A(n_1159), .B(n_1077), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1175), .B(n_1155), .Y(n_1288) );
INVx2_ASAP7_75t_SL g1289 ( .A(n_1161), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1202), .B(n_1135), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1175), .B(n_1142), .Y(n_1291) );
HB1xp67_ASAP7_75t_L g1292 ( .A(n_1230), .Y(n_1292) );
INVx3_ASAP7_75t_L g1293 ( .A(n_1254), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1285), .B(n_1227), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1234), .Y(n_1295) );
INVx1_ASAP7_75t_SL g1296 ( .A(n_1278), .Y(n_1296) );
OR2x2_ASAP7_75t_L g1297 ( .A(n_1236), .B(n_1231), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1249), .B(n_1227), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1241), .B(n_1203), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_1264), .B(n_1203), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1249), .B(n_1290), .Y(n_1301) );
OR2x2_ASAP7_75t_L g1302 ( .A(n_1287), .B(n_1231), .Y(n_1302) );
NOR3xp33_ASAP7_75t_L g1303 ( .A(n_1238), .B(n_1183), .C(n_1187), .Y(n_1303) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1234), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1243), .B(n_1191), .Y(n_1305) );
OR2x6_ASAP7_75t_L g1306 ( .A(n_1272), .B(n_1254), .Y(n_1306) );
CKINVDCx16_ASAP7_75t_R g1307 ( .A(n_1276), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1263), .Y(n_1308) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1275), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1239), .B(n_1219), .Y(n_1310) );
OAI22xp5_ASAP7_75t_L g1311 ( .A1(n_1246), .A2(n_1224), .B1(n_1178), .B2(n_1212), .Y(n_1311) );
INVxp67_ASAP7_75t_SL g1312 ( .A(n_1258), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1288), .B(n_1219), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1281), .Y(n_1314) );
NAND2xp33_ASAP7_75t_L g1315 ( .A(n_1267), .B(n_1168), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1284), .Y(n_1316) );
INVx2_ASAP7_75t_L g1317 ( .A(n_1242), .Y(n_1317) );
OR2x2_ASAP7_75t_L g1318 ( .A(n_1235), .B(n_1291), .Y(n_1318) );
INVx1_ASAP7_75t_SL g1319 ( .A(n_1260), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1240), .B(n_1225), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1240), .B(n_1225), .Y(n_1321) );
BUFx2_ASAP7_75t_L g1322 ( .A(n_1254), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1245), .B(n_1191), .Y(n_1323) );
AOI21xp5_ASAP7_75t_L g1324 ( .A1(n_1282), .A2(n_1145), .B(n_1178), .Y(n_1324) );
INVxp67_ASAP7_75t_L g1325 ( .A(n_1250), .Y(n_1325) );
NAND2xp67_ASAP7_75t_L g1326 ( .A(n_1268), .B(n_1228), .Y(n_1326) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1286), .Y(n_1327) );
OR2x2_ASAP7_75t_L g1328 ( .A(n_1259), .B(n_1206), .Y(n_1328) );
OR2x2_ASAP7_75t_L g1329 ( .A(n_1279), .B(n_1206), .Y(n_1329) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_1266), .B(n_1208), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1240), .B(n_1211), .Y(n_1331) );
INVx1_ASAP7_75t_SL g1332 ( .A(n_1255), .Y(n_1332) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1269), .Y(n_1333) );
INVx2_ASAP7_75t_L g1334 ( .A(n_1242), .Y(n_1334) );
INVx2_ASAP7_75t_L g1335 ( .A(n_1258), .Y(n_1335) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1252), .Y(n_1336) );
INVx1_ASAP7_75t_SL g1337 ( .A(n_1319), .Y(n_1337) );
AOI22xp5_ASAP7_75t_L g1338 ( .A1(n_1311), .A2(n_1237), .B1(n_1246), .B2(n_1247), .Y(n_1338) );
AOI221x1_ASAP7_75t_L g1339 ( .A1(n_1303), .A2(n_1274), .B1(n_1271), .B2(n_1237), .C(n_1253), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1301), .B(n_1233), .Y(n_1340) );
INVx2_ASAP7_75t_L g1341 ( .A(n_1335), .Y(n_1341) );
NAND2x1_ASAP7_75t_L g1342 ( .A(n_1306), .B(n_1168), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1300), .B(n_1187), .Y(n_1343) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1295), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1304), .B(n_1190), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1313), .B(n_1190), .Y(n_1346) );
AOI21xp5_ASAP7_75t_L g1347 ( .A1(n_1315), .A2(n_1280), .B(n_1283), .Y(n_1347) );
NAND4xp25_ASAP7_75t_L g1348 ( .A(n_1324), .B(n_1253), .C(n_1248), .D(n_1251), .Y(n_1348) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1308), .Y(n_1349) );
AOI21xp33_ASAP7_75t_SL g1350 ( .A1(n_1307), .A2(n_1248), .B(n_1289), .Y(n_1350) );
INVxp67_ASAP7_75t_L g1351 ( .A(n_1322), .Y(n_1351) );
O2A1O1Ixp33_ASAP7_75t_L g1352 ( .A1(n_1315), .A2(n_1262), .B(n_1154), .C(n_1208), .Y(n_1352) );
NAND2xp5_ASAP7_75t_L g1353 ( .A(n_1313), .B(n_1167), .Y(n_1353) );
AOI22xp5_ASAP7_75t_L g1354 ( .A1(n_1325), .A2(n_1168), .B1(n_1265), .B2(n_1244), .Y(n_1354) );
OAI21xp33_ASAP7_75t_L g1355 ( .A1(n_1326), .A2(n_1301), .B(n_1298), .Y(n_1355) );
OAI22xp5_ASAP7_75t_L g1356 ( .A1(n_1306), .A2(n_1268), .B1(n_1256), .B2(n_1261), .Y(n_1356) );
INVx1_ASAP7_75t_SL g1357 ( .A(n_1332), .Y(n_1357) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1309), .Y(n_1358) );
OAI21xp5_ASAP7_75t_SL g1359 ( .A1(n_1322), .A2(n_1228), .B(n_1244), .Y(n_1359) );
AOI221xp5_ASAP7_75t_L g1360 ( .A1(n_1336), .A2(n_1167), .B1(n_1179), .B2(n_1267), .C(n_1209), .Y(n_1360) );
AOI22xp5_ASAP7_75t_L g1361 ( .A1(n_1333), .A2(n_1168), .B1(n_1244), .B2(n_1270), .Y(n_1361) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_1331), .A2(n_1168), .B1(n_1211), .B2(n_1229), .Y(n_1362) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1314), .Y(n_1363) );
AOI32xp33_ASAP7_75t_L g1364 ( .A1(n_1296), .A2(n_1256), .A3(n_1273), .B1(n_1204), .B2(n_1289), .Y(n_1364) );
AOI22xp33_ASAP7_75t_L g1365 ( .A1(n_1331), .A2(n_1168), .B1(n_1211), .B2(n_1229), .Y(n_1365) );
NAND2xp5_ASAP7_75t_L g1366 ( .A(n_1343), .B(n_1298), .Y(n_1366) );
NAND2xp5_ASAP7_75t_SL g1367 ( .A(n_1364), .B(n_1293), .Y(n_1367) );
OAI22xp33_ASAP7_75t_L g1368 ( .A1(n_1338), .A2(n_1306), .B1(n_1293), .B2(n_1256), .Y(n_1368) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1358), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1363), .Y(n_1370) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1349), .Y(n_1371) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1344), .Y(n_1372) );
OAI22xp5_ASAP7_75t_L g1373 ( .A1(n_1350), .A2(n_1293), .B1(n_1329), .B2(n_1318), .Y(n_1373) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1345), .Y(n_1374) );
OAI222xp33_ASAP7_75t_L g1375 ( .A1(n_1337), .A2(n_1318), .B1(n_1329), .B2(n_1302), .C1(n_1328), .C2(n_1297), .Y(n_1375) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1346), .Y(n_1376) );
OAI22xp5_ASAP7_75t_L g1377 ( .A1(n_1355), .A2(n_1328), .B1(n_1297), .B2(n_1302), .Y(n_1377) );
AOI221xp5_ASAP7_75t_L g1378 ( .A1(n_1348), .A2(n_1299), .B1(n_1294), .B2(n_1323), .C(n_1305), .Y(n_1378) );
OAI22xp33_ASAP7_75t_L g1379 ( .A1(n_1342), .A2(n_1204), .B1(n_1330), .B2(n_1257), .Y(n_1379) );
OAI31xp33_ASAP7_75t_L g1380 ( .A1(n_1357), .A2(n_1320), .A3(n_1321), .B(n_1294), .Y(n_1380) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1341), .Y(n_1381) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1353), .Y(n_1382) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1340), .Y(n_1383) );
NOR2xp33_ASAP7_75t_L g1384 ( .A(n_1351), .B(n_1310), .Y(n_1384) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1352), .Y(n_1385) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1369), .Y(n_1386) );
AOI221x1_ASAP7_75t_L g1387 ( .A1(n_1385), .A2(n_1347), .B1(n_1356), .B2(n_1327), .C(n_1316), .Y(n_1387) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1370), .Y(n_1388) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1371), .Y(n_1389) );
AOI211xp5_ASAP7_75t_L g1390 ( .A1(n_1368), .A2(n_1373), .B(n_1367), .C(n_1375), .Y(n_1390) );
OA22x2_ASAP7_75t_L g1391 ( .A1(n_1377), .A2(n_1359), .B1(n_1339), .B2(n_1354), .Y(n_1391) );
NOR2xp67_ASAP7_75t_L g1392 ( .A(n_1384), .B(n_1347), .Y(n_1392) );
OAI32xp33_ASAP7_75t_L g1393 ( .A1(n_1384), .A2(n_1330), .A3(n_1352), .B1(n_1326), .B2(n_1365), .Y(n_1393) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1372), .Y(n_1394) );
NOR4xp25_ASAP7_75t_L g1395 ( .A(n_1368), .B(n_1360), .C(n_1310), .D(n_1232), .Y(n_1395) );
AOI221xp5_ASAP7_75t_L g1396 ( .A1(n_1378), .A2(n_1320), .B1(n_1321), .B2(n_1312), .C(n_1362), .Y(n_1396) );
AOI22xp5_ASAP7_75t_L g1397 ( .A1(n_1379), .A2(n_1168), .B1(n_1361), .B2(n_1115), .Y(n_1397) );
AOI221xp5_ASAP7_75t_L g1398 ( .A1(n_1376), .A2(n_1179), .B1(n_1211), .B2(n_1335), .C(n_1098), .Y(n_1398) );
AOI211xp5_ASAP7_75t_L g1399 ( .A1(n_1393), .A2(n_1379), .B(n_1380), .C(n_1382), .Y(n_1399) );
AOI322xp5_ASAP7_75t_L g1400 ( .A1(n_1396), .A2(n_1383), .A3(n_1366), .B1(n_1374), .B2(n_1381), .C1(n_1115), .C2(n_1283), .Y(n_1400) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1386), .Y(n_1401) );
AOI22xp5_ASAP7_75t_L g1402 ( .A1(n_1391), .A2(n_1115), .B1(n_1082), .B2(n_1277), .Y(n_1402) );
NAND2xp5_ASAP7_75t_SL g1403 ( .A(n_1395), .B(n_1334), .Y(n_1403) );
NAND3xp33_ASAP7_75t_L g1404 ( .A(n_1390), .B(n_1226), .C(n_1232), .Y(n_1404) );
AOI221xp5_ASAP7_75t_L g1405 ( .A1(n_1388), .A2(n_1334), .B1(n_1317), .B2(n_1221), .C(n_1220), .Y(n_1405) );
OAI21xp33_ASAP7_75t_L g1406 ( .A1(n_1392), .A2(n_1317), .B(n_1215), .Y(n_1406) );
NOR2x1_ASAP7_75t_L g1407 ( .A(n_1404), .B(n_1394), .Y(n_1407) );
OAI211xp5_ASAP7_75t_L g1408 ( .A1(n_1402), .A2(n_1387), .B(n_1397), .C(n_1398), .Y(n_1408) );
CKINVDCx5p33_ASAP7_75t_R g1409 ( .A(n_1401), .Y(n_1409) );
NOR4xp25_ASAP7_75t_SL g1410 ( .A(n_1406), .B(n_1389), .C(n_1397), .D(n_1151), .Y(n_1410) );
NAND2x1p5_ASAP7_75t_L g1411 ( .A(n_1403), .B(n_1204), .Y(n_1411) );
NAND5xp2_ASAP7_75t_L g1412 ( .A(n_1399), .B(n_1107), .C(n_1106), .D(n_1220), .E(n_1216), .Y(n_1412) );
AOI22xp5_ASAP7_75t_L g1413 ( .A1(n_1409), .A2(n_1405), .B1(n_1400), .B2(n_1082), .Y(n_1413) );
AOI222xp33_ASAP7_75t_L g1414 ( .A1(n_1408), .A2(n_1221), .B1(n_1215), .B2(n_1216), .C1(n_1292), .C2(n_1218), .Y(n_1414) );
OR4x2_ASAP7_75t_L g1415 ( .A(n_1412), .B(n_1135), .C(n_1177), .D(n_1218), .Y(n_1415) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1407), .Y(n_1416) );
AOI221x1_ASAP7_75t_L g1417 ( .A1(n_1416), .A2(n_1414), .B1(n_1410), .B2(n_1415), .C(n_1413), .Y(n_1417) );
AO21x2_ASAP7_75t_L g1418 ( .A1(n_1416), .A2(n_1411), .B(n_1094), .Y(n_1418) );
XNOR2xp5_ASAP7_75t_L g1419 ( .A(n_1417), .B(n_1135), .Y(n_1419) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_1419), .B(n_1418), .Y(n_1420) );
AOI22xp33_ASAP7_75t_L g1421 ( .A1(n_1420), .A2(n_1418), .B1(n_1196), .B2(n_1195), .Y(n_1421) );
AOI322xp5_ASAP7_75t_L g1422 ( .A1(n_1421), .A2(n_1109), .A3(n_1124), .B1(n_1196), .B2(n_1195), .C1(n_1193), .C2(n_1180), .Y(n_1422) );
AOI221xp5_ASAP7_75t_L g1423 ( .A1(n_1422), .A2(n_1193), .B1(n_1176), .B2(n_1197), .C(n_1186), .Y(n_1423) );
endmodule