module real_jpeg_13069_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_3),
.A2(n_37),
.B(n_38),
.C(n_44),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_3),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_3),
.B(n_128),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_3),
.B(n_41),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_SL g177 ( 
.A1(n_3),
.A2(n_41),
.B(n_163),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_3),
.B(n_25),
.C(n_87),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_3),
.A2(n_40),
.B1(n_53),
.B2(n_57),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_3),
.A2(n_24),
.B1(n_28),
.B2(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_3),
.B(n_63),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_71),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_5),
.A2(n_53),
.B1(n_57),
.B2(n_71),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_5),
.A2(n_25),
.B1(n_32),
.B2(n_71),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_6),
.A2(n_25),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_6),
.A2(n_31),
.B1(n_53),
.B2(n_57),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_7),
.A2(n_25),
.B1(n_32),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_7),
.A2(n_34),
.B1(n_53),
.B2(n_57),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_9),
.A2(n_25),
.B1(n_32),
.B2(n_62),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_9),
.A2(n_53),
.B1(n_57),
.B2(n_62),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_12),
.A2(n_25),
.B1(n_32),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_12),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_12),
.A2(n_53),
.B1(n_57),
.B2(n_81),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_81),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_69),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_13),
.A2(n_53),
.B1(n_57),
.B2(n_69),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_13),
.A2(n_25),
.B1(n_32),
.B2(n_69),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_50),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_14),
.A2(n_50),
.B1(n_53),
.B2(n_57),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_14),
.A2(n_25),
.B1(n_32),
.B2(n_50),
.Y(n_194)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_132),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_111),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_19),
.B(n_111),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_72),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_48),
.C(n_64),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_21),
.B(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_35),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_22),
.A2(n_35),
.B1(n_36),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_22),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_23),
.A2(n_78),
.B(n_99),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_23),
.A2(n_29),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_24),
.B(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_24),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_24),
.A2(n_28),
.B1(n_192),
.B2(n_200),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_24),
.A2(n_77),
.B(n_194),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_25),
.A2(n_32),
.B1(n_87),
.B2(n_88),
.Y(n_90)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_28),
.B(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_28),
.B(n_40),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_29),
.B(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_29),
.A2(n_30),
.B(n_79),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_32),
.B(n_198),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_33),
.Y(n_97)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_37),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_37),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_37),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B(n_41),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_40),
.B(n_90),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_42),
.B1(n_55),
.B2(n_56),
.Y(n_58)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND3xp33_ASAP7_75t_SL g164 ( 
.A(n_42),
.B(n_55),
.C(n_57),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_48),
.B(n_64),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_51),
.B(n_59),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_49),
.A2(n_51),
.B1(n_52),
.B2(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_51),
.A2(n_61),
.B(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_51),
.A2(n_52),
.B1(n_123),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_51),
.A2(n_52),
.B1(n_147),
.B2(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_58),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_52)
);

INVx5_ASAP7_75t_SL g57 ( 
.A(n_53),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_57),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_53),
.A2(n_56),
.B(n_162),
.C(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_53),
.B(n_186),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_63),
.B(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_70),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_65),
.A2(n_66),
.B1(n_70),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_68),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_94),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_82),
.B2(n_93),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B1(n_91),
.B2(n_92),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_90),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_85),
.A2(n_91),
.B1(n_157),
.B2(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_85),
.A2(n_91),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_85),
.A2(n_91),
.B1(n_179),
.B2(n_189),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_91),
.B(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_91),
.B(n_119),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_103),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_100),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_107),
.B2(n_110),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.C(n_129),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_112),
.B(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_114),
.B(n_129),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_121),
.C(n_124),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_116),
.B1(n_121),
.B2(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B(n_120),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_117),
.A2(n_156),
.B(n_158),
.Y(n_155)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_124),
.B(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_228),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_223),
.B(n_224),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_167),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_152),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_137),
.B(n_152),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_150),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_141),
.B1(n_148),
.B2(n_149),
.Y(n_138)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_141),
.B(n_148),
.C(n_150),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.C(n_146),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_154)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_146),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.C(n_159),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_155),
.A2(n_159),
.B1(n_160),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_165),
.B1(n_166),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_180),
.B(n_222),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_169),
.B(n_172),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.C(n_178),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_216),
.B(n_221),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_206),
.B(n_215),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_195),
.B(n_205),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_190),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_190),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_187),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_201),
.B(n_204),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_208),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_211),
.C(n_214),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_213),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_220),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_227),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);


endmodule