module fake_netlist_1_12376_n_31 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_31);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx8_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
NAND2xp5_ASAP7_75t_SL g14 ( .A(n_8), .B(n_11), .Y(n_14) );
BUFx2_ASAP7_75t_L g15 ( .A(n_3), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_5), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_5), .Y(n_18) );
NOR3xp33_ASAP7_75t_SL g19 ( .A(n_18), .B(n_1), .C(n_2), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
A2O1A1Ixp33_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_15), .B(n_17), .C(n_18), .Y(n_21) );
AOI22xp33_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_15), .B1(n_13), .B2(n_14), .Y(n_22) );
OAI33xp33_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_19), .A3(n_13), .B1(n_3), .B2(n_4), .B3(n_6), .Y(n_23) );
OR2x2_ASAP7_75t_L g24 ( .A(n_23), .B(n_22), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_24), .B(n_1), .Y(n_25) );
OAI21x1_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_9), .B(n_12), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_13), .B1(n_4), .B2(n_6), .Y(n_27) );
BUFx12f_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
CKINVDCx5p33_ASAP7_75t_R g29 ( .A(n_26), .Y(n_29) );
OAI22x1_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_2), .B1(n_7), .B2(n_10), .Y(n_30) );
AOI222xp33_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_7), .B1(n_28), .B2(n_23), .C1(n_29), .C2(n_13), .Y(n_31) );
endmodule