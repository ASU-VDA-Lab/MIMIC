module fake_netlist_6_2577_n_4421 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_466, n_506, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_493, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_514, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4421);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_493;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_514;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4421;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3813;
wire n_3660;
wire n_801;
wire n_3766;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3783;
wire n_700;
wire n_3773;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_3844;
wire n_4388;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_4395;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4168;
wire n_783;
wire n_4372;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_4370;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_4050;
wire n_3706;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_873;
wire n_1371;
wire n_1285;
wire n_2974;
wire n_2886;
wire n_3946;
wire n_4213;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_852;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_836;
wire n_3345;
wire n_2074;
wire n_4417;
wire n_2447;
wire n_522;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_4308;
wire n_616;
wire n_658;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_4325;
wire n_2212;
wire n_3929;
wire n_758;
wire n_516;
wire n_3494;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_4187;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_538;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3737;
wire n_3624;
wire n_3077;
wire n_3979;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_539;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_1404;
wire n_638;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_4414;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_4262;
wire n_4392;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_1815;
wire n_659;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_913;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4071;
wire n_4255;
wire n_4403;
wire n_3506;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_551;
wire n_1986;
wire n_699;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_564;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4349;
wire n_824;
wire n_686;
wire n_4102;
wire n_4297;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_577;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_619;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_572;
wire n_4314;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_606;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_3910;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4415;
wire n_4296;
wire n_4009;
wire n_2633;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_630;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_541;
wire n_2669;
wire n_2925;
wire n_4094;
wire n_3728;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_792;
wire n_2522;
wire n_3949;
wire n_4364;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_4393;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_982;
wire n_4257;
wire n_2674;
wire n_2832;
wire n_4226;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_932;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_4366;
wire n_3446;
wire n_4158;
wire n_4377;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_905;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_993;
wire n_2692;
wire n_3842;
wire n_689;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_966;
wire n_3888;
wire n_2908;
wire n_3168;
wire n_764;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4161;
wire n_4130;
wire n_4337;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3055;
wire n_3092;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_4369;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_1014;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_882;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_586;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_4375;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1912;
wire n_1563;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_702;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_4386;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_690;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_3917;
wire n_1654;
wire n_816;
wire n_4371;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_4043;
wire n_825;
wire n_4313;
wire n_728;
wire n_4353;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_4381;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_4418;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_696;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_593;
wire n_4169;
wire n_4055;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_3271;
wire n_950;
wire n_4362;
wire n_4248;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_4361;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_4367;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_590;
wire n_4394;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_3073;
wire n_2431;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_595;
wire n_1767;
wire n_627;
wire n_3253;
wire n_1779;
wire n_524;
wire n_1465;
wire n_3337;
wire n_3450;
wire n_3431;
wire n_3209;
wire n_4002;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_4288;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4289;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_815;
wire n_3953;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_4385;
wire n_1952;
wire n_865;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_4191;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_963;
wire n_639;
wire n_2767;
wire n_794;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1139;
wire n_1714;
wire n_872;
wire n_3922;
wire n_3179;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_2537;
wire n_2897;
wire n_3970;
wire n_4389;
wire n_4345;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_3171;
wire n_1913;
wire n_791;
wire n_4216;
wire n_3608;
wire n_837;
wire n_4315;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3426;
wire n_1788;
wire n_3158;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2643;
wire n_2590;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_765;
wire n_987;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_705;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_3887;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_4096;
wire n_1431;
wire n_4123;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_4286;
wire n_1809;
wire n_3119;
wire n_4280;
wire n_2958;
wire n_1577;
wire n_2948;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_4379;
wire n_3731;
wire n_1822;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_4218;
wire n_4402;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4264;
wire n_2857;
wire n_3693;
wire n_3788;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2896;
wire n_526;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_4079;
wire n_2494;
wire n_2959;
wire n_3674;
wire n_2501;
wire n_3325;
wire n_3203;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_4175;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_1507;
wire n_2482;
wire n_552;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_745;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_1774;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1398;
wire n_1201;
wire n_884;
wire n_716;
wire n_2354;
wire n_2682;
wire n_3103;
wire n_3032;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_3393;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_2442;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3480;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_958;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_4401;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_4368;
wire n_1478;
wire n_589;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_3591;
wire n_767;
wire n_3641;
wire n_1314;
wire n_600;
wire n_964;
wire n_1837;
wire n_2218;
wire n_831;
wire n_2788;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1564;
wire n_1736;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_3944;
wire n_3909;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_4387;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_3481;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_2990;
wire n_3847;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3323;
wire n_3364;
wire n_3226;
wire n_4020;
wire n_4176;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_4404;
wire n_651;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_4261;
wire n_1745;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_3742;
wire n_4410;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_3243;
wire n_4034;
wire n_4056;
wire n_3683;
wire n_1617;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_4206;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_4132;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_858;
wire n_4149;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_4355;
wire n_2276;
wire n_960;
wire n_956;
wire n_3234;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_3016;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_1129;
wire n_3870;
wire n_4030;
wire n_4126;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_1869;
wire n_664;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_587;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_828;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_4357;
wire n_607;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_4374;
wire n_2201;
wire n_725;
wire n_952;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3276;
wire n_1934;
wire n_3250;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_617;
wire n_3886;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_4420;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3926;
wire n_3797;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_4405;
wire n_610;
wire n_4234;
wire n_4304;
wire n_4413;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_1847;
wire n_2052;
wire n_3634;
wire n_2302;
wire n_517;
wire n_4211;
wire n_4182;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_1037;
wire n_1397;
wire n_621;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_923;
wire n_1409;
wire n_4230;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_4274;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4270;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_710;
wire n_1108;
wire n_1818;
wire n_3730;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_4397;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_4155;
wire n_2740;
wire n_746;
wire n_4238;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_4406;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_4380;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_4398;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4109;
wire n_4192;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4159;
wire n_4195;
wire n_3784;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_1870;
wire n_2964;
wire n_4174;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3475;
wire n_662;
wire n_3501;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_711;
wire n_579;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_4258;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_1823;
wire n_776;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_4135;
wire n_2871;
wire n_4209;
wire n_4279;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_3858;
wire n_4183;
wire n_1489;
wire n_4321;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_543;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_4040;
wire n_804;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_1548;
wire n_799;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_4343;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_652;
wire n_2154;
wire n_2727;
wire n_3377;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_4378;
wire n_4407;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3932;
wire n_3469;
wire n_3958;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_4358;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_655;
wire n_1045;
wire n_1650;
wire n_1794;
wire n_1962;
wire n_706;
wire n_1236;
wire n_786;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_4317;
wire n_834;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_743;
wire n_766;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2671;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_2888;
wire n_3711;
wire n_3776;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_817;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_841;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_4376;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3458;
wire n_3216;
wire n_3515;
wire n_1150;
wire n_4203;
wire n_3808;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_4365;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_591;
wire n_3758;
wire n_1879;
wire n_853;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_680;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2163;
wire n_2186;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_4408;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_4295;
wire n_1120;
wire n_832;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_691;
wire n_535;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_918;
wire n_748;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_957;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_4352;
wire n_744;
wire n_971;
wire n_4391;
wire n_4416;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_1303;
wire n_761;
wire n_2769;
wire n_4342;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_611;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_4106;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4027;
wire n_4373;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_647;
wire n_4160;
wire n_4231;
wire n_844;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2255;
wire n_2112;
wire n_1737;
wire n_1464;
wire n_653;
wire n_2430;
wire n_1414;
wire n_3486;
wire n_4086;
wire n_908;
wire n_752;
wire n_2649;
wire n_2721;
wire n_944;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_1028;
wire n_576;
wire n_3836;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_4409;
wire n_2744;
wire n_4309;
wire n_4363;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_2444;
wire n_839;
wire n_2743;
wire n_3962;
wire n_1973;
wire n_708;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_4166;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1821;
wire n_1537;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3256;
wire n_3868;
wire n_1276;
wire n_3802;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4142;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_1584;
wire n_771;
wire n_2425;
wire n_924;
wire n_3461;
wire n_3408;
wire n_1582;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_719;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_4383;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_2666;
wire n_4105;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_4244;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_1362;
wire n_1156;
wire n_829;
wire n_4259;
wire n_3123;
wire n_2600;
wire n_984;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_570;
wire n_859;
wire n_2033;
wire n_3086;
wire n_4104;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_3285;
wire n_519;
wire n_4208;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_4346;
wire n_4351;
wire n_1144;
wire n_2071;
wire n_3863;
wire n_3669;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_4316;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4390;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_4396;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_3989;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_1606;
wire n_4332;
wire n_810;
wire n_4108;
wire n_1133;
wire n_635;
wire n_1194;
wire n_3374;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_4051;
wire n_1051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_4293;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_3709;
wire n_753;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_3187;
wire n_2540;
wire n_4412;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_4148;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_679;
wire n_4057;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_633;
wire n_1170;
wire n_1629;
wire n_665;
wire n_2221;
wire n_588;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_3903;
wire n_730;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3333;
wire n_3274;
wire n_3186;
wire n_1322;
wire n_640;
wire n_4129;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_3079;
wire n_4360;
wire n_2098;
wire n_3085;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_4039;
wire n_3584;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_4275;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_900;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_827;
wire n_531;
wire n_2912;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g516 ( 
.A(n_464),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_16),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_293),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_174),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_110),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_449),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_508),
.Y(n_522)
);

BUFx10_ASAP7_75t_L g523 ( 
.A(n_282),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_79),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_11),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_492),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_54),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_218),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_142),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_305),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_314),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_337),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_16),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_388),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_99),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_323),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_177),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_46),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_453),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_291),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_420),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_216),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_29),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_338),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_511),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_472),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_364),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_180),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_117),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_128),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_226),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_347),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_96),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_412),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_121),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_368),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_198),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_274),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_141),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_182),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_151),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_319),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_282),
.Y(n_563)
);

CKINVDCx14_ASAP7_75t_R g564 ( 
.A(n_283),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_233),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_503),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_24),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_358),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_476),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_184),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_447),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_324),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_129),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_77),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_159),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_260),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_482),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_135),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_137),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_491),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_167),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_178),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_378),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_263),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_449),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_324),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_467),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_151),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_67),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_337),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_318),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_454),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_448),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_183),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_237),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_310),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_312),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_386),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_104),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_351),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_253),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_411),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_448),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_88),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_312),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_425),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_222),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_167),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_309),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_201),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_303),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_73),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_462),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_176),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_13),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_290),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_451),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_269),
.Y(n_618)
);

BUFx5_ASAP7_75t_L g619 ( 
.A(n_49),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_410),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_367),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_323),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_138),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_490),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_299),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_375),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_33),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_72),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_294),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_58),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_119),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_497),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_43),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_501),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_58),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_35),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_209),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_85),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_357),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_259),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_438),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_386),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_339),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_468),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_257),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_120),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_426),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_433),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_173),
.Y(n_649)
);

BUFx2_ASAP7_75t_SL g650 ( 
.A(n_426),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_236),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_189),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_162),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_232),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_240),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_42),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_455),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_439),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_128),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_418),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_436),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_66),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_289),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_245),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_376),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_400),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_88),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_493),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_378),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_315),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_181),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_32),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_147),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_420),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_247),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_86),
.Y(n_676)
);

BUFx5_ASAP7_75t_L g677 ( 
.A(n_415),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_321),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_106),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_146),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_204),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_366),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_90),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_171),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_163),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_260),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_286),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_404),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_374),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_407),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_44),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_259),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_221),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_233),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_113),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_164),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_325),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_333),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_327),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_155),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_89),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_303),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_89),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_365),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_429),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_349),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_331),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_112),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_358),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_190),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_170),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_494),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_243),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_445),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_9),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_249),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_335),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_56),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_44),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_291),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_141),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_83),
.Y(n_722)
);

INVx1_ASAP7_75t_SL g723 ( 
.A(n_91),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_456),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_137),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_188),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_339),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_427),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_311),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_295),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_111),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_269),
.Y(n_732)
);

CKINVDCx16_ASAP7_75t_R g733 ( 
.A(n_162),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_111),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_316),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_286),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_413),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_77),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_24),
.Y(n_739)
);

BUFx10_ASAP7_75t_L g740 ( 
.A(n_108),
.Y(n_740)
);

BUFx5_ASAP7_75t_L g741 ( 
.A(n_145),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_380),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_417),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_389),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_444),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_314),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_11),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_40),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_352),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_310),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_478),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_346),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_143),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_75),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_447),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_227),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_144),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_355),
.Y(n_758)
);

BUFx10_ASAP7_75t_L g759 ( 
.A(n_254),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_41),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_248),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_331),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_185),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_183),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_396),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_485),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_180),
.Y(n_767)
);

BUFx10_ASAP7_75t_L g768 ( 
.A(n_370),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_135),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_22),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_365),
.Y(n_771)
);

BUFx10_ASAP7_75t_L g772 ( 
.A(n_347),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_357),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_7),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_374),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_199),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_387),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_408),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_220),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_423),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_504),
.Y(n_781)
);

CKINVDCx16_ASAP7_75t_R g782 ( 
.A(n_458),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_481),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_82),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_441),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_178),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_255),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_42),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_372),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_280),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_270),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_345),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_60),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_117),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_179),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_325),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_93),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_515),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_428),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_267),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_62),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_170),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_138),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_175),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_338),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_277),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_26),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_299),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_271),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_361),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_196),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_107),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_496),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_502),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_248),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_446),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_0),
.Y(n_817)
);

CKINVDCx16_ASAP7_75t_R g818 ( 
.A(n_87),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_175),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_333),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_50),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_402),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_15),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_221),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_205),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_394),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_507),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_21),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_290),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_360),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_119),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_432),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_436),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_332),
.Y(n_834)
);

CKINVDCx14_ASAP7_75t_R g835 ( 
.A(n_413),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_526),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_619),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_619),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_619),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_573),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_619),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_619),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_619),
.Y(n_843)
);

NOR2xp67_ASAP7_75t_L g844 ( 
.A(n_622),
.B(n_0),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_619),
.Y(n_845)
);

INVxp67_ASAP7_75t_SL g846 ( 
.A(n_622),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_619),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_619),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_545),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_801),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_677),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_546),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_677),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_677),
.Y(n_854)
);

INVxp33_ASAP7_75t_SL g855 ( 
.A(n_614),
.Y(n_855)
);

INVxp33_ASAP7_75t_L g856 ( 
.A(n_700),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_677),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_677),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_677),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_677),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_569),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_622),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_677),
.Y(n_863)
);

CKINVDCx16_ASAP7_75t_R g864 ( 
.A(n_733),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_677),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_741),
.Y(n_866)
);

INVxp67_ASAP7_75t_SL g867 ( 
.A(n_622),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_517),
.B(n_1),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_741),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_573),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_741),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_741),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_668),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_741),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_646),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_741),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_741),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_613),
.Y(n_878)
);

INVxp67_ASAP7_75t_SL g879 ( 
.A(n_668),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_646),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_741),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_741),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_568),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_675),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_580),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_568),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_568),
.Y(n_887)
);

INVxp33_ASAP7_75t_SL g888 ( 
.A(n_675),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_568),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_568),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_568),
.Y(n_891)
);

CKINVDCx16_ASAP7_75t_R g892 ( 
.A(n_733),
.Y(n_892)
);

CKINVDCx14_ASAP7_75t_R g893 ( 
.A(n_564),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_604),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_604),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_604),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_624),
.Y(n_897)
);

INVxp67_ASAP7_75t_SL g898 ( 
.A(n_668),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_604),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_657),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_604),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_604),
.Y(n_902)
);

INVxp33_ASAP7_75t_L g903 ( 
.A(n_742),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_516),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_698),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_698),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_742),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_698),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_781),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_698),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_698),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_698),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_703),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_516),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_522),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_703),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_703),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_703),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_634),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_703),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_703),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_726),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_726),
.Y(n_923)
);

INVxp33_ASAP7_75t_L g924 ( 
.A(n_809),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_726),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_726),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_813),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_726),
.Y(n_928)
);

INVxp33_ASAP7_75t_SL g929 ( 
.A(n_809),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_726),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_796),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_796),
.Y(n_932)
);

INVxp67_ASAP7_75t_SL g933 ( 
.A(n_796),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_796),
.Y(n_934)
);

INVxp33_ASAP7_75t_SL g935 ( 
.A(n_519),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_814),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_796),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_796),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_536),
.Y(n_939)
);

INVxp33_ASAP7_75t_L g940 ( 
.A(n_517),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_536),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_590),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_590),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_835),
.B(n_1),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_596),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_801),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_827),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_520),
.Y(n_948)
);

BUFx2_ASAP7_75t_SL g949 ( 
.A(n_644),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_782),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_596),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_626),
.Y(n_952)
);

CKINVDCx14_ASAP7_75t_R g953 ( 
.A(n_523),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_626),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_662),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_662),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_666),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_666),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_671),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_525),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_818),
.Y(n_961)
);

INVxp33_ASAP7_75t_L g962 ( 
.A(n_518),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_671),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_587),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_650),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_521),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_810),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_810),
.Y(n_968)
);

CKINVDCx14_ASAP7_75t_R g969 ( 
.A(n_523),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_823),
.Y(n_970)
);

INVxp67_ASAP7_75t_SL g971 ( 
.A(n_801),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_782),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_535),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_650),
.Y(n_974)
);

INVxp33_ASAP7_75t_SL g975 ( 
.A(n_528),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_823),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_812),
.Y(n_977)
);

INVxp33_ASAP7_75t_L g978 ( 
.A(n_518),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_812),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_812),
.Y(n_980)
);

BUFx5_ASAP7_75t_L g981 ( 
.A(n_522),
.Y(n_981)
);

INVxp67_ASAP7_75t_SL g982 ( 
.A(n_701),
.Y(n_982)
);

INVxp33_ASAP7_75t_L g983 ( 
.A(n_524),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_524),
.Y(n_984)
);

INVxp33_ASAP7_75t_SL g985 ( 
.A(n_529),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_527),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_946),
.B(n_701),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_883),
.Y(n_988)
);

BUFx8_ASAP7_75t_SL g989 ( 
.A(n_973),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_888),
.A2(n_818),
.B1(n_832),
.B2(n_541),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_883),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_964),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_836),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_886),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_971),
.B(n_779),
.Y(n_995)
);

INVx5_ASAP7_75t_L g996 ( 
.A(n_964),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_929),
.A2(n_855),
.B1(n_884),
.B2(n_840),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_849),
.B(n_644),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_894),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_873),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_964),
.Y(n_1001)
);

INVx5_ASAP7_75t_L g1002 ( 
.A(n_964),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_886),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_852),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_964),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_894),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_906),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_893),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_861),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_935),
.B(n_975),
.Y(n_1010)
);

INVx5_ASAP7_75t_L g1011 ( 
.A(n_853),
.Y(n_1011)
);

OAI22x1_ASAP7_75t_R g1012 ( 
.A1(n_950),
.A2(n_603),
.B1(n_660),
.B2(n_572),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_906),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_853),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_873),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_878),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_933),
.B(n_566),
.Y(n_1017)
);

OA21x2_ASAP7_75t_L g1018 ( 
.A1(n_887),
.A2(n_577),
.B(n_566),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_863),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_887),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_863),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_885),
.Y(n_1022)
);

BUFx12f_ASAP7_75t_L g1023 ( 
.A(n_897),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_850),
.B(n_779),
.Y(n_1024)
);

AOI22x1_ASAP7_75t_SL g1025 ( 
.A1(n_972),
.A2(n_714),
.B1(n_721),
.B2(n_710),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_977),
.Y(n_1026)
);

INVx6_ASAP7_75t_L g1027 ( 
.A(n_981),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_900),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_850),
.B(n_802),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_889),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_881),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_889),
.Y(n_1032)
);

OA21x2_ASAP7_75t_L g1033 ( 
.A1(n_890),
.A2(n_895),
.B(n_891),
.Y(n_1033)
);

OA21x2_ASAP7_75t_L g1034 ( 
.A1(n_890),
.A2(n_632),
.B(n_577),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_944),
.A2(n_819),
.B1(n_588),
.B2(n_663),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_891),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_895),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_896),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_896),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_881),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_919),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_899),
.Y(n_1042)
);

BUFx8_ASAP7_75t_SL g1043 ( 
.A(n_880),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_899),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_909),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_977),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_901),
.Y(n_1047)
);

OA21x2_ASAP7_75t_L g1048 ( 
.A1(n_901),
.A2(n_712),
.B(n_632),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_846),
.B(n_712),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_902),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_862),
.B(n_724),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_979),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_903),
.A2(n_806),
.B1(n_533),
.B2(n_537),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_837),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_837),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_979),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_927),
.B(n_947),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_902),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_948),
.Y(n_1059)
);

INVx6_ASAP7_75t_L g1060 ( 
.A(n_981),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_905),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_905),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_908),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_908),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_980),
.Y(n_1065)
);

AND2x6_ASAP7_75t_L g1066 ( 
.A(n_838),
.B(n_587),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_864),
.A2(n_530),
.B1(n_542),
.B2(n_538),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_838),
.A2(n_751),
.B(n_724),
.Y(n_1068)
);

BUFx8_ASAP7_75t_SL g1069 ( 
.A(n_880),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_879),
.B(n_751),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_910),
.Y(n_1071)
);

OAI22x1_ASAP7_75t_R g1072 ( 
.A1(n_936),
.A2(n_548),
.B1(n_551),
.B2(n_550),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_892),
.A2(n_554),
.B1(n_555),
.B2(n_544),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_SL g1074 ( 
.A(n_961),
.B(n_523),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_898),
.B(n_802),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_910),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_960),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_911),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_911),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_912),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_985),
.A2(n_557),
.B1(n_558),
.B2(n_556),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_912),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_913),
.Y(n_1083)
);

OAI22x1_ASAP7_75t_L g1084 ( 
.A1(n_870),
.A2(n_579),
.B1(n_669),
.B2(n_656),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_913),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_981),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_867),
.B(n_783),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_916),
.Y(n_1088)
);

OA21x2_ASAP7_75t_L g1089 ( 
.A1(n_916),
.A2(n_798),
.B(n_783),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_949),
.B(n_798),
.Y(n_1090)
);

OAI22x1_ASAP7_75t_R g1091 ( 
.A1(n_966),
.A2(n_562),
.B1(n_570),
.B2(n_561),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_953),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_949),
.B(n_579),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_969),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_875),
.Y(n_1095)
);

BUFx12f_ASAP7_75t_L g1096 ( 
.A(n_868),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_917),
.Y(n_1097)
);

INVx6_ASAP7_75t_L g1098 ( 
.A(n_981),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_980),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_907),
.Y(n_1100)
);

BUFx8_ASAP7_75t_SL g1101 ( 
.A(n_904),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_917),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_918),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_918),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_920),
.Y(n_1105)
);

OA21x2_ASAP7_75t_L g1106 ( 
.A1(n_920),
.A2(n_834),
.B(n_833),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_921),
.Y(n_1107)
);

INVx5_ASAP7_75t_L g1108 ( 
.A(n_904),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_844),
.B(n_914),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_921),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_922),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_922),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_989),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_1092),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_1101),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_1022),
.Y(n_1116)
);

INVxp67_ASAP7_75t_SL g1117 ( 
.A(n_1015),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1026),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_1041),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1026),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1031),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1031),
.Y(n_1122)
);

NAND2xp33_ASAP7_75t_L g1123 ( 
.A(n_1066),
.B(n_587),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1026),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1031),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1046),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_992),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1046),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1046),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1052),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_1015),
.B(n_941),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_992),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_992),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_992),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1052),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_1095),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_1043),
.Y(n_1137)
);

INVxp67_ASAP7_75t_L g1138 ( 
.A(n_1074),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_993),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1052),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_R g1141 ( 
.A(n_1077),
.B(n_574),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_999),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1056),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1094),
.B(n_924),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1000),
.B(n_923),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_1004),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1056),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1009),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_1069),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_992),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_992),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1001),
.Y(n_1152)
);

CKINVDCx8_ASAP7_75t_R g1153 ( 
.A(n_1094),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1016),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_1028),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_1045),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1023),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_999),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1056),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1015),
.B(n_941),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1065),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1065),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1000),
.B(n_982),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_1012),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1001),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1023),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1023),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1065),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1099),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1099),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1099),
.B(n_943),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1024),
.B(n_965),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_1100),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1102),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1102),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1024),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1102),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_1096),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1054),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_997),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_1001),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1054),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1054),
.Y(n_1183)
);

INVxp33_ASAP7_75t_L g1184 ( 
.A(n_997),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1059),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_1017),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_999),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1054),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1001),
.Y(n_1189)
);

CKINVDCx20_ASAP7_75t_R g1190 ( 
.A(n_1012),
.Y(n_1190)
);

BUFx8_ASAP7_75t_L g1191 ( 
.A(n_1008),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1008),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_990),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_990),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1007),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1007),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_1029),
.Y(n_1197)
);

XNOR2xp5_ASAP7_75t_L g1198 ( 
.A(n_1025),
.B(n_856),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1055),
.Y(n_1199)
);

NAND2xp33_ASAP7_75t_L g1200 ( 
.A(n_1066),
.B(n_587),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1025),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1059),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1010),
.B(n_974),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_1072),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1055),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1001),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_1096),
.Y(n_1207)
);

CKINVDCx20_ASAP7_75t_R g1208 ( 
.A(n_1072),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1096),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1007),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1013),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_998),
.B(n_962),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_SL g1213 ( 
.A(n_1057),
.B(n_534),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1055),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_SL g1215 ( 
.A(n_1053),
.B(n_690),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1081),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1001),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1035),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1029),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1005),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1035),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1013),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1075),
.B(n_940),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1005),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1067),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1005),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1005),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1005),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_1073),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1075),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1055),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1005),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_987),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_987),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_995),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_1091),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_988),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_995),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_1091),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_988),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1070),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1013),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1084),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_991),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1019),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1084),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_991),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_994),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_1087),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_994),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1093),
.B(n_523),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1049),
.B(n_923),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1003),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1003),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1020),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1020),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1030),
.Y(n_1257)
);

BUFx12f_ASAP7_75t_L g1258 ( 
.A(n_1049),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1049),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1030),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1049),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1032),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1032),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1051),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1036),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1019),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1036),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1014),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1037),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1014),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1037),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1051),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1051),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1014),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1051),
.B(n_925),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1014),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1017),
.B(n_925),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1017),
.B(n_926),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1047),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1019),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1109),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1038),
.Y(n_1282)
);

OA21x2_ASAP7_75t_L g1283 ( 
.A1(n_1068),
.A2(n_841),
.B(n_839),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1047),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1047),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1038),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1039),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1068),
.A2(n_841),
.B(n_839),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_1090),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_1109),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1017),
.B(n_926),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1109),
.B(n_928),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1039),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1064),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1019),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1050),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1109),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1050),
.Y(n_1298)
);

INVx1_ASAP7_75t_SL g1299 ( 
.A(n_1106),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1019),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1061),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_R g1302 ( 
.A(n_1108),
.B(n_575),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1061),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1062),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1108),
.B(n_740),
.Y(n_1305)
);

OA21x2_ASAP7_75t_L g1306 ( 
.A1(n_1062),
.A2(n_843),
.B(n_842),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_1106),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1108),
.B(n_978),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1106),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1071),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1071),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1103),
.Y(n_1312)
);

NOR2xp67_ASAP7_75t_L g1313 ( 
.A(n_1108),
.B(n_915),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_R g1314 ( 
.A(n_1108),
.B(n_576),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_1019),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1021),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1064),
.Y(n_1317)
);

INVxp67_ASAP7_75t_L g1318 ( 
.A(n_1106),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1108),
.B(n_943),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1033),
.A2(n_843),
.B(n_842),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1018),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1064),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1103),
.Y(n_1323)
);

INVx6_ASAP7_75t_L g1324 ( 
.A(n_1042),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1104),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1104),
.B(n_983),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1105),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1105),
.B(n_954),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1112),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1112),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1042),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1042),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1066),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1042),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1042),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1021),
.B(n_928),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1076),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1066),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1241),
.B(n_704),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1186),
.Y(n_1340)
);

BUFx4f_ASAP7_75t_L g1341 ( 
.A(n_1258),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1306),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1306),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1306),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1307),
.A2(n_1018),
.B1(n_1048),
.B2(n_1034),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1121),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1186),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1121),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1122),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1259),
.B(n_587),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1307),
.A2(n_1018),
.B1(n_1048),
.B2(n_1034),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1122),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1125),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1125),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1264),
.B(n_1021),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1212),
.B(n_713),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1245),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1223),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1118),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1142),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1120),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1124),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1142),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1126),
.Y(n_1364)
);

NAND2xp33_ASAP7_75t_L g1365 ( 
.A(n_1259),
.B(n_587),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1163),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1128),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1261),
.B(n_766),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1158),
.Y(n_1369)
);

INVx8_ASAP7_75t_L g1370 ( 
.A(n_1258),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1158),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1113),
.Y(n_1372)
);

INVx4_ASAP7_75t_L g1373 ( 
.A(n_1245),
.Y(n_1373)
);

OR2x6_ASAP7_75t_L g1374 ( 
.A(n_1273),
.B(n_868),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1219),
.B(n_720),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1230),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1131),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1289),
.B(n_723),
.Y(n_1378)
);

INVx4_ASAP7_75t_L g1379 ( 
.A(n_1245),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1187),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1180),
.B(n_826),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1187),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1261),
.B(n_766),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1131),
.Y(n_1384)
);

INVx2_ASAP7_75t_SL g1385 ( 
.A(n_1131),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1318),
.A2(n_1033),
.B(n_1018),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1213),
.B(n_578),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1195),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1195),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1233),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1309),
.A2(n_1275),
.B(n_1252),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1272),
.B(n_766),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1160),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1196),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1129),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1264),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_SL g1397 ( 
.A(n_1160),
.Y(n_1397)
);

NAND2xp33_ASAP7_75t_SL g1398 ( 
.A(n_1229),
.B(n_1216),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1272),
.B(n_766),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1196),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1172),
.B(n_1089),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1171),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1171),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1171),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1174),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1210),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1210),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1211),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1115),
.Y(n_1409)
);

INVx4_ASAP7_75t_L g1410 ( 
.A(n_1245),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1175),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_1160),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1234),
.B(n_1235),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1177),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1211),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1321),
.A2(n_1218),
.B1(n_1221),
.B2(n_1215),
.Y(n_1416)
);

CKINVDCx6p67_ASAP7_75t_R g1417 ( 
.A(n_1137),
.Y(n_1417)
);

NAND2xp33_ASAP7_75t_SL g1418 ( 
.A(n_1216),
.B(n_656),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1130),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1222),
.Y(n_1420)
);

BUFx8_ASAP7_75t_SL g1421 ( 
.A(n_1137),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1179),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1245),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1176),
.B(n_1089),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1182),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1135),
.B(n_1021),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1222),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_1144),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1238),
.B(n_766),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1140),
.B(n_1143),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1242),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1242),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1147),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1183),
.Y(n_1434)
);

INVx8_ASAP7_75t_L g1435 ( 
.A(n_1321),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1173),
.Y(n_1436)
);

INVxp67_ASAP7_75t_SL g1437 ( 
.A(n_1266),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1266),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1266),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1188),
.Y(n_1440)
);

AOI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1218),
.A2(n_1089),
.B1(n_1034),
.B2(n_1048),
.Y(n_1441)
);

INVxp33_ASAP7_75t_SL g1442 ( 
.A(n_1136),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1159),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1199),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1205),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1281),
.B(n_766),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1214),
.Y(n_1447)
);

INVx2_ASAP7_75t_SL g1448 ( 
.A(n_1197),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1281),
.B(n_981),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1161),
.B(n_1021),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1279),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1325),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1290),
.B(n_981),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1221),
.A2(n_1089),
.B1(n_1034),
.B2(n_1048),
.Y(n_1454)
);

NAND2xp33_ASAP7_75t_SL g1455 ( 
.A(n_1141),
.B(n_669),
.Y(n_1455)
);

AND2x6_ASAP7_75t_L g1456 ( 
.A(n_1299),
.B(n_527),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1279),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1284),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_1119),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1266),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1231),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1284),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1162),
.B(n_1021),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1285),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1285),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1294),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1290),
.B(n_981),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1294),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1317),
.Y(n_1469)
);

BUFx10_ASAP7_75t_L g1470 ( 
.A(n_1114),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1266),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1317),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1322),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1322),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1337),
.Y(n_1475)
);

INVxp33_ASAP7_75t_L g1476 ( 
.A(n_1184),
.Y(n_1476)
);

BUFx4f_ASAP7_75t_L g1477 ( 
.A(n_1168),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1337),
.Y(n_1478)
);

OAI21xp33_ASAP7_75t_SL g1479 ( 
.A1(n_1251),
.A2(n_816),
.B(n_794),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1277),
.B(n_1033),
.C(n_847),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1320),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1320),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1237),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1240),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1249),
.A2(n_1033),
.B1(n_1066),
.B2(n_816),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1244),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1247),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1297),
.B(n_981),
.Y(n_1488)
);

CKINVDCx6p67_ASAP7_75t_R g1489 ( 
.A(n_1149),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1203),
.B(n_1138),
.Y(n_1490)
);

INVx4_ASAP7_75t_L g1491 ( 
.A(n_1280),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1248),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1250),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1253),
.Y(n_1494)
);

AND3x1_ASAP7_75t_L g1495 ( 
.A(n_1326),
.B(n_794),
.C(n_532),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1280),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1254),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1255),
.Y(n_1498)
);

OAI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1297),
.A2(n_532),
.B1(n_539),
.B2(n_531),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1256),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1169),
.B(n_1040),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1243),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1257),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1325),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1260),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1170),
.B(n_1040),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1262),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1263),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1280),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1265),
.Y(n_1510)
);

AND2x2_ASAP7_75t_SL g1511 ( 
.A(n_1123),
.B(n_531),
.Y(n_1511)
);

INVx5_ASAP7_75t_L g1512 ( 
.A(n_1280),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1308),
.B(n_1267),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1269),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_SL g1515 ( 
.A(n_1327),
.B(n_981),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1271),
.B(n_1040),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1280),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1282),
.Y(n_1518)
);

NOR2x1p5_ASAP7_75t_L g1519 ( 
.A(n_1207),
.B(n_539),
.Y(n_1519)
);

AOI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1249),
.A2(n_1066),
.B1(n_583),
.B2(n_585),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1286),
.Y(n_1521)
);

BUFx6f_ASAP7_75t_L g1522 ( 
.A(n_1295),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1287),
.Y(n_1523)
);

INVx4_ASAP7_75t_L g1524 ( 
.A(n_1295),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1293),
.Y(n_1525)
);

AND2x6_ASAP7_75t_L g1526 ( 
.A(n_1315),
.B(n_540),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1296),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1298),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1301),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1303),
.B(n_1040),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1304),
.B(n_1040),
.Y(n_1531)
);

NAND3xp33_ASAP7_75t_L g1532 ( 
.A(n_1278),
.B(n_847),
.C(n_845),
.Y(n_1532)
);

AND3x2_ASAP7_75t_L g1533 ( 
.A(n_1178),
.B(n_543),
.C(n_540),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1310),
.B(n_1040),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1291),
.A2(n_1066),
.B1(n_848),
.B2(n_851),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1311),
.B(n_1086),
.Y(n_1536)
);

INVx4_ASAP7_75t_L g1537 ( 
.A(n_1295),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1327),
.B(n_1329),
.Y(n_1538)
);

OAI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1225),
.A2(n_547),
.B1(n_549),
.B2(n_543),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1225),
.A2(n_1066),
.B1(n_589),
.B2(n_592),
.Y(n_1540)
);

INVx8_ASAP7_75t_L g1541 ( 
.A(n_1333),
.Y(n_1541)
);

BUFx4f_ASAP7_75t_L g1542 ( 
.A(n_1312),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1329),
.B(n_581),
.Y(n_1543)
);

OR2x6_ASAP7_75t_L g1544 ( 
.A(n_1292),
.B(n_547),
.Y(n_1544)
);

INVxp33_ASAP7_75t_L g1545 ( 
.A(n_1198),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1323),
.B(n_1086),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1243),
.B(n_984),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1330),
.Y(n_1548)
);

NOR2x1p5_ASAP7_75t_L g1549 ( 
.A(n_1207),
.B(n_549),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1328),
.Y(n_1550)
);

INVxp67_ASAP7_75t_L g1551 ( 
.A(n_1202),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1246),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1268),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1117),
.A2(n_848),
.B1(n_851),
.B2(n_845),
.Y(n_1554)
);

BUFx6f_ASAP7_75t_L g1555 ( 
.A(n_1295),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1145),
.B(n_1086),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1115),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1295),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1268),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1315),
.B(n_1086),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1288),
.Y(n_1561)
);

OR2x6_ASAP7_75t_L g1562 ( 
.A(n_1305),
.B(n_552),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1270),
.Y(n_1563)
);

INVx8_ASAP7_75t_L g1564 ( 
.A(n_1333),
.Y(n_1564)
);

NAND2xp33_ASAP7_75t_SL g1565 ( 
.A(n_1246),
.B(n_598),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1288),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1270),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1185),
.B(n_1202),
.Y(n_1568)
);

INVx5_ASAP7_75t_L g1569 ( 
.A(n_1300),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1139),
.B(n_593),
.Y(n_1570)
);

INVx4_ASAP7_75t_L g1571 ( 
.A(n_1300),
.Y(n_1571)
);

AOI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1336),
.A2(n_857),
.B(n_854),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1274),
.Y(n_1573)
);

AND2x6_ASAP7_75t_L g1574 ( 
.A(n_1315),
.B(n_552),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1274),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1283),
.B(n_984),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1139),
.B(n_595),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1146),
.B(n_597),
.Y(n_1578)
);

CKINVDCx6p67_ASAP7_75t_R g1579 ( 
.A(n_1149),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1276),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1146),
.B(n_600),
.Y(n_1581)
);

INVx2_ASAP7_75t_SL g1582 ( 
.A(n_1283),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1276),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1283),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1319),
.Y(n_1585)
);

INVx3_ASAP7_75t_L g1586 ( 
.A(n_1340),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1402),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1402),
.Y(n_1588)
);

INVxp33_ASAP7_75t_L g1589 ( 
.A(n_1568),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1403),
.Y(n_1590)
);

NOR2xp67_ASAP7_75t_L g1591 ( 
.A(n_1551),
.B(n_1148),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1366),
.B(n_1356),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1490),
.A2(n_1338),
.B1(n_1194),
.B2(n_1193),
.Y(n_1593)
);

AND2x6_ASAP7_75t_SL g1594 ( 
.A(n_1570),
.B(n_553),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1403),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1404),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1404),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1585),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1366),
.A2(n_1338),
.B1(n_1194),
.B2(n_1193),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_L g1600 ( 
.A(n_1522),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1378),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1585),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1346),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1339),
.B(n_1148),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_1522),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1396),
.B(n_1300),
.Y(n_1606)
);

NOR3xp33_ASAP7_75t_L g1607 ( 
.A(n_1387),
.B(n_1192),
.C(n_1155),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1515),
.A2(n_1154),
.B1(n_1156),
.B2(n_1155),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1346),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1396),
.B(n_1300),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1483),
.B(n_1300),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1347),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_SL g1613 ( 
.A(n_1470),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1476),
.B(n_1154),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1542),
.B(n_1156),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1348),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1370),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_L g1618 ( 
.A(n_1541),
.B(n_1209),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1483),
.B(n_1316),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1542),
.B(n_1340),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1428),
.B(n_1209),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1358),
.B(n_1153),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1542),
.B(n_1316),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1347),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1375),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1381),
.B(n_1153),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1375),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1486),
.B(n_1316),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1422),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1381),
.B(n_1114),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1522),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1348),
.Y(n_1632)
);

BUFx6f_ASAP7_75t_L g1633 ( 
.A(n_1522),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1486),
.B(n_1316),
.Y(n_1634)
);

BUFx3_ASAP7_75t_L g1635 ( 
.A(n_1370),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1340),
.B(n_1316),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1477),
.B(n_1192),
.Y(n_1637)
);

NAND3xp33_ASAP7_75t_L g1638 ( 
.A(n_1543),
.B(n_1416),
.C(n_1577),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1451),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1487),
.B(n_1134),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1370),
.Y(n_1641)
);

INVxp33_ASAP7_75t_L g1642 ( 
.A(n_1568),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1422),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1477),
.B(n_1331),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1487),
.B(n_1134),
.Y(n_1645)
);

NAND3xp33_ASAP7_75t_L g1646 ( 
.A(n_1416),
.B(n_1581),
.C(n_1578),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1492),
.B(n_1134),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1349),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1425),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1384),
.B(n_1119),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1477),
.B(n_1332),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1421),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1436),
.B(n_1116),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_1522),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1349),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1425),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1555),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_L g1658 ( 
.A(n_1372),
.B(n_1157),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1401),
.B(n_1334),
.Y(n_1659)
);

BUFx6f_ASAP7_75t_L g1660 ( 
.A(n_1555),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1492),
.B(n_1224),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1434),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1434),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1440),
.Y(n_1664)
);

BUFx6f_ASAP7_75t_L g1665 ( 
.A(n_1555),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1440),
.Y(n_1666)
);

NAND3xp33_ASAP7_75t_L g1667 ( 
.A(n_1538),
.B(n_1166),
.C(n_1157),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1452),
.B(n_1116),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1493),
.B(n_1228),
.Y(n_1669)
);

BUFx5_ASAP7_75t_L g1670 ( 
.A(n_1584),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1352),
.Y(n_1671)
);

CKINVDCx20_ASAP7_75t_R g1672 ( 
.A(n_1372),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1448),
.B(n_1166),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1555),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1444),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_SL g1676 ( 
.A(n_1442),
.B(n_1167),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1555),
.Y(n_1677)
);

BUFx6f_ASAP7_75t_L g1678 ( 
.A(n_1558),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1493),
.B(n_1228),
.Y(n_1679)
);

NAND2x1_ASAP7_75t_L g1680 ( 
.A(n_1373),
.B(n_1217),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1352),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1444),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1376),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1494),
.B(n_1228),
.Y(n_1684)
);

OR2x6_ASAP7_75t_L g1685 ( 
.A(n_1370),
.B(n_1191),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1448),
.B(n_1452),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1353),
.Y(n_1687)
);

AOI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1401),
.A2(n_1385),
.B1(n_1393),
.B2(n_1377),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1353),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1494),
.B(n_1232),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1456),
.A2(n_559),
.B1(n_560),
.B2(n_553),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1497),
.B(n_1232),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1504),
.B(n_1167),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1445),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1445),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1504),
.B(n_1335),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1558),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_SL g1698 ( 
.A(n_1424),
.B(n_1127),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1447),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1447),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1461),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1376),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1497),
.B(n_1217),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1424),
.B(n_1127),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1370),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1461),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1377),
.B(n_1385),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1374),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1390),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1393),
.B(n_1127),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1412),
.B(n_1127),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1547),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1498),
.B(n_1217),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1498),
.B(n_1224),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1503),
.B(n_1224),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1503),
.B(n_1232),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1412),
.B(n_1127),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1485),
.B(n_1132),
.Y(n_1718)
);

BUFx6f_ASAP7_75t_L g1719 ( 
.A(n_1558),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1384),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1451),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1485),
.B(n_1132),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_1547),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1354),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1523),
.B(n_1132),
.Y(n_1725)
);

INVxp67_ASAP7_75t_L g1726 ( 
.A(n_1390),
.Y(n_1726)
);

INVx4_ASAP7_75t_L g1727 ( 
.A(n_1397),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1413),
.B(n_1513),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1374),
.B(n_1236),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1354),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1456),
.A2(n_560),
.B1(n_563),
.B2(n_559),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1523),
.B(n_1132),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1405),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1525),
.B(n_1548),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1525),
.B(n_1132),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1374),
.B(n_1236),
.Y(n_1736)
);

NOR3xp33_ASAP7_75t_L g1737 ( 
.A(n_1398),
.B(n_1201),
.C(n_606),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1548),
.B(n_1133),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1484),
.B(n_1133),
.Y(n_1739)
);

INVxp67_ASAP7_75t_L g1740 ( 
.A(n_1418),
.Y(n_1740)
);

BUFx6f_ASAP7_75t_L g1741 ( 
.A(n_1558),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1360),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1405),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1457),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1374),
.B(n_1239),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1484),
.B(n_1133),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1411),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_SL g1748 ( 
.A(n_1470),
.Y(n_1748)
);

AO221x1_ASAP7_75t_L g1749 ( 
.A1(n_1539),
.A2(n_567),
.B1(n_571),
.B2(n_565),
.C(n_563),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1374),
.B(n_1239),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1533),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1500),
.B(n_1133),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1411),
.Y(n_1753)
);

BUFx5_ASAP7_75t_L g1754 ( 
.A(n_1584),
.Y(n_1754)
);

NAND2xp33_ASAP7_75t_L g1755 ( 
.A(n_1541),
.B(n_1302),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_SL g1756 ( 
.A(n_1558),
.B(n_1133),
.Y(n_1756)
);

NAND3xp33_ASAP7_75t_L g1757 ( 
.A(n_1520),
.B(n_1191),
.C(n_1201),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1414),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1536),
.B(n_1150),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1546),
.B(n_1150),
.Y(n_1760)
);

XOR2xp5_ASAP7_75t_L g1761 ( 
.A(n_1409),
.B(n_1557),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1414),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1576),
.B(n_1150),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1360),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1500),
.B(n_1150),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1455),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1359),
.Y(n_1767)
);

BUFx6f_ASAP7_75t_SL g1768 ( 
.A(n_1470),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1359),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1505),
.B(n_1150),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1550),
.B(n_1164),
.Y(n_1771)
);

NOR2xp67_ASAP7_75t_L g1772 ( 
.A(n_1409),
.B(n_986),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1550),
.B(n_601),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1363),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1363),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1361),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1361),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1369),
.Y(n_1778)
);

NAND2xp33_ASAP7_75t_L g1779 ( 
.A(n_1541),
.B(n_1314),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1362),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1362),
.Y(n_1781)
);

NOR2xp67_ASAP7_75t_L g1782 ( 
.A(n_1557),
.B(n_986),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1369),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1505),
.B(n_1151),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1576),
.B(n_1151),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1364),
.Y(n_1786)
);

NAND2xp33_ASAP7_75t_L g1787 ( 
.A(n_1541),
.B(n_1151),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1371),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1507),
.B(n_1151),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1520),
.B(n_608),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_R g1791 ( 
.A(n_1565),
.B(n_1164),
.Y(n_1791)
);

NOR3xp33_ASAP7_75t_L g1792 ( 
.A(n_1479),
.B(n_612),
.C(n_609),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1417),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1364),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1507),
.B(n_1151),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_L g1796 ( 
.A(n_1540),
.B(n_1191),
.C(n_1204),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1457),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1419),
.Y(n_1798)
);

NOR2xp67_ASAP7_75t_L g1799 ( 
.A(n_1540),
.B(n_1319),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1458),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1508),
.B(n_1152),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1508),
.B(n_1152),
.Y(n_1802)
);

BUFx6f_ASAP7_75t_SL g1803 ( 
.A(n_1470),
.Y(n_1803)
);

AOI221x1_ASAP7_75t_L g1804 ( 
.A1(n_1367),
.A2(n_932),
.B1(n_934),
.B2(n_931),
.C(n_930),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1433),
.B(n_615),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1510),
.B(n_1152),
.Y(n_1806)
);

INVxp67_ASAP7_75t_L g1807 ( 
.A(n_1502),
.Y(n_1807)
);

INVxp67_ASAP7_75t_L g1808 ( 
.A(n_1502),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_SL g1809 ( 
.A(n_1510),
.B(n_1152),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1367),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1395),
.Y(n_1811)
);

AOI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1499),
.A2(n_571),
.B1(n_582),
.B2(n_567),
.C(n_565),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1514),
.B(n_1152),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1514),
.B(n_1165),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1518),
.B(n_1165),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1544),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1518),
.B(n_1521),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1521),
.B(n_1165),
.Y(n_1818)
);

NOR2xp67_ASAP7_75t_L g1819 ( 
.A(n_1527),
.B(n_1319),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1527),
.B(n_1528),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1371),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1528),
.B(n_1165),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1395),
.Y(n_1823)
);

NOR3xp33_ASAP7_75t_L g1824 ( 
.A(n_1479),
.B(n_617),
.C(n_616),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1433),
.B(n_618),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_L g1826 ( 
.A(n_1443),
.B(n_620),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_SL g1827 ( 
.A(n_1442),
.B(n_1204),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1380),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1529),
.B(n_1165),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1553),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1529),
.B(n_1181),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1443),
.B(n_621),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1670),
.B(n_1391),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1587),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1588),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1638),
.B(n_1341),
.Y(n_1836)
);

INVxp67_ASAP7_75t_L g1837 ( 
.A(n_1627),
.Y(n_1837)
);

AO22x2_ASAP7_75t_L g1838 ( 
.A1(n_1646),
.A2(n_1459),
.B1(n_1429),
.B2(n_1495),
.Y(n_1838)
);

INVx1_ASAP7_75t_SL g1839 ( 
.A(n_1702),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1595),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1597),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1598),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1639),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1670),
.B(n_1391),
.Y(n_1844)
);

NAND2x1p5_ASAP7_75t_L g1845 ( 
.A(n_1617),
.B(n_1373),
.Y(n_1845)
);

BUFx6f_ASAP7_75t_L g1846 ( 
.A(n_1617),
.Y(n_1846)
);

CKINVDCx20_ASAP7_75t_R g1847 ( 
.A(n_1672),
.Y(n_1847)
);

NOR2x1p5_ASAP7_75t_L g1848 ( 
.A(n_1757),
.B(n_1417),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1602),
.Y(n_1849)
);

AO22x2_ASAP7_75t_L g1850 ( 
.A1(n_1796),
.A2(n_1495),
.B1(n_584),
.B2(n_586),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1590),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1670),
.B(n_1391),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1596),
.Y(n_1853)
);

AO22x2_ASAP7_75t_L g1854 ( 
.A1(n_1601),
.A2(n_584),
.B1(n_586),
.B2(n_582),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1830),
.Y(n_1855)
);

CKINVDCx20_ASAP7_75t_R g1856 ( 
.A(n_1652),
.Y(n_1856)
);

INVx2_ASAP7_75t_SL g1857 ( 
.A(n_1712),
.Y(n_1857)
);

AO22x2_ASAP7_75t_L g1858 ( 
.A1(n_1723),
.A2(n_594),
.B1(n_599),
.B2(n_591),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1639),
.Y(n_1859)
);

AO22x2_ASAP7_75t_L g1860 ( 
.A1(n_1733),
.A2(n_594),
.B1(n_599),
.B2(n_591),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1629),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1643),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1649),
.Y(n_1863)
);

BUFx2_ASAP7_75t_L g1864 ( 
.A(n_1650),
.Y(n_1864)
);

CKINVDCx16_ASAP7_75t_R g1865 ( 
.A(n_1827),
.Y(n_1865)
);

AO22x2_ASAP7_75t_L g1866 ( 
.A1(n_1743),
.A2(n_605),
.B1(n_607),
.B2(n_602),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1656),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1662),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1670),
.B(n_1456),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1663),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1664),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1670),
.B(n_1456),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1666),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1670),
.B(n_1456),
.Y(n_1874)
);

AO22x2_ASAP7_75t_L g1875 ( 
.A1(n_1747),
.A2(n_605),
.B1(n_607),
.B2(n_602),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1721),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1721),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1744),
.Y(n_1878)
);

OR2x6_ASAP7_75t_L g1879 ( 
.A(n_1685),
.B(n_1435),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1675),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1604),
.B(n_1552),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1604),
.B(n_1552),
.Y(n_1882)
);

AO22x2_ASAP7_75t_L g1883 ( 
.A1(n_1753),
.A2(n_1758),
.B1(n_1767),
.B2(n_1762),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1682),
.Y(n_1884)
);

AO22x2_ASAP7_75t_L g1885 ( 
.A1(n_1769),
.A2(n_611),
.B1(n_625),
.B2(n_610),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1694),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1695),
.Y(n_1887)
);

INVx4_ASAP7_75t_L g1888 ( 
.A(n_1798),
.Y(n_1888)
);

OR2x6_ASAP7_75t_L g1889 ( 
.A(n_1685),
.B(n_1435),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1728),
.A2(n_1435),
.B1(n_1456),
.B2(n_1544),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1699),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1744),
.Y(n_1892)
);

BUFx2_ASAP7_75t_L g1893 ( 
.A(n_1650),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1700),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1701),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1706),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1793),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1776),
.Y(n_1898)
);

AO22x2_ASAP7_75t_L g1899 ( 
.A1(n_1777),
.A2(n_611),
.B1(n_625),
.B2(n_610),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1797),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1780),
.Y(n_1901)
);

AO22x2_ASAP7_75t_L g1902 ( 
.A1(n_1781),
.A2(n_629),
.B1(n_631),
.B2(n_627),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1786),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1625),
.B(n_1519),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1630),
.B(n_1626),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1794),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1810),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1811),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1797),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1592),
.B(n_1341),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1823),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1820),
.Y(n_1912)
);

AOI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1728),
.A2(n_1435),
.B1(n_1456),
.B2(n_1544),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1800),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1800),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1626),
.B(n_1341),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1754),
.B(n_1342),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1754),
.B(n_1342),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1603),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1754),
.B(n_1343),
.Y(n_1920)
);

BUFx6f_ASAP7_75t_SL g1921 ( 
.A(n_1685),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1754),
.B(n_1343),
.Y(n_1922)
);

NOR2xp67_ASAP7_75t_L g1923 ( 
.A(n_1734),
.B(n_1480),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1635),
.B(n_1419),
.Y(n_1924)
);

INVxp67_ASAP7_75t_SL g1925 ( 
.A(n_1754),
.Y(n_1925)
);

AO22x2_ASAP7_75t_L g1926 ( 
.A1(n_1637),
.A2(n_629),
.B1(n_631),
.B2(n_627),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1612),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1754),
.B(n_1344),
.Y(n_1928)
);

AO22x2_ASAP7_75t_L g1929 ( 
.A1(n_1637),
.A2(n_649),
.B1(n_651),
.B2(n_636),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1624),
.Y(n_1930)
);

CKINVDCx20_ASAP7_75t_R g1931 ( 
.A(n_1761),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1609),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1616),
.Y(n_1933)
);

NOR2xp67_ASAP7_75t_L g1934 ( 
.A(n_1586),
.B(n_1766),
.Y(n_1934)
);

INVx3_ASAP7_75t_L g1935 ( 
.A(n_1798),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1632),
.Y(n_1936)
);

BUFx8_ASAP7_75t_L g1937 ( 
.A(n_1613),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1648),
.Y(n_1938)
);

INVx3_ASAP7_75t_L g1939 ( 
.A(n_1798),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1655),
.Y(n_1940)
);

AO22x2_ASAP7_75t_L g1941 ( 
.A1(n_1718),
.A2(n_649),
.B1(n_651),
.B2(n_636),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1671),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1681),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1586),
.B(n_1344),
.Y(n_1944)
);

AO22x2_ASAP7_75t_L g1945 ( 
.A1(n_1718),
.A2(n_655),
.B1(n_658),
.B2(n_654),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1686),
.B(n_1435),
.Y(n_1946)
);

NAND2x1p5_ASAP7_75t_L g1947 ( 
.A(n_1635),
.B(n_1373),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1687),
.Y(n_1948)
);

AOI22xp33_ASAP7_75t_L g1949 ( 
.A1(n_1790),
.A2(n_1544),
.B1(n_1419),
.B2(n_1397),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1653),
.B(n_1430),
.Y(n_1950)
);

INVxp67_ASAP7_75t_L g1951 ( 
.A(n_1686),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1689),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1724),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1630),
.B(n_1545),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1668),
.B(n_1519),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1641),
.B(n_1705),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1730),
.Y(n_1957)
);

INVxp33_ASAP7_75t_L g1958 ( 
.A(n_1614),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1742),
.Y(n_1959)
);

AOI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1790),
.A2(n_1544),
.B1(n_1554),
.B2(n_1526),
.Y(n_1960)
);

AO22x2_ASAP7_75t_L g1961 ( 
.A1(n_1722),
.A2(n_655),
.B1(n_658),
.B2(n_654),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1764),
.Y(n_1962)
);

BUFx8_ASAP7_75t_L g1963 ( 
.A(n_1613),
.Y(n_1963)
);

OAI221xp5_ASAP7_75t_L g1964 ( 
.A1(n_1691),
.A2(n_673),
.B1(n_679),
.B2(n_672),
.C(n_665),
.Y(n_1964)
);

AND2x4_ASAP7_75t_L g1965 ( 
.A(n_1641),
.B(n_1549),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1774),
.Y(n_1966)
);

OAI21xp33_ASAP7_75t_L g1967 ( 
.A1(n_1691),
.A2(n_1454),
.B(n_1441),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1817),
.B(n_1582),
.Y(n_1968)
);

AO22x2_ASAP7_75t_L g1969 ( 
.A1(n_1722),
.A2(n_672),
.B1(n_673),
.B2(n_665),
.Y(n_1969)
);

AO22x2_ASAP7_75t_L g1970 ( 
.A1(n_1607),
.A2(n_680),
.B1(n_681),
.B2(n_679),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1608),
.B(n_1467),
.Y(n_1971)
);

AO22x2_ASAP7_75t_L g1972 ( 
.A1(n_1615),
.A2(n_681),
.B1(n_684),
.B2(n_680),
.Y(n_1972)
);

AOI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1817),
.A2(n_1574),
.B1(n_1526),
.B2(n_1453),
.Y(n_1973)
);

AO22x2_ASAP7_75t_L g1974 ( 
.A1(n_1615),
.A2(n_685),
.B1(n_687),
.B2(n_684),
.Y(n_1974)
);

AO22x2_ASAP7_75t_L g1975 ( 
.A1(n_1807),
.A2(n_1808),
.B1(n_1824),
.B2(n_1792),
.Y(n_1975)
);

NAND2x1p5_ASAP7_75t_L g1976 ( 
.A(n_1705),
.B(n_1373),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1775),
.Y(n_1977)
);

NAND2x1p5_ASAP7_75t_L g1978 ( 
.A(n_1798),
.B(n_1379),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1727),
.B(n_1549),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1591),
.B(n_1449),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1621),
.B(n_1589),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1642),
.B(n_1562),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1659),
.B(n_1582),
.Y(n_1983)
);

INVx3_ASAP7_75t_L g1984 ( 
.A(n_1600),
.Y(n_1984)
);

AO22x2_ASAP7_75t_L g1985 ( 
.A1(n_1696),
.A2(n_1771),
.B1(n_1720),
.B2(n_1804),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1778),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1783),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1788),
.Y(n_1988)
);

AO22x2_ASAP7_75t_L g1989 ( 
.A1(n_1696),
.A2(n_687),
.B1(n_689),
.B2(n_685),
.Y(n_1989)
);

CKINVDCx20_ASAP7_75t_R g1990 ( 
.A(n_1791),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1821),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1828),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1659),
.B(n_1541),
.Y(n_1993)
);

AO22x2_ASAP7_75t_L g1994 ( 
.A1(n_1667),
.A2(n_691),
.B1(n_696),
.B2(n_689),
.Y(n_1994)
);

AOI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1688),
.A2(n_1526),
.B1(n_1574),
.B2(n_1488),
.Y(n_1995)
);

OAI22xp33_ASAP7_75t_L g1996 ( 
.A1(n_1593),
.A2(n_1816),
.B1(n_1599),
.B2(n_1799),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1698),
.B(n_1564),
.Y(n_1997)
);

AND2x4_ASAP7_75t_L g1998 ( 
.A(n_1727),
.B(n_1708),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1622),
.B(n_1564),
.Y(n_1999)
);

CKINVDCx20_ASAP7_75t_R g2000 ( 
.A(n_1791),
.Y(n_2000)
);

AO22x2_ASAP7_75t_L g2001 ( 
.A1(n_1683),
.A2(n_696),
.B1(n_697),
.B2(n_691),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1622),
.B(n_1562),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1698),
.B(n_1564),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1640),
.Y(n_2004)
);

AO22x2_ASAP7_75t_L g2005 ( 
.A1(n_1709),
.A2(n_711),
.B1(n_719),
.B2(n_697),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1645),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1647),
.Y(n_2007)
);

AO22x2_ASAP7_75t_L g2008 ( 
.A1(n_1726),
.A2(n_719),
.B1(n_725),
.B2(n_711),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1661),
.Y(n_2009)
);

AO22x2_ASAP7_75t_L g2010 ( 
.A1(n_1737),
.A2(n_1623),
.B1(n_1704),
.B2(n_1740),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1669),
.Y(n_2011)
);

NOR2xp67_ASAP7_75t_L g2012 ( 
.A(n_1620),
.B(n_1480),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1679),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1684),
.Y(n_2014)
);

NAND2x1p5_ASAP7_75t_L g2015 ( 
.A(n_1600),
.B(n_1605),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1690),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1692),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1703),
.Y(n_2018)
);

AO22x2_ASAP7_75t_L g2019 ( 
.A1(n_1623),
.A2(n_727),
.B1(n_729),
.B2(n_725),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1713),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1714),
.Y(n_2021)
);

HB1xp67_ASAP7_75t_L g2022 ( 
.A(n_1600),
.Y(n_2022)
);

AO22x2_ASAP7_75t_L g2023 ( 
.A1(n_1704),
.A2(n_729),
.B1(n_734),
.B2(n_727),
.Y(n_2023)
);

NOR2xp67_ASAP7_75t_L g2024 ( 
.A(n_1620),
.B(n_1532),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1773),
.B(n_1562),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_1748),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1715),
.Y(n_2027)
);

NOR2xp67_ASAP7_75t_L g2028 ( 
.A(n_1819),
.B(n_1532),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1716),
.Y(n_2029)
);

AO22x2_ASAP7_75t_L g2030 ( 
.A1(n_1763),
.A2(n_737),
.B1(n_738),
.B2(n_734),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1739),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1746),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1725),
.Y(n_2033)
);

AND2x4_ASAP7_75t_L g2034 ( 
.A(n_1751),
.B(n_1562),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1752),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1732),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1614),
.B(n_1190),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1735),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1738),
.Y(n_2039)
);

AND2x2_ASAP7_75t_SL g2040 ( 
.A(n_1618),
.B(n_1511),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1611),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_1693),
.B(n_1190),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_SL g2043 ( 
.A(n_1693),
.B(n_1564),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1619),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1847),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1905),
.B(n_1773),
.Y(n_2046)
);

CKINVDCx11_ASAP7_75t_R g2047 ( 
.A(n_1856),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1843),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_1958),
.B(n_1676),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_2025),
.B(n_1628),
.Y(n_2050)
);

AOI21xp5_ASAP7_75t_L g2051 ( 
.A1(n_1925),
.A2(n_1787),
.B(n_2043),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_L g2052 ( 
.A(n_1881),
.B(n_1805),
.Y(n_2052)
);

OAI21xp5_ASAP7_75t_L g2053 ( 
.A1(n_2012),
.A2(n_1707),
.B(n_1651),
.Y(n_2053)
);

OAI21xp33_ASAP7_75t_L g2054 ( 
.A1(n_1882),
.A2(n_1825),
.B(n_1805),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1859),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1951),
.B(n_1825),
.Y(n_2056)
);

AOI21xp5_ASAP7_75t_L g2057 ( 
.A1(n_1925),
.A2(n_1410),
.B(n_1379),
.Y(n_2057)
);

NAND3xp33_ASAP7_75t_L g2058 ( 
.A(n_1954),
.B(n_2042),
.C(n_1832),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1865),
.B(n_1673),
.Y(n_2059)
);

AOI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_1917),
.A2(n_1410),
.B(n_1379),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1917),
.A2(n_1410),
.B(n_1379),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1876),
.Y(n_2062)
);

OAI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_1949),
.A2(n_1564),
.B1(n_1673),
.B2(n_1634),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_1918),
.A2(n_1438),
.B(n_1410),
.Y(n_2064)
);

NOR3xp33_ASAP7_75t_SL g2065 ( 
.A(n_1836),
.B(n_1736),
.C(n_1729),
.Y(n_2065)
);

AOI21x1_ASAP7_75t_L g2066 ( 
.A1(n_1946),
.A2(n_1760),
.B(n_1759),
.Y(n_2066)
);

INVxp67_ASAP7_75t_L g2067 ( 
.A(n_1839),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_L g2068 ( 
.A(n_1951),
.B(n_1826),
.Y(n_2068)
);

A2O1A1Ixp33_ASAP7_75t_L g2069 ( 
.A1(n_1960),
.A2(n_1832),
.B(n_1826),
.C(n_1772),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1912),
.B(n_1782),
.Y(n_2070)
);

OAI21x1_ASAP7_75t_L g2071 ( 
.A1(n_1869),
.A2(n_1760),
.B(n_1759),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1981),
.B(n_1729),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_2002),
.B(n_1950),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_1998),
.B(n_1658),
.Y(n_2074)
);

BUFx4f_ASAP7_75t_L g2075 ( 
.A(n_1879),
.Y(n_2075)
);

AOI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1918),
.A2(n_1491),
.B(n_1438),
.Y(n_2076)
);

INVxp67_ASAP7_75t_L g2077 ( 
.A(n_1839),
.Y(n_2077)
);

AOI21xp5_ASAP7_75t_L g2078 ( 
.A1(n_1920),
.A2(n_1491),
.B(n_1438),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1955),
.B(n_1736),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1883),
.Y(n_2080)
);

AOI21xp5_ASAP7_75t_L g2081 ( 
.A1(n_1920),
.A2(n_1491),
.B(n_1438),
.Y(n_2081)
);

INVx3_ASAP7_75t_L g2082 ( 
.A(n_1845),
.Y(n_2082)
);

AOI21xp5_ASAP7_75t_L g2083 ( 
.A1(n_1922),
.A2(n_1524),
.B(n_1491),
.Y(n_2083)
);

AOI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_1922),
.A2(n_1537),
.B(n_1524),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_SL g2085 ( 
.A(n_1996),
.B(n_1837),
.Y(n_2085)
);

OAI22xp5_ASAP7_75t_L g2086 ( 
.A1(n_1890),
.A2(n_1610),
.B1(n_1606),
.B2(n_1707),
.Y(n_2086)
);

AOI21xp5_ASAP7_75t_L g2087 ( 
.A1(n_1928),
.A2(n_1537),
.B(n_1524),
.Y(n_2087)
);

O2A1O1Ixp33_ASAP7_75t_L g2088 ( 
.A1(n_1916),
.A2(n_1910),
.B(n_1996),
.C(n_1971),
.Y(n_2088)
);

AOI21x1_ASAP7_75t_L g2089 ( 
.A1(n_1999),
.A2(n_1651),
.B(n_1644),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2033),
.B(n_1731),
.Y(n_2090)
);

INVx4_ASAP7_75t_L g2091 ( 
.A(n_1846),
.Y(n_2091)
);

AOI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_1928),
.A2(n_1537),
.B(n_1524),
.Y(n_2092)
);

AOI33xp33_ASAP7_75t_L g2093 ( 
.A1(n_1904),
.A2(n_1812),
.A3(n_1731),
.B1(n_746),
.B2(n_738),
.B3(n_748),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1883),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_2036),
.B(n_1749),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1861),
.Y(n_2096)
);

A2O1A1Ixp33_ASAP7_75t_L g2097 ( 
.A1(n_1960),
.A2(n_1967),
.B(n_1913),
.C(n_1890),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1913),
.B(n_1644),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2038),
.B(n_1763),
.Y(n_2099)
);

AOI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_1833),
.A2(n_1571),
.B(n_1537),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_1998),
.B(n_1710),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2039),
.B(n_1785),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_SL g2103 ( 
.A(n_1923),
.B(n_1600),
.Y(n_2103)
);

OAI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_1964),
.A2(n_1208),
.B1(n_1750),
.B2(n_1745),
.Y(n_2104)
);

AOI21x1_ASAP7_75t_L g2105 ( 
.A1(n_1869),
.A2(n_1795),
.B(n_1789),
.Y(n_2105)
);

AOI22xp5_ASAP7_75t_L g2106 ( 
.A1(n_2037),
.A2(n_1208),
.B1(n_1750),
.B2(n_1745),
.Y(n_2106)
);

OAI21x1_ASAP7_75t_L g2107 ( 
.A1(n_1872),
.A2(n_1818),
.B(n_1770),
.Y(n_2107)
);

AOI21xp5_ASAP7_75t_L g2108 ( 
.A1(n_1833),
.A2(n_1571),
.B(n_1844),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2041),
.B(n_1785),
.Y(n_2109)
);

HB1xp67_ASAP7_75t_L g2110 ( 
.A(n_2022),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_1982),
.B(n_1864),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2044),
.B(n_1350),
.Y(n_2112)
);

NOR2xp33_ASAP7_75t_L g2113 ( 
.A(n_1837),
.B(n_1594),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2004),
.B(n_1368),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1877),
.Y(n_2115)
);

AOI22x1_ASAP7_75t_L g2116 ( 
.A1(n_2010),
.A2(n_1475),
.B1(n_1478),
.B2(n_1437),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2006),
.B(n_2007),
.Y(n_2117)
);

AOI21xp5_ASAP7_75t_L g2118 ( 
.A1(n_1844),
.A2(n_1571),
.B(n_1755),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_1893),
.B(n_1562),
.Y(n_2119)
);

BUFx2_ASAP7_75t_L g2120 ( 
.A(n_1857),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1862),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2009),
.B(n_1383),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_L g2123 ( 
.A(n_1863),
.B(n_1392),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2011),
.B(n_1399),
.Y(n_2124)
);

A2O1A1Ixp33_ASAP7_75t_L g2125 ( 
.A1(n_1967),
.A2(n_1365),
.B(n_1446),
.C(n_1779),
.Y(n_2125)
);

AOI21xp5_ASAP7_75t_L g2126 ( 
.A1(n_1852),
.A2(n_1571),
.B(n_1569),
.Y(n_2126)
);

AO21x1_ASAP7_75t_L g2127 ( 
.A1(n_1872),
.A2(n_1795),
.B(n_1789),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2013),
.B(n_1345),
.Y(n_2128)
);

INVxp67_ASAP7_75t_L g2129 ( 
.A(n_1867),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2014),
.B(n_1351),
.Y(n_2130)
);

NOR2xp33_ASAP7_75t_L g2131 ( 
.A(n_1868),
.B(n_1748),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_SL g2132 ( 
.A(n_2034),
.B(n_1605),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2016),
.B(n_1765),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2017),
.B(n_1784),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_2020),
.B(n_1801),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_L g2136 ( 
.A(n_1870),
.B(n_1768),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1871),
.Y(n_2137)
);

NOR2xp33_ASAP7_75t_L g2138 ( 
.A(n_1873),
.B(n_1768),
.Y(n_2138)
);

NAND2x1p5_ASAP7_75t_L g2139 ( 
.A(n_1956),
.B(n_1605),
.Y(n_2139)
);

AND2x4_ASAP7_75t_L g2140 ( 
.A(n_1965),
.B(n_1710),
.Y(n_2140)
);

AOI21xp5_ASAP7_75t_L g2141 ( 
.A1(n_1852),
.A2(n_1569),
.B(n_1512),
.Y(n_2141)
);

O2A1O1Ixp33_ASAP7_75t_L g2142 ( 
.A1(n_1980),
.A2(n_1822),
.B(n_1829),
.C(n_1809),
.Y(n_2142)
);

AOI21xp5_ASAP7_75t_L g2143 ( 
.A1(n_1993),
.A2(n_1569),
.B(n_1512),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2021),
.B(n_1802),
.Y(n_2144)
);

AOI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_1993),
.A2(n_1569),
.B(n_1512),
.Y(n_2145)
);

NOR3xp33_ASAP7_75t_L g2146 ( 
.A(n_1964),
.B(n_1530),
.C(n_1516),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1878),
.Y(n_2147)
);

OAI321xp33_ASAP7_75t_L g2148 ( 
.A1(n_1927),
.A2(n_747),
.A3(n_746),
.B1(n_749),
.B2(n_748),
.C(n_737),
.Y(n_2148)
);

INVx6_ASAP7_75t_L g2149 ( 
.A(n_1846),
.Y(n_2149)
);

AOI21xp5_ASAP7_75t_L g2150 ( 
.A1(n_1997),
.A2(n_1569),
.B(n_1512),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1880),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1892),
.Y(n_2152)
);

AOI33xp33_ASAP7_75t_L g2153 ( 
.A1(n_1884),
.A2(n_753),
.A3(n_747),
.B1(n_758),
.B2(n_756),
.B3(n_749),
.Y(n_2153)
);

NOR2xp33_ASAP7_75t_L g2154 ( 
.A(n_1886),
.B(n_1803),
.Y(n_2154)
);

OAI21xp5_ASAP7_75t_L g2155 ( 
.A1(n_2012),
.A2(n_1355),
.B(n_1806),
.Y(n_2155)
);

NOR2xp33_ASAP7_75t_L g2156 ( 
.A(n_1887),
.B(n_1803),
.Y(n_2156)
);

BUFx12f_ASAP7_75t_L g2157 ( 
.A(n_1937),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2027),
.B(n_1813),
.Y(n_2158)
);

BUFx3_ASAP7_75t_L g2159 ( 
.A(n_1937),
.Y(n_2159)
);

INVx6_ASAP7_75t_L g2160 ( 
.A(n_1846),
.Y(n_2160)
);

BUFx8_ASAP7_75t_L g2161 ( 
.A(n_1921),
.Y(n_2161)
);

AO22x1_ASAP7_75t_L g2162 ( 
.A1(n_1965),
.A2(n_628),
.B1(n_630),
.B2(n_623),
.Y(n_2162)
);

A2O1A1Ixp33_ASAP7_75t_L g2163 ( 
.A1(n_2024),
.A2(n_1717),
.B(n_1711),
.C(n_1814),
.Y(n_2163)
);

O2A1O1Ixp5_ASAP7_75t_L g2164 ( 
.A1(n_1874),
.A2(n_1822),
.B(n_1829),
.C(n_1809),
.Y(n_2164)
);

O2A1O1Ixp5_ASAP7_75t_SL g2165 ( 
.A1(n_1855),
.A2(n_1831),
.B(n_753),
.C(n_758),
.Y(n_2165)
);

OAI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_2040),
.A2(n_1815),
.B1(n_1741),
.B2(n_1719),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_SL g2167 ( 
.A(n_2034),
.B(n_1719),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1900),
.Y(n_2168)
);

INVx3_ASAP7_75t_L g2169 ( 
.A(n_1845),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1891),
.Y(n_2170)
);

O2A1O1Ixp33_ASAP7_75t_L g2171 ( 
.A1(n_1930),
.A2(n_1831),
.B(n_756),
.C(n_764),
.Y(n_2171)
);

AOI21xp5_ASAP7_75t_L g2172 ( 
.A1(n_1997),
.A2(n_1512),
.B(n_1569),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2018),
.B(n_1511),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_SL g2174 ( 
.A(n_1924),
.B(n_1605),
.Y(n_2174)
);

NOR2xp33_ASAP7_75t_L g2175 ( 
.A(n_1894),
.B(n_1397),
.Y(n_2175)
);

AOI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_2003),
.A2(n_1512),
.B(n_1556),
.Y(n_2176)
);

AOI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_2003),
.A2(n_1566),
.B(n_1561),
.Y(n_2177)
);

AND2x2_ASAP7_75t_SL g2178 ( 
.A(n_1874),
.B(n_1511),
.Y(n_2178)
);

AOI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_1923),
.A2(n_1566),
.B(n_1561),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_1970),
.B(n_1489),
.Y(n_2180)
);

AOI21xp5_ASAP7_75t_L g2181 ( 
.A1(n_1944),
.A2(n_1482),
.B(n_1481),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2029),
.B(n_1553),
.Y(n_2182)
);

AOI21xp5_ASAP7_75t_L g2183 ( 
.A1(n_1944),
.A2(n_1482),
.B(n_1481),
.Y(n_2183)
);

OAI21xp5_ASAP7_75t_L g2184 ( 
.A1(n_2024),
.A2(n_1717),
.B(n_1711),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1895),
.B(n_1559),
.Y(n_2185)
);

AOI21xp5_ASAP7_75t_L g2186 ( 
.A1(n_1968),
.A2(n_1636),
.B(n_1633),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_L g2187 ( 
.A(n_1896),
.B(n_1489),
.Y(n_2187)
);

INVx3_ASAP7_75t_L g2188 ( 
.A(n_1947),
.Y(n_2188)
);

INVx3_ASAP7_75t_L g2189 ( 
.A(n_1947),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_1970),
.B(n_1579),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1898),
.B(n_1559),
.Y(n_2191)
);

AOI21xp5_ASAP7_75t_L g2192 ( 
.A1(n_1968),
.A2(n_1636),
.B(n_1633),
.Y(n_2192)
);

HB1xp67_ASAP7_75t_L g2193 ( 
.A(n_2022),
.Y(n_2193)
);

AOI21x1_ASAP7_75t_L g2194 ( 
.A1(n_2010),
.A2(n_1534),
.B(n_1531),
.Y(n_2194)
);

OAI22xp5_ASAP7_75t_L g2195 ( 
.A1(n_1924),
.A2(n_1633),
.B1(n_1654),
.B2(n_1631),
.Y(n_2195)
);

OR2x2_ASAP7_75t_L g2196 ( 
.A(n_1901),
.B(n_1579),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1903),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_L g2198 ( 
.A(n_1906),
.B(n_1756),
.Y(n_2198)
);

AOI21xp5_ASAP7_75t_L g2199 ( 
.A1(n_1983),
.A2(n_1633),
.B(n_1631),
.Y(n_2199)
);

OAI21xp5_ASAP7_75t_L g2200 ( 
.A1(n_2028),
.A2(n_1450),
.B(n_1426),
.Y(n_2200)
);

AOI21xp33_ASAP7_75t_L g2201 ( 
.A1(n_1838),
.A2(n_1501),
.B(n_1463),
.Y(n_2201)
);

O2A1O1Ixp5_ASAP7_75t_L g2202 ( 
.A1(n_1983),
.A2(n_1756),
.B(n_1572),
.C(n_1506),
.Y(n_2202)
);

INVx3_ASAP7_75t_L g2203 ( 
.A(n_1976),
.Y(n_2203)
);

OAI22xp5_ASAP7_75t_L g2204 ( 
.A1(n_1907),
.A2(n_1674),
.B1(n_1677),
.B2(n_1665),
.Y(n_2204)
);

NAND3xp33_ASAP7_75t_L g2205 ( 
.A(n_1897),
.B(n_635),
.C(n_633),
.Y(n_2205)
);

INVxp67_ASAP7_75t_SL g2206 ( 
.A(n_1978),
.Y(n_2206)
);

AOI21xp5_ASAP7_75t_L g2207 ( 
.A1(n_2028),
.A2(n_1654),
.B(n_1631),
.Y(n_2207)
);

AOI21xp5_ASAP7_75t_L g2208 ( 
.A1(n_2031),
.A2(n_1654),
.B(n_1631),
.Y(n_2208)
);

AOI21xp5_ASAP7_75t_L g2209 ( 
.A1(n_2032),
.A2(n_1657),
.B(n_1654),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1908),
.Y(n_2210)
);

AOI21xp5_ASAP7_75t_L g2211 ( 
.A1(n_2035),
.A2(n_1660),
.B(n_1657),
.Y(n_2211)
);

AOI21xp5_ASAP7_75t_L g2212 ( 
.A1(n_1978),
.A2(n_1660),
.B(n_1657),
.Y(n_2212)
);

AO22x1_ASAP7_75t_L g2213 ( 
.A1(n_1979),
.A2(n_638),
.B1(n_639),
.B2(n_637),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_1909),
.Y(n_2214)
);

AOI21xp5_ASAP7_75t_L g2215 ( 
.A1(n_1995),
.A2(n_1660),
.B(n_1657),
.Y(n_2215)
);

A2O1A1Ixp33_ASAP7_75t_L g2216 ( 
.A1(n_1934),
.A2(n_1454),
.B(n_1441),
.C(n_1563),
.Y(n_2216)
);

AOI21xp5_ASAP7_75t_L g2217 ( 
.A1(n_1995),
.A2(n_1665),
.B(n_1660),
.Y(n_2217)
);

AOI21xp5_ASAP7_75t_L g2218 ( 
.A1(n_1973),
.A2(n_1674),
.B(n_1665),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1911),
.B(n_1563),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_1834),
.B(n_1567),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_1835),
.B(n_1567),
.Y(n_2221)
);

AND2x6_ASAP7_75t_L g2222 ( 
.A(n_1973),
.B(n_1665),
.Y(n_2222)
);

NOR2x1_ASAP7_75t_L g2223 ( 
.A(n_1888),
.B(n_1674),
.Y(n_2223)
);

AOI21xp5_ASAP7_75t_L g2224 ( 
.A1(n_1976),
.A2(n_1677),
.B(n_1674),
.Y(n_2224)
);

HB1xp67_ASAP7_75t_L g2225 ( 
.A(n_2015),
.Y(n_2225)
);

AOI21xp5_ASAP7_75t_L g2226 ( 
.A1(n_2015),
.A2(n_1678),
.B(n_1677),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_1914),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1840),
.B(n_1573),
.Y(n_2228)
);

NOR2xp33_ASAP7_75t_SL g2229 ( 
.A(n_1931),
.B(n_1677),
.Y(n_2229)
);

OAI21xp5_ASAP7_75t_L g2230 ( 
.A1(n_1934),
.A2(n_1853),
.B(n_1851),
.Y(n_2230)
);

A2O1A1Ixp33_ASAP7_75t_L g2231 ( 
.A1(n_1841),
.A2(n_1575),
.B(n_1580),
.C(n_1573),
.Y(n_2231)
);

AOI21xp5_ASAP7_75t_L g2232 ( 
.A1(n_1915),
.A2(n_1697),
.B(n_1678),
.Y(n_2232)
);

AOI21xp5_ASAP7_75t_L g2233 ( 
.A1(n_1956),
.A2(n_1697),
.B(n_1678),
.Y(n_2233)
);

OA22x2_ASAP7_75t_L g2234 ( 
.A1(n_1979),
.A2(n_641),
.B1(n_642),
.B2(n_640),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1842),
.B(n_1575),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1849),
.B(n_1580),
.Y(n_2236)
);

AOI21xp5_ASAP7_75t_L g2237 ( 
.A1(n_1941),
.A2(n_1697),
.B(n_1678),
.Y(n_2237)
);

OAI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_1838),
.A2(n_1741),
.B1(n_1719),
.B2(n_1697),
.Y(n_2238)
);

HB1xp67_ASAP7_75t_L g2239 ( 
.A(n_1935),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1926),
.B(n_1475),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_1926),
.B(n_1478),
.Y(n_2241)
);

NOR2xp33_ASAP7_75t_L g2242 ( 
.A(n_1936),
.B(n_1719),
.Y(n_2242)
);

AOI21xp5_ASAP7_75t_L g2243 ( 
.A1(n_1941),
.A2(n_1741),
.B(n_1560),
.Y(n_2243)
);

AOI21xp5_ASAP7_75t_L g2244 ( 
.A1(n_1945),
.A2(n_1741),
.B(n_1386),
.Y(n_2244)
);

NOR2xp33_ASAP7_75t_L g2245 ( 
.A(n_1938),
.B(n_1583),
.Y(n_2245)
);

HB1xp67_ASAP7_75t_L g2246 ( 
.A(n_1935),
.Y(n_2246)
);

NAND2x2_ASAP7_75t_L g2247 ( 
.A(n_1848),
.B(n_740),
.Y(n_2247)
);

AOI21xp5_ASAP7_75t_L g2248 ( 
.A1(n_1945),
.A2(n_1680),
.B(n_1423),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_1929),
.B(n_1583),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_1929),
.B(n_1989),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_1919),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_1989),
.B(n_1458),
.Y(n_2252)
);

AOI22x1_ASAP7_75t_L g2253 ( 
.A1(n_1961),
.A2(n_1464),
.B1(n_1465),
.B2(n_1462),
.Y(n_2253)
);

OAI22xp5_ASAP7_75t_L g2254 ( 
.A1(n_1879),
.A2(n_1423),
.B1(n_1439),
.B2(n_1357),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1940),
.Y(n_2255)
);

NAND2x1p5_ASAP7_75t_L g2256 ( 
.A(n_1888),
.B(n_1496),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_1984),
.Y(n_2257)
);

OAI21xp5_ASAP7_75t_L g2258 ( 
.A1(n_1942),
.A2(n_1464),
.B(n_1462),
.Y(n_2258)
);

A2O1A1Ixp33_ASAP7_75t_L g2259 ( 
.A1(n_1948),
.A2(n_1466),
.B(n_1468),
.C(n_1465),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1959),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_L g2261 ( 
.A(n_1966),
.B(n_1466),
.Y(n_2261)
);

INVx3_ASAP7_75t_L g2262 ( 
.A(n_1939),
.Y(n_2262)
);

AOI21xp5_ASAP7_75t_L g2263 ( 
.A1(n_1961),
.A2(n_1471),
.B(n_1423),
.Y(n_2263)
);

BUFx2_ASAP7_75t_SL g2264 ( 
.A(n_1921),
.Y(n_2264)
);

INVx2_ASAP7_75t_SL g2265 ( 
.A(n_2026),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1977),
.Y(n_2266)
);

AOI21xp5_ASAP7_75t_L g2267 ( 
.A1(n_1969),
.A2(n_1439),
.B(n_1357),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1986),
.Y(n_2268)
);

OAI21xp5_ASAP7_75t_L g2269 ( 
.A1(n_1988),
.A2(n_1992),
.B(n_1991),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_1972),
.B(n_1468),
.Y(n_2270)
);

OAI21xp33_ASAP7_75t_L g2271 ( 
.A1(n_2001),
.A2(n_645),
.B(n_643),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_1850),
.B(n_740),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1932),
.Y(n_2273)
);

NOR2xp33_ASAP7_75t_L g2274 ( 
.A(n_1933),
.B(n_1469),
.Y(n_2274)
);

INVxp67_ASAP7_75t_L g2275 ( 
.A(n_1985),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1972),
.B(n_1469),
.Y(n_2276)
);

AOI21xp5_ASAP7_75t_L g2277 ( 
.A1(n_2051),
.A2(n_1969),
.B(n_1889),
.Y(n_2277)
);

AOI22xp33_ASAP7_75t_L g2278 ( 
.A1(n_2052),
.A2(n_1850),
.B1(n_1994),
.B2(n_1854),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2096),
.Y(n_2279)
);

AOI21xp5_ASAP7_75t_L g2280 ( 
.A1(n_2069),
.A2(n_1889),
.B(n_1879),
.Y(n_2280)
);

O2A1O1Ixp33_ASAP7_75t_SL g2281 ( 
.A1(n_2104),
.A2(n_1939),
.B(n_1952),
.C(n_1943),
.Y(n_2281)
);

O2A1O1Ixp33_ASAP7_75t_L g2282 ( 
.A1(n_2054),
.A2(n_764),
.B(n_765),
.C(n_761),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_L g2283 ( 
.A(n_2052),
.B(n_1990),
.Y(n_2283)
);

INVx1_ASAP7_75t_SL g2284 ( 
.A(n_2120),
.Y(n_2284)
);

NOR4xp25_ASAP7_75t_SL g2285 ( 
.A(n_2148),
.B(n_2019),
.C(n_1974),
.D(n_2023),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2046),
.B(n_1994),
.Y(n_2286)
);

OA22x2_ASAP7_75t_L g2287 ( 
.A1(n_2106),
.A2(n_2085),
.B1(n_2059),
.B2(n_2272),
.Y(n_2287)
);

AOI21xp5_ASAP7_75t_L g2288 ( 
.A1(n_2057),
.A2(n_1889),
.B(n_2019),
.Y(n_2288)
);

NOR2xp33_ASAP7_75t_L g2289 ( 
.A(n_2058),
.B(n_2000),
.Y(n_2289)
);

AOI21xp5_ASAP7_75t_L g2290 ( 
.A1(n_2118),
.A2(n_1975),
.B(n_2023),
.Y(n_2290)
);

NOR2xp33_ASAP7_75t_L g2291 ( 
.A(n_2104),
.B(n_1953),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2251),
.Y(n_2292)
);

OAI22xp5_ASAP7_75t_L g2293 ( 
.A1(n_2068),
.A2(n_1975),
.B1(n_1985),
.B2(n_1974),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_2056),
.B(n_1963),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2273),
.Y(n_2295)
);

INVx4_ASAP7_75t_L g2296 ( 
.A(n_2149),
.Y(n_2296)
);

AOI221xp5_ASAP7_75t_L g2297 ( 
.A1(n_2271),
.A2(n_2001),
.B1(n_2008),
.B2(n_2005),
.C(n_1854),
.Y(n_2297)
);

AOI21xp5_ASAP7_75t_L g2298 ( 
.A1(n_2108),
.A2(n_2030),
.B(n_1439),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2068),
.B(n_1858),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_L g2300 ( 
.A(n_2073),
.B(n_1957),
.Y(n_2300)
);

AOI21xp5_ASAP7_75t_L g2301 ( 
.A1(n_2125),
.A2(n_2030),
.B(n_1460),
.Y(n_2301)
);

O2A1O1Ixp33_ASAP7_75t_L g2302 ( 
.A1(n_2088),
.A2(n_765),
.B(n_785),
.C(n_761),
.Y(n_2302)
);

NAND3xp33_ASAP7_75t_SL g2303 ( 
.A(n_2065),
.B(n_648),
.C(n_647),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_SL g2304 ( 
.A(n_2070),
.B(n_1963),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2117),
.B(n_1858),
.Y(n_2305)
);

AOI21xp5_ASAP7_75t_L g2306 ( 
.A1(n_2100),
.A2(n_1460),
.B(n_1357),
.Y(n_2306)
);

AOI21xp5_ASAP7_75t_L g2307 ( 
.A1(n_2097),
.A2(n_1471),
.B(n_1460),
.Y(n_2307)
);

BUFx2_ASAP7_75t_R g2308 ( 
.A(n_2045),
.Y(n_2308)
);

NOR2xp33_ASAP7_75t_L g2309 ( 
.A(n_2072),
.B(n_1962),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2067),
.B(n_2005),
.Y(n_2310)
);

AO22x1_ASAP7_75t_L g2311 ( 
.A1(n_2161),
.A2(n_653),
.B1(n_659),
.B2(n_652),
.Y(n_2311)
);

BUFx3_ASAP7_75t_L g2312 ( 
.A(n_2149),
.Y(n_2312)
);

HB1xp67_ASAP7_75t_L g2313 ( 
.A(n_2080),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2121),
.Y(n_2314)
);

BUFx2_ASAP7_75t_L g2315 ( 
.A(n_2067),
.Y(n_2315)
);

AOI21xp5_ASAP7_75t_L g2316 ( 
.A1(n_2060),
.A2(n_1496),
.B(n_1471),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_2065),
.B(n_1987),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_SL g2318 ( 
.A(n_2230),
.B(n_1984),
.Y(n_2318)
);

OR2x2_ASAP7_75t_L g2319 ( 
.A(n_2111),
.B(n_939),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_L g2320 ( 
.A(n_2077),
.B(n_1472),
.Y(n_2320)
);

OAI21x1_ASAP7_75t_L g2321 ( 
.A1(n_2107),
.A2(n_1572),
.B(n_1509),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2137),
.Y(n_2322)
);

AOI21xp5_ASAP7_75t_L g2323 ( 
.A1(n_2061),
.A2(n_1509),
.B(n_1496),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_2079),
.B(n_1472),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2077),
.B(n_2008),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2227),
.Y(n_2326)
);

AOI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_2064),
.A2(n_1517),
.B(n_1509),
.Y(n_2327)
);

NOR2xp33_ASAP7_75t_L g2328 ( 
.A(n_2049),
.B(n_1473),
.Y(n_2328)
);

INVx4_ASAP7_75t_L g2329 ( 
.A(n_2149),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2151),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2153),
.B(n_1860),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2170),
.Y(n_2332)
);

NOR2x1_ASAP7_75t_R g2333 ( 
.A(n_2047),
.B(n_661),
.Y(n_2333)
);

AOI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_2076),
.A2(n_2081),
.B(n_2078),
.Y(n_2334)
);

BUFx2_ASAP7_75t_L g2335 ( 
.A(n_2196),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2093),
.B(n_1860),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_L g2337 ( 
.A(n_2050),
.B(n_1473),
.Y(n_2337)
);

OR2x2_ASAP7_75t_L g2338 ( 
.A(n_2110),
.B(n_939),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2133),
.B(n_2134),
.Y(n_2339)
);

INVx3_ASAP7_75t_L g2340 ( 
.A(n_2139),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2197),
.Y(n_2341)
);

AOI21xp5_ASAP7_75t_L g2342 ( 
.A1(n_2083),
.A2(n_1517),
.B(n_1474),
.Y(n_2342)
);

O2A1O1Ixp5_ASAP7_75t_L g2343 ( 
.A1(n_2194),
.A2(n_1474),
.B(n_1517),
.C(n_1382),
.Y(n_2343)
);

OAI22xp5_ASAP7_75t_L g2344 ( 
.A1(n_2075),
.A2(n_1875),
.B1(n_1885),
.B2(n_1866),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_L g2345 ( 
.A(n_2050),
.B(n_1380),
.Y(n_2345)
);

A2O1A1Ixp33_ASAP7_75t_L g2346 ( 
.A1(n_2123),
.A2(n_790),
.B(n_795),
.C(n_785),
.Y(n_2346)
);

NOR2xp33_ASAP7_75t_L g2347 ( 
.A(n_2229),
.B(n_1382),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2135),
.B(n_1866),
.Y(n_2348)
);

INVx5_ASAP7_75t_L g2349 ( 
.A(n_2160),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2144),
.B(n_1875),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_2187),
.B(n_740),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2158),
.B(n_1885),
.Y(n_2352)
);

AOI21x1_ASAP7_75t_L g2353 ( 
.A1(n_2066),
.A2(n_1902),
.B(n_1899),
.Y(n_2353)
);

AOI21xp5_ASAP7_75t_L g2354 ( 
.A1(n_2084),
.A2(n_1389),
.B(n_1388),
.Y(n_2354)
);

AOI21x1_ASAP7_75t_L g2355 ( 
.A1(n_2098),
.A2(n_2176),
.B(n_2248),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2129),
.B(n_1899),
.Y(n_2356)
);

AND2x4_ASAP7_75t_L g2357 ( 
.A(n_2074),
.B(n_1388),
.Y(n_2357)
);

AOI21xp5_ASAP7_75t_L g2358 ( 
.A1(n_2087),
.A2(n_1394),
.B(n_1389),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2210),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_2187),
.B(n_759),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2048),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2129),
.B(n_1902),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2255),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2260),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2055),
.Y(n_2365)
);

AOI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2092),
.A2(n_1400),
.B(n_1394),
.Y(n_2366)
);

CKINVDCx20_ASAP7_75t_R g2367 ( 
.A(n_2161),
.Y(n_2367)
);

CKINVDCx11_ASAP7_75t_R g2368 ( 
.A(n_2157),
.Y(n_2368)
);

AOI21xp5_ASAP7_75t_L g2369 ( 
.A1(n_2215),
.A2(n_2217),
.B(n_2086),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2099),
.B(n_664),
.Y(n_2370)
);

AOI21xp5_ASAP7_75t_L g2371 ( 
.A1(n_2218),
.A2(n_1406),
.B(n_1400),
.Y(n_2371)
);

INVx3_ASAP7_75t_L g2372 ( 
.A(n_2139),
.Y(n_2372)
);

HB1xp67_ASAP7_75t_L g2373 ( 
.A(n_2094),
.Y(n_2373)
);

NOR3xp33_ASAP7_75t_SL g2374 ( 
.A(n_2113),
.B(n_670),
.C(n_667),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2102),
.B(n_674),
.Y(n_2375)
);

INVx4_ASAP7_75t_L g2376 ( 
.A(n_2160),
.Y(n_2376)
);

O2A1O1Ixp33_ASAP7_75t_L g2377 ( 
.A1(n_2113),
.A2(n_2132),
.B(n_2167),
.C(n_2095),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_SL g2378 ( 
.A(n_2265),
.B(n_1526),
.Y(n_2378)
);

NOR2xp33_ASAP7_75t_L g2379 ( 
.A(n_2114),
.B(n_2122),
.Y(n_2379)
);

NOR2xp33_ASAP7_75t_L g2380 ( 
.A(n_2124),
.B(n_1406),
.Y(n_2380)
);

AND2x4_ASAP7_75t_L g2381 ( 
.A(n_2074),
.B(n_1407),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2266),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_2175),
.B(n_759),
.Y(n_2383)
);

NOR2xp33_ASAP7_75t_SL g2384 ( 
.A(n_2075),
.B(n_1526),
.Y(n_2384)
);

OR2x6_ASAP7_75t_L g2385 ( 
.A(n_2264),
.B(n_1407),
.Y(n_2385)
);

AOI21xp5_ASAP7_75t_L g2386 ( 
.A1(n_2098),
.A2(n_1415),
.B(n_1408),
.Y(n_2386)
);

BUFx6f_ASAP7_75t_L g2387 ( 
.A(n_2257),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2062),
.Y(n_2388)
);

AOI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_2244),
.A2(n_1415),
.B(n_1408),
.Y(n_2389)
);

AOI221xp5_ASAP7_75t_L g2390 ( 
.A1(n_2250),
.A2(n_682),
.B1(n_683),
.B2(n_678),
.C(n_676),
.Y(n_2390)
);

NAND3xp33_ASAP7_75t_L g2391 ( 
.A(n_2205),
.B(n_688),
.C(n_686),
.Y(n_2391)
);

NOR3xp33_ASAP7_75t_L g2392 ( 
.A(n_2213),
.B(n_795),
.C(n_790),
.Y(n_2392)
);

AOI21xp5_ASAP7_75t_L g2393 ( 
.A1(n_2155),
.A2(n_1427),
.B(n_1420),
.Y(n_2393)
);

CKINVDCx5p33_ASAP7_75t_R g2394 ( 
.A(n_2159),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2115),
.Y(n_2395)
);

A2O1A1Ixp33_ASAP7_75t_L g2396 ( 
.A1(n_2123),
.A2(n_800),
.B(n_803),
.C(n_797),
.Y(n_2396)
);

NOR2xp33_ASAP7_75t_L g2397 ( 
.A(n_2112),
.B(n_1420),
.Y(n_2397)
);

NOR2xp33_ASAP7_75t_L g2398 ( 
.A(n_2173),
.B(n_1427),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2109),
.B(n_692),
.Y(n_2399)
);

INVx1_ASAP7_75t_SL g2400 ( 
.A(n_2160),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2119),
.B(n_693),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2090),
.B(n_694),
.Y(n_2402)
);

AOI21xp5_ASAP7_75t_L g2403 ( 
.A1(n_2126),
.A2(n_1432),
.B(n_1431),
.Y(n_2403)
);

AOI22xp33_ASAP7_75t_L g2404 ( 
.A1(n_2234),
.A2(n_768),
.B1(n_772),
.B2(n_759),
.Y(n_2404)
);

OAI22xp5_ASAP7_75t_L g2405 ( 
.A1(n_2175),
.A2(n_699),
.B1(n_702),
.B2(n_695),
.Y(n_2405)
);

NOR2xp33_ASAP7_75t_L g2406 ( 
.A(n_2140),
.B(n_1431),
.Y(n_2406)
);

OAI21x1_ASAP7_75t_L g2407 ( 
.A1(n_2177),
.A2(n_1432),
.B(n_1078),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2140),
.B(n_705),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2268),
.Y(n_2409)
);

BUFx3_ASAP7_75t_L g2410 ( 
.A(n_2091),
.Y(n_2410)
);

HB1xp67_ASAP7_75t_L g2411 ( 
.A(n_2110),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2147),
.Y(n_2412)
);

AND2x4_ASAP7_75t_L g2413 ( 
.A(n_2091),
.B(n_1526),
.Y(n_2413)
);

BUFx6f_ASAP7_75t_L g2414 ( 
.A(n_2257),
.Y(n_2414)
);

O2A1O1Ixp33_ASAP7_75t_L g2415 ( 
.A1(n_2063),
.A2(n_800),
.B(n_803),
.C(n_797),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2101),
.B(n_706),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2101),
.B(n_707),
.Y(n_2417)
);

AOI21xp5_ASAP7_75t_L g2418 ( 
.A1(n_2163),
.A2(n_1200),
.B(n_1123),
.Y(n_2418)
);

INVx1_ASAP7_75t_SL g2419 ( 
.A(n_2193),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_SL g2420 ( 
.A(n_2131),
.B(n_759),
.Y(n_2420)
);

NOR2xp33_ASAP7_75t_L g2421 ( 
.A(n_2193),
.B(n_708),
.Y(n_2421)
);

AOI21xp5_ASAP7_75t_L g2422 ( 
.A1(n_2184),
.A2(n_1200),
.B(n_1535),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_SL g2423 ( 
.A(n_2131),
.B(n_768),
.Y(n_2423)
);

INVx2_ASAP7_75t_SL g2424 ( 
.A(n_2257),
.Y(n_2424)
);

AOI21xp5_ASAP7_75t_L g2425 ( 
.A1(n_2103),
.A2(n_1189),
.B(n_1181),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2198),
.B(n_709),
.Y(n_2426)
);

BUFx6f_ASAP7_75t_L g2427 ( 
.A(n_2257),
.Y(n_2427)
);

INVx3_ASAP7_75t_L g2428 ( 
.A(n_2262),
.Y(n_2428)
);

A2O1A1Ixp33_ASAP7_75t_L g2429 ( 
.A1(n_2053),
.A2(n_815),
.B(n_820),
.C(n_807),
.Y(n_2429)
);

OAI22xp5_ASAP7_75t_L g2430 ( 
.A1(n_2136),
.A2(n_716),
.B1(n_717),
.B2(n_715),
.Y(n_2430)
);

BUFx10_ASAP7_75t_L g2431 ( 
.A(n_2136),
.Y(n_2431)
);

NAND3xp33_ASAP7_75t_SL g2432 ( 
.A(n_2138),
.B(n_722),
.C(n_718),
.Y(n_2432)
);

AOI21xp5_ASAP7_75t_L g2433 ( 
.A1(n_2103),
.A2(n_1189),
.B(n_1181),
.Y(n_2433)
);

A2O1A1Ixp33_ASAP7_75t_L g2434 ( 
.A1(n_2198),
.A2(n_815),
.B(n_820),
.C(n_807),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2152),
.Y(n_2435)
);

INVx4_ASAP7_75t_L g2436 ( 
.A(n_2082),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_SL g2437 ( 
.A(n_2138),
.B(n_768),
.Y(n_2437)
);

OAI21xp33_ASAP7_75t_L g2438 ( 
.A1(n_2234),
.A2(n_730),
.B(n_728),
.Y(n_2438)
);

BUFx6f_ASAP7_75t_L g2439 ( 
.A(n_2262),
.Y(n_2439)
);

OR2x2_ASAP7_75t_L g2440 ( 
.A(n_2168),
.B(n_942),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2182),
.B(n_731),
.Y(n_2441)
);

NOR2xp33_ASAP7_75t_L g2442 ( 
.A(n_2178),
.B(n_732),
.Y(n_2442)
);

AOI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2128),
.A2(n_1189),
.B(n_1181),
.Y(n_2443)
);

NOR2xp33_ASAP7_75t_L g2444 ( 
.A(n_2178),
.B(n_735),
.Y(n_2444)
);

AOI21xp5_ASAP7_75t_L g2445 ( 
.A1(n_2130),
.A2(n_1189),
.B(n_1181),
.Y(n_2445)
);

A2O1A1Ixp33_ASAP7_75t_L g2446 ( 
.A1(n_2154),
.A2(n_831),
.B(n_833),
.C(n_822),
.Y(n_2446)
);

AOI21xp5_ASAP7_75t_L g2447 ( 
.A1(n_2206),
.A2(n_1206),
.B(n_1189),
.Y(n_2447)
);

BUFx4f_ASAP7_75t_L g2448 ( 
.A(n_2180),
.Y(n_2448)
);

AOI21xp5_ASAP7_75t_L g2449 ( 
.A1(n_2206),
.A2(n_1220),
.B(n_1206),
.Y(n_2449)
);

AOI21xp5_ASAP7_75t_L g2450 ( 
.A1(n_2200),
.A2(n_1220),
.B(n_1206),
.Y(n_2450)
);

INVxp67_ASAP7_75t_L g2451 ( 
.A(n_2239),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2214),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2239),
.Y(n_2453)
);

NAND3xp33_ASAP7_75t_SL g2454 ( 
.A(n_2154),
.B(n_739),
.C(n_736),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2162),
.B(n_743),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2246),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2185),
.B(n_744),
.Y(n_2457)
);

AND2x2_ASAP7_75t_L g2458 ( 
.A(n_2190),
.B(n_2246),
.Y(n_2458)
);

BUFx2_ASAP7_75t_L g2459 ( 
.A(n_2225),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2191),
.B(n_745),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2219),
.B(n_750),
.Y(n_2461)
);

A2O1A1Ixp33_ASAP7_75t_L g2462 ( 
.A1(n_2156),
.A2(n_831),
.B(n_834),
.C(n_822),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_SL g2463 ( 
.A(n_2156),
.B(n_768),
.Y(n_2463)
);

AOI22xp33_ASAP7_75t_L g2464 ( 
.A1(n_2146),
.A2(n_772),
.B1(n_754),
.B2(n_755),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_SL g2465 ( 
.A(n_2269),
.B(n_2220),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2221),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_SL g2467 ( 
.A(n_2228),
.B(n_772),
.Y(n_2467)
);

INVx2_ASAP7_75t_SL g2468 ( 
.A(n_2247),
.Y(n_2468)
);

O2A1O1Ixp33_ASAP7_75t_SL g2469 ( 
.A1(n_2216),
.A2(n_931),
.B(n_932),
.C(n_930),
.Y(n_2469)
);

A2O1A1Ixp33_ASAP7_75t_L g2470 ( 
.A1(n_2142),
.A2(n_757),
.B(n_760),
.C(n_752),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2235),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2236),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2274),
.Y(n_2473)
);

NOR3xp33_ASAP7_75t_SL g2474 ( 
.A(n_2238),
.B(n_763),
.C(n_762),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2274),
.Y(n_2475)
);

O2A1O1Ixp33_ASAP7_75t_L g2476 ( 
.A1(n_2201),
.A2(n_945),
.B(n_951),
.C(n_942),
.Y(n_2476)
);

OR2x2_ASAP7_75t_L g2477 ( 
.A(n_2240),
.B(n_945),
.Y(n_2477)
);

BUFx6f_ASAP7_75t_L g2478 ( 
.A(n_2174),
.Y(n_2478)
);

A2O1A1Ixp33_ASAP7_75t_L g2479 ( 
.A1(n_2171),
.A2(n_769),
.B(n_770),
.C(n_767),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2261),
.B(n_771),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2245),
.Y(n_2481)
);

INVx4_ASAP7_75t_L g2482 ( 
.A(n_2082),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_SL g2483 ( 
.A(n_2146),
.B(n_954),
.Y(n_2483)
);

INVx1_ASAP7_75t_SL g2484 ( 
.A(n_2225),
.Y(n_2484)
);

A2O1A1Ixp33_ASAP7_75t_L g2485 ( 
.A1(n_2237),
.A2(n_773),
.B(n_775),
.C(n_774),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2261),
.Y(n_2486)
);

OAI21x1_ASAP7_75t_L g2487 ( 
.A1(n_2071),
.A2(n_1078),
.B(n_1076),
.Y(n_2487)
);

BUFx2_ASAP7_75t_L g2488 ( 
.A(n_2223),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2245),
.Y(n_2489)
);

NOR3xp33_ASAP7_75t_SL g2490 ( 
.A(n_2254),
.B(n_777),
.C(n_776),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2256),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2256),
.Y(n_2492)
);

OAI22xp5_ASAP7_75t_L g2493 ( 
.A1(n_2116),
.A2(n_778),
.B1(n_784),
.B2(n_780),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2105),
.Y(n_2494)
);

BUFx3_ASAP7_75t_L g2495 ( 
.A(n_2169),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2249),
.Y(n_2496)
);

INVx2_ASAP7_75t_SL g2497 ( 
.A(n_2247),
.Y(n_2497)
);

O2A1O1Ixp33_ASAP7_75t_L g2498 ( 
.A1(n_2241),
.A2(n_2276),
.B(n_2270),
.C(n_2252),
.Y(n_2498)
);

NAND2x1p5_ASAP7_75t_L g2499 ( 
.A(n_2169),
.B(n_2188),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2242),
.Y(n_2500)
);

HB1xp67_ASAP7_75t_L g2501 ( 
.A(n_2275),
.Y(n_2501)
);

AOI21xp5_ASAP7_75t_L g2502 ( 
.A1(n_2141),
.A2(n_1220),
.B(n_1206),
.Y(n_2502)
);

AOI21xp5_ASAP7_75t_L g2503 ( 
.A1(n_2243),
.A2(n_1220),
.B(n_1206),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_SL g2504 ( 
.A(n_2242),
.B(n_772),
.Y(n_2504)
);

O2A1O1Ixp5_ASAP7_75t_L g2505 ( 
.A1(n_2127),
.A2(n_952),
.B(n_955),
.C(n_951),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2231),
.Y(n_2506)
);

AOI21xp5_ASAP7_75t_L g2507 ( 
.A1(n_2179),
.A2(n_1226),
.B(n_1220),
.Y(n_2507)
);

A2O1A1Ixp33_ASAP7_75t_L g2508 ( 
.A1(n_2164),
.A2(n_787),
.B(n_788),
.C(n_786),
.Y(n_2508)
);

OR2x6_ASAP7_75t_L g2509 ( 
.A(n_2188),
.B(n_1324),
.Y(n_2509)
);

AOI21xp5_ASAP7_75t_L g2510 ( 
.A1(n_2186),
.A2(n_1227),
.B(n_1226),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2233),
.B(n_789),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_SL g2512 ( 
.A(n_2166),
.B(n_791),
.Y(n_2512)
);

BUFx4f_ASAP7_75t_SL g2513 ( 
.A(n_2189),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2192),
.B(n_2189),
.Y(n_2514)
);

NAND2xp33_ASAP7_75t_SL g2515 ( 
.A(n_2203),
.B(n_792),
.Y(n_2515)
);

AOI21xp5_ASAP7_75t_L g2516 ( 
.A1(n_2224),
.A2(n_1227),
.B(n_1226),
.Y(n_2516)
);

BUFx6f_ASAP7_75t_L g2517 ( 
.A(n_2222),
.Y(n_2517)
);

HB1xp67_ASAP7_75t_L g2518 ( 
.A(n_2275),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2258),
.Y(n_2519)
);

NAND3xp33_ASAP7_75t_L g2520 ( 
.A(n_2165),
.B(n_799),
.C(n_793),
.Y(n_2520)
);

OAI22x1_ASAP7_75t_L g2521 ( 
.A1(n_2253),
.A2(n_805),
.B1(n_808),
.B2(n_804),
.Y(n_2521)
);

INVx8_ASAP7_75t_L g2522 ( 
.A(n_2203),
.Y(n_2522)
);

AOI21xp5_ASAP7_75t_L g2523 ( 
.A1(n_2212),
.A2(n_1227),
.B(n_1226),
.Y(n_2523)
);

AO22x1_ASAP7_75t_L g2524 ( 
.A1(n_2222),
.A2(n_817),
.B1(n_821),
.B2(n_811),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_2207),
.B(n_824),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_SL g2526 ( 
.A(n_2208),
.B(n_825),
.Y(n_2526)
);

INVx5_ASAP7_75t_L g2527 ( 
.A(n_2222),
.Y(n_2527)
);

O2A1O1Ixp33_ASAP7_75t_L g2528 ( 
.A1(n_2164),
.A2(n_955),
.B(n_956),
.C(n_952),
.Y(n_2528)
);

AOI21xp5_ASAP7_75t_L g2529 ( 
.A1(n_2181),
.A2(n_2183),
.B(n_2199),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2259),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_SL g2531 ( 
.A(n_2209),
.B(n_828),
.Y(n_2531)
);

AOI21xp5_ASAP7_75t_L g2532 ( 
.A1(n_2143),
.A2(n_1227),
.B(n_1226),
.Y(n_2532)
);

AND2x2_ASAP7_75t_L g2533 ( 
.A(n_2195),
.B(n_956),
.Y(n_2533)
);

CKINVDCx20_ASAP7_75t_R g2534 ( 
.A(n_2204),
.Y(n_2534)
);

AND2x4_ASAP7_75t_L g2535 ( 
.A(n_2226),
.B(n_1526),
.Y(n_2535)
);

NOR2x1_ASAP7_75t_L g2536 ( 
.A(n_2211),
.B(n_957),
.Y(n_2536)
);

AOI22xp5_ASAP7_75t_L g2537 ( 
.A1(n_2222),
.A2(n_1574),
.B1(n_830),
.B2(n_829),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2089),
.Y(n_2538)
);

AOI21xp5_ASAP7_75t_L g2539 ( 
.A1(n_2145),
.A2(n_1227),
.B(n_1313),
.Y(n_2539)
);

OAI21xp5_ASAP7_75t_L g2540 ( 
.A1(n_2202),
.A2(n_1574),
.B(n_958),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2222),
.B(n_1574),
.Y(n_2541)
);

AOI21xp5_ASAP7_75t_L g2542 ( 
.A1(n_2369),
.A2(n_2232),
.B(n_2172),
.Y(n_2542)
);

OAI21x1_ASAP7_75t_L g2543 ( 
.A1(n_2334),
.A2(n_2150),
.B(n_2202),
.Y(n_2543)
);

OAI21x1_ASAP7_75t_L g2544 ( 
.A1(n_2529),
.A2(n_2267),
.B(n_2263),
.Y(n_2544)
);

AOI21xp5_ASAP7_75t_L g2545 ( 
.A1(n_2280),
.A2(n_1078),
.B(n_1076),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2313),
.Y(n_2546)
);

OAI21x1_ASAP7_75t_L g2547 ( 
.A1(n_2487),
.A2(n_1082),
.B(n_1080),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2458),
.B(n_957),
.Y(n_2548)
);

INVx2_ASAP7_75t_SL g2549 ( 
.A(n_2312),
.Y(n_2549)
);

NOR2xp67_ASAP7_75t_L g2550 ( 
.A(n_2391),
.B(n_457),
.Y(n_2550)
);

OAI21xp33_ASAP7_75t_L g2551 ( 
.A1(n_2464),
.A2(n_959),
.B(n_958),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2313),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2379),
.B(n_959),
.Y(n_2553)
);

OA21x2_ASAP7_75t_L g2554 ( 
.A1(n_2343),
.A2(n_967),
.B(n_963),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2330),
.Y(n_2555)
);

INVx5_ASAP7_75t_L g2556 ( 
.A(n_2385),
.Y(n_2556)
);

OAI21x1_ASAP7_75t_L g2557 ( 
.A1(n_2443),
.A2(n_1082),
.B(n_1080),
.Y(n_2557)
);

AOI21xp5_ASAP7_75t_L g2558 ( 
.A1(n_2469),
.A2(n_1082),
.B(n_1080),
.Y(n_2558)
);

AOI21x1_ASAP7_75t_L g2559 ( 
.A1(n_2353),
.A2(n_967),
.B(n_963),
.Y(n_2559)
);

OAI21xp5_ASAP7_75t_L g2560 ( 
.A1(n_2290),
.A2(n_1574),
.B(n_970),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2373),
.Y(n_2561)
);

OAI21x1_ASAP7_75t_L g2562 ( 
.A1(n_2445),
.A2(n_1107),
.B(n_1083),
.Y(n_2562)
);

OAI21xp5_ASAP7_75t_L g2563 ( 
.A1(n_2464),
.A2(n_1574),
.B(n_970),
.Y(n_2563)
);

AOI21xp5_ASAP7_75t_L g2564 ( 
.A1(n_2527),
.A2(n_1107),
.B(n_1083),
.Y(n_2564)
);

NOR2x1_ASAP7_75t_L g2565 ( 
.A(n_2481),
.B(n_968),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2309),
.B(n_968),
.Y(n_2566)
);

AOI21xp5_ASAP7_75t_L g2567 ( 
.A1(n_2527),
.A2(n_2465),
.B(n_2422),
.Y(n_2567)
);

AOI21xp5_ASAP7_75t_L g2568 ( 
.A1(n_2527),
.A2(n_1107),
.B(n_1083),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_SL g2569 ( 
.A(n_2486),
.B(n_976),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2332),
.Y(n_2570)
);

OR2x2_ASAP7_75t_L g2571 ( 
.A(n_2411),
.B(n_976),
.Y(n_2571)
);

OAI22xp5_ASAP7_75t_L g2572 ( 
.A1(n_2278),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2373),
.Y(n_2573)
);

OAI21xp5_ASAP7_75t_L g2574 ( 
.A1(n_2415),
.A2(n_937),
.B(n_934),
.Y(n_2574)
);

AOI31xp67_ASAP7_75t_L g2575 ( 
.A1(n_2287),
.A2(n_1324),
.A3(n_938),
.B(n_937),
.Y(n_2575)
);

OAI21x1_ASAP7_75t_L g2576 ( 
.A1(n_2355),
.A2(n_2389),
.B(n_2321),
.Y(n_2576)
);

OAI22xp5_ASAP7_75t_L g2577 ( 
.A1(n_2278),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_2577)
);

OAI21xp5_ASAP7_75t_L g2578 ( 
.A1(n_2302),
.A2(n_938),
.B(n_857),
.Y(n_2578)
);

OR2x2_ASAP7_75t_L g2579 ( 
.A(n_2411),
.B(n_854),
.Y(n_2579)
);

AO31x2_ASAP7_75t_L g2580 ( 
.A1(n_2293),
.A2(n_859),
.A3(n_860),
.B(n_858),
.Y(n_2580)
);

OR2x2_ASAP7_75t_L g2581 ( 
.A(n_2310),
.B(n_858),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2501),
.Y(n_2582)
);

NAND3x1_ASAP7_75t_L g2583 ( 
.A(n_2392),
.B(n_5),
.C(n_6),
.Y(n_2583)
);

OAI21x1_ASAP7_75t_L g2584 ( 
.A1(n_2403),
.A2(n_860),
.B(n_859),
.Y(n_2584)
);

OAI21x1_ASAP7_75t_L g2585 ( 
.A1(n_2407),
.A2(n_866),
.B(n_865),
.Y(n_2585)
);

AO31x2_ASAP7_75t_L g2586 ( 
.A1(n_2277),
.A2(n_866),
.A3(n_869),
.B(n_865),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2466),
.B(n_5),
.Y(n_2587)
);

AOI22xp5_ASAP7_75t_L g2588 ( 
.A1(n_2289),
.A2(n_871),
.B1(n_872),
.B2(n_869),
.Y(n_2588)
);

AOI21xp5_ASAP7_75t_L g2589 ( 
.A1(n_2527),
.A2(n_872),
.B(n_871),
.Y(n_2589)
);

OAI21x1_ASAP7_75t_L g2590 ( 
.A1(n_2306),
.A2(n_876),
.B(n_874),
.Y(n_2590)
);

AO21x2_ASAP7_75t_L g2591 ( 
.A1(n_2288),
.A2(n_876),
.B(n_874),
.Y(n_2591)
);

AOI21xp5_ASAP7_75t_L g2592 ( 
.A1(n_2450),
.A2(n_2339),
.B(n_2540),
.Y(n_2592)
);

INVxp67_ASAP7_75t_SL g2593 ( 
.A(n_2451),
.Y(n_2593)
);

OAI22x1_ASAP7_75t_L g2594 ( 
.A1(n_2442),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_2594)
);

O2A1O1Ixp33_ASAP7_75t_SL g2595 ( 
.A1(n_2351),
.A2(n_2360),
.B(n_2423),
.C(n_2420),
.Y(n_2595)
);

AND2x2_ASAP7_75t_L g2596 ( 
.A(n_2309),
.B(n_459),
.Y(n_2596)
);

AND2x4_ASAP7_75t_L g2597 ( 
.A(n_2459),
.B(n_460),
.Y(n_2597)
);

NOR2xp67_ASAP7_75t_SL g2598 ( 
.A(n_2468),
.B(n_1006),
.Y(n_2598)
);

AOI21xp5_ASAP7_75t_L g2599 ( 
.A1(n_2301),
.A2(n_882),
.B(n_877),
.Y(n_2599)
);

BUFx2_ASAP7_75t_L g2600 ( 
.A(n_2315),
.Y(n_2600)
);

AOI21xp5_ASAP7_75t_L g2601 ( 
.A1(n_2447),
.A2(n_882),
.B(n_877),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2501),
.Y(n_2602)
);

OAI21x1_ASAP7_75t_L g2603 ( 
.A1(n_2502),
.A2(n_1324),
.B(n_1006),
.Y(n_2603)
);

OAI21x1_ASAP7_75t_L g2604 ( 
.A1(n_2503),
.A2(n_1006),
.B(n_1042),
.Y(n_2604)
);

OAI21x1_ASAP7_75t_L g2605 ( 
.A1(n_2532),
.A2(n_2539),
.B(n_2358),
.Y(n_2605)
);

AO31x2_ASAP7_75t_L g2606 ( 
.A1(n_2538),
.A2(n_463),
.A3(n_465),
.B(n_461),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2518),
.Y(n_2607)
);

NOR2x1_ASAP7_75t_L g2608 ( 
.A(n_2432),
.B(n_1006),
.Y(n_2608)
);

NOR2xp33_ASAP7_75t_SL g2609 ( 
.A(n_2308),
.B(n_8),
.Y(n_2609)
);

O2A1O1Ixp33_ASAP7_75t_SL g2610 ( 
.A1(n_2437),
.A2(n_12),
.B(n_9),
.C(n_10),
.Y(n_2610)
);

AOI21xp5_ASAP7_75t_L g2611 ( 
.A1(n_2449),
.A2(n_1006),
.B(n_1002),
.Y(n_2611)
);

INVx2_ASAP7_75t_SL g2612 ( 
.A(n_2349),
.Y(n_2612)
);

INVx5_ASAP7_75t_L g2613 ( 
.A(n_2385),
.Y(n_2613)
);

CKINVDCx6p67_ASAP7_75t_R g2614 ( 
.A(n_2368),
.Y(n_2614)
);

OAI22xp5_ASAP7_75t_L g2615 ( 
.A1(n_2404),
.A2(n_13),
.B1(n_10),
.B2(n_12),
.Y(n_2615)
);

AND2x2_ASAP7_75t_L g2616 ( 
.A(n_2300),
.B(n_466),
.Y(n_2616)
);

AO31x2_ASAP7_75t_L g2617 ( 
.A1(n_2298),
.A2(n_470),
.A3(n_471),
.B(n_469),
.Y(n_2617)
);

AOI211x1_ASAP7_75t_L g2618 ( 
.A1(n_2438),
.A2(n_17),
.B(n_14),
.C(n_15),
.Y(n_2618)
);

O2A1O1Ixp33_ASAP7_75t_SL g2619 ( 
.A1(n_2463),
.A2(n_18),
.B(n_14),
.C(n_17),
.Y(n_2619)
);

INVx4_ASAP7_75t_L g2620 ( 
.A(n_2349),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2518),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2379),
.B(n_18),
.Y(n_2622)
);

AO31x2_ASAP7_75t_L g2623 ( 
.A1(n_2494),
.A2(n_474),
.A3(n_475),
.B(n_473),
.Y(n_2623)
);

AND2x2_ASAP7_75t_L g2624 ( 
.A(n_2300),
.B(n_477),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2326),
.Y(n_2625)
);

BUFx3_ASAP7_75t_L g2626 ( 
.A(n_2335),
.Y(n_2626)
);

BUFx6f_ASAP7_75t_L g2627 ( 
.A(n_2349),
.Y(n_2627)
);

AND2x4_ASAP7_75t_L g2628 ( 
.A(n_2340),
.B(n_479),
.Y(n_2628)
);

OAI21x1_ASAP7_75t_L g2629 ( 
.A1(n_2354),
.A2(n_2366),
.B(n_2342),
.Y(n_2629)
);

AND2x2_ASAP7_75t_L g2630 ( 
.A(n_2299),
.B(n_480),
.Y(n_2630)
);

NOR2x1_ASAP7_75t_SL g2631 ( 
.A(n_2517),
.B(n_1006),
.Y(n_2631)
);

OAI21x1_ASAP7_75t_L g2632 ( 
.A1(n_2316),
.A2(n_1058),
.B(n_1044),
.Y(n_2632)
);

OAI21x1_ASAP7_75t_L g2633 ( 
.A1(n_2323),
.A2(n_1058),
.B(n_1044),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2442),
.B(n_483),
.Y(n_2634)
);

OAI22x1_ASAP7_75t_L g2635 ( 
.A1(n_2444),
.A2(n_2383),
.B1(n_2356),
.B2(n_2362),
.Y(n_2635)
);

INVxp67_ASAP7_75t_L g2636 ( 
.A(n_2284),
.Y(n_2636)
);

OAI22xp5_ASAP7_75t_L g2637 ( 
.A1(n_2404),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_2637)
);

NAND2xp33_ASAP7_75t_R g2638 ( 
.A(n_2374),
.B(n_2394),
.Y(n_2638)
);

AO21x2_ASAP7_75t_L g2639 ( 
.A1(n_2483),
.A2(n_19),
.B(n_20),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2279),
.Y(n_2640)
);

OAI21x1_ASAP7_75t_L g2641 ( 
.A1(n_2327),
.A2(n_1058),
.B(n_1044),
.Y(n_2641)
);

BUFx6f_ASAP7_75t_L g2642 ( 
.A(n_2349),
.Y(n_2642)
);

OAI21x1_ASAP7_75t_L g2643 ( 
.A1(n_2343),
.A2(n_1058),
.B(n_1044),
.Y(n_2643)
);

OAI22xp5_ASAP7_75t_L g2644 ( 
.A1(n_2297),
.A2(n_25),
.B1(n_22),
.B2(n_23),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2473),
.B(n_23),
.Y(n_2645)
);

OAI21xp5_ASAP7_75t_L g2646 ( 
.A1(n_2470),
.A2(n_1011),
.B(n_25),
.Y(n_2646)
);

INVxp67_ASAP7_75t_SL g2647 ( 
.A(n_2451),
.Y(n_2647)
);

OAI21x1_ASAP7_75t_SL g2648 ( 
.A1(n_2377),
.A2(n_26),
.B(n_27),
.Y(n_2648)
);

OA22x2_ASAP7_75t_L g2649 ( 
.A1(n_2344),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2314),
.Y(n_2650)
);

CKINVDCx20_ASAP7_75t_R g2651 ( 
.A(n_2367),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2322),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2475),
.B(n_2489),
.Y(n_2653)
);

A2O1A1Ixp33_ASAP7_75t_L g2654 ( 
.A1(n_2444),
.A2(n_31),
.B(n_28),
.C(n_30),
.Y(n_2654)
);

INVx3_ASAP7_75t_L g2655 ( 
.A(n_2387),
.Y(n_2655)
);

AOI31xp67_ASAP7_75t_L g2656 ( 
.A1(n_2287),
.A2(n_486),
.A3(n_487),
.B(n_484),
.Y(n_2656)
);

OR2x2_ASAP7_75t_L g2657 ( 
.A(n_2325),
.B(n_30),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2471),
.B(n_31),
.Y(n_2658)
);

OR2x2_ASAP7_75t_L g2659 ( 
.A(n_2496),
.B(n_32),
.Y(n_2659)
);

OAI21x1_ASAP7_75t_SL g2660 ( 
.A1(n_2331),
.A2(n_33),
.B(n_34),
.Y(n_2660)
);

OAI21x1_ASAP7_75t_L g2661 ( 
.A1(n_2371),
.A2(n_2510),
.B(n_2393),
.Y(n_2661)
);

OAI22xp5_ASAP7_75t_L g2662 ( 
.A1(n_2336),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_2662)
);

AOI21xp5_ASAP7_75t_L g2663 ( 
.A1(n_2418),
.A2(n_1002),
.B(n_996),
.Y(n_2663)
);

OAI21xp5_ASAP7_75t_L g2664 ( 
.A1(n_2508),
.A2(n_1011),
.B(n_36),
.Y(n_2664)
);

AOI21xp5_ASAP7_75t_L g2665 ( 
.A1(n_2514),
.A2(n_1002),
.B(n_996),
.Y(n_2665)
);

OAI21x1_ASAP7_75t_L g2666 ( 
.A1(n_2507),
.A2(n_1058),
.B(n_1044),
.Y(n_2666)
);

AO31x2_ASAP7_75t_L g2667 ( 
.A1(n_2521),
.A2(n_489),
.A3(n_495),
.B(n_488),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2341),
.Y(n_2668)
);

OAI21x1_ASAP7_75t_L g2669 ( 
.A1(n_2386),
.A2(n_1058),
.B(n_1044),
.Y(n_2669)
);

AO21x1_ASAP7_75t_L g2670 ( 
.A1(n_2317),
.A2(n_2504),
.B(n_2512),
.Y(n_2670)
);

A2O1A1Ixp33_ASAP7_75t_L g2671 ( 
.A1(n_2392),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_2671)
);

OAI21x1_ASAP7_75t_L g2672 ( 
.A1(n_2425),
.A2(n_1079),
.B(n_1063),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2359),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2363),
.Y(n_2674)
);

OAI21x1_ASAP7_75t_L g2675 ( 
.A1(n_2433),
.A2(n_2505),
.B(n_2307),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2472),
.B(n_37),
.Y(n_2676)
);

OAI21x1_ASAP7_75t_L g2677 ( 
.A1(n_2505),
.A2(n_1079),
.B(n_1063),
.Y(n_2677)
);

OAI21x1_ASAP7_75t_L g2678 ( 
.A1(n_2516),
.A2(n_1079),
.B(n_1063),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2364),
.Y(n_2679)
);

HB1xp67_ASAP7_75t_L g2680 ( 
.A(n_2419),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_SL g2681 ( 
.A(n_2283),
.B(n_1063),
.Y(n_2681)
);

INVxp67_ASAP7_75t_L g2682 ( 
.A(n_2421),
.Y(n_2682)
);

OAI21x1_ASAP7_75t_L g2683 ( 
.A1(n_2523),
.A2(n_2528),
.B(n_2536),
.Y(n_2683)
);

OAI21x1_ASAP7_75t_L g2684 ( 
.A1(n_2530),
.A2(n_1079),
.B(n_1063),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2500),
.B(n_38),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2453),
.B(n_39),
.Y(n_2686)
);

OR2x2_ASAP7_75t_L g2687 ( 
.A(n_2319),
.B(n_40),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2382),
.Y(n_2688)
);

NAND2x1p5_ASAP7_75t_L g2689 ( 
.A(n_2517),
.B(n_1063),
.Y(n_2689)
);

O2A1O1Ixp5_ASAP7_75t_L g2690 ( 
.A1(n_2524),
.A2(n_45),
.B(n_41),
.C(n_43),
.Y(n_2690)
);

OA21x2_ASAP7_75t_L g2691 ( 
.A1(n_2485),
.A2(n_45),
.B(n_46),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2409),
.Y(n_2692)
);

AOI21xp5_ASAP7_75t_L g2693 ( 
.A1(n_2281),
.A2(n_1002),
.B(n_996),
.Y(n_2693)
);

OA21x2_ASAP7_75t_L g2694 ( 
.A1(n_2483),
.A2(n_47),
.B(n_48),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2456),
.Y(n_2695)
);

NOR2xp33_ASAP7_75t_L g2696 ( 
.A(n_2283),
.B(n_498),
.Y(n_2696)
);

AOI22xp5_ASAP7_75t_L g2697 ( 
.A1(n_2289),
.A2(n_1085),
.B1(n_1088),
.B2(n_1079),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2305),
.B(n_47),
.Y(n_2698)
);

OAI21x1_ASAP7_75t_L g2699 ( 
.A1(n_2506),
.A2(n_1085),
.B(n_1079),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2348),
.B(n_48),
.Y(n_2700)
);

BUFx6f_ASAP7_75t_L g2701 ( 
.A(n_2387),
.Y(n_2701)
);

OAI22xp5_ASAP7_75t_L g2702 ( 
.A1(n_2285),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_2702)
);

NOR2xp33_ASAP7_75t_L g2703 ( 
.A(n_2432),
.B(n_2454),
.Y(n_2703)
);

NOR2x1_ASAP7_75t_L g2704 ( 
.A(n_2454),
.B(n_1085),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2350),
.B(n_51),
.Y(n_2705)
);

OR2x2_ASAP7_75t_L g2706 ( 
.A(n_2286),
.B(n_52),
.Y(n_2706)
);

NOR2xp33_ASAP7_75t_L g2707 ( 
.A(n_2426),
.B(n_499),
.Y(n_2707)
);

NAND3xp33_ASAP7_75t_L g2708 ( 
.A(n_2390),
.B(n_1088),
.C(n_1085),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2352),
.B(n_52),
.Y(n_2709)
);

AO31x2_ASAP7_75t_L g2710 ( 
.A1(n_2519),
.A2(n_505),
.A3(n_506),
.B(n_500),
.Y(n_2710)
);

INVx3_ASAP7_75t_L g2711 ( 
.A(n_2387),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2498),
.B(n_53),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2361),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2365),
.Y(n_2714)
);

CKINVDCx11_ASAP7_75t_R g2715 ( 
.A(n_2431),
.Y(n_2715)
);

OAI21x1_ASAP7_75t_L g2716 ( 
.A1(n_2318),
.A2(n_1088),
.B(n_1085),
.Y(n_2716)
);

AOI21xp5_ASAP7_75t_L g2717 ( 
.A1(n_2318),
.A2(n_1002),
.B(n_996),
.Y(n_2717)
);

AOI21xp5_ASAP7_75t_L g2718 ( 
.A1(n_2525),
.A2(n_1002),
.B(n_996),
.Y(n_2718)
);

NAND2x1p5_ASAP7_75t_L g2719 ( 
.A(n_2517),
.B(n_1085),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2291),
.B(n_53),
.Y(n_2720)
);

OAI22xp5_ASAP7_75t_L g2721 ( 
.A1(n_2517),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2291),
.B(n_55),
.Y(n_2722)
);

BUFx2_ASAP7_75t_L g2723 ( 
.A(n_2387),
.Y(n_2723)
);

OAI22xp5_ASAP7_75t_L g2724 ( 
.A1(n_2534),
.A2(n_60),
.B1(n_57),
.B2(n_59),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2398),
.B(n_2337),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2388),
.Y(n_2726)
);

AOI21xp5_ASAP7_75t_L g2727 ( 
.A1(n_2384),
.A2(n_996),
.B(n_1011),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_SL g2728 ( 
.A(n_2431),
.B(n_1088),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_2400),
.Y(n_2729)
);

NOR3xp33_ASAP7_75t_SL g2730 ( 
.A(n_2303),
.B(n_57),
.C(n_59),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2398),
.B(n_61),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2337),
.B(n_61),
.Y(n_2732)
);

OAI21xp5_ASAP7_75t_L g2733 ( 
.A1(n_2429),
.A2(n_1011),
.B(n_62),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2345),
.B(n_63),
.Y(n_2734)
);

NOR2xp33_ASAP7_75t_L g2735 ( 
.A(n_2480),
.B(n_509),
.Y(n_2735)
);

AOI21xp5_ASAP7_75t_L g2736 ( 
.A1(n_2526),
.A2(n_1011),
.B(n_1088),
.Y(n_2736)
);

NAND3xp33_ASAP7_75t_L g2737 ( 
.A(n_2346),
.B(n_1097),
.C(n_1088),
.Y(n_2737)
);

INVx5_ASAP7_75t_L g2738 ( 
.A(n_2385),
.Y(n_2738)
);

INVx3_ASAP7_75t_SL g2739 ( 
.A(n_2304),
.Y(n_2739)
);

AOI21xp5_ASAP7_75t_L g2740 ( 
.A1(n_2531),
.A2(n_1011),
.B(n_1097),
.Y(n_2740)
);

OAI21xp5_ASAP7_75t_L g2741 ( 
.A1(n_2317),
.A2(n_63),
.B(n_64),
.Y(n_2741)
);

AO22x2_ASAP7_75t_L g2742 ( 
.A1(n_2303),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2345),
.B(n_65),
.Y(n_2743)
);

OR2x2_ASAP7_75t_L g2744 ( 
.A(n_2477),
.B(n_67),
.Y(n_2744)
);

AOI21x1_ASAP7_75t_L g2745 ( 
.A1(n_2533),
.A2(n_1110),
.B(n_1097),
.Y(n_2745)
);

AO21x2_ASAP7_75t_L g2746 ( 
.A1(n_2474),
.A2(n_68),
.B(n_69),
.Y(n_2746)
);

NAND2xp33_ASAP7_75t_L g2747 ( 
.A(n_2374),
.B(n_1097),
.Y(n_2747)
);

HB1xp67_ASAP7_75t_L g2748 ( 
.A(n_2484),
.Y(n_2748)
);

OAI21x1_ASAP7_75t_L g2749 ( 
.A1(n_2541),
.A2(n_1110),
.B(n_1097),
.Y(n_2749)
);

AO32x2_ASAP7_75t_L g2750 ( 
.A1(n_2493),
.A2(n_70),
.A3(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_2750)
);

NAND3x1_ASAP7_75t_L g2751 ( 
.A(n_2455),
.B(n_2402),
.C(n_2421),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2380),
.B(n_70),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2370),
.B(n_71),
.Y(n_2753)
);

BUFx6f_ASAP7_75t_L g2754 ( 
.A(n_2414),
.Y(n_2754)
);

AO32x2_ASAP7_75t_L g2755 ( 
.A1(n_2405),
.A2(n_74),
.A3(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_2755)
);

CKINVDCx20_ASAP7_75t_R g2756 ( 
.A(n_2513),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_L g2757 ( 
.A(n_2333),
.B(n_510),
.Y(n_2757)
);

NAND3x1_ASAP7_75t_L g2758 ( 
.A(n_2401),
.B(n_74),
.C(n_76),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2292),
.Y(n_2759)
);

AND2x4_ASAP7_75t_L g2760 ( 
.A(n_2340),
.B(n_512),
.Y(n_2760)
);

OAI21x1_ASAP7_75t_L g2761 ( 
.A1(n_2476),
.A2(n_1110),
.B(n_1097),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2328),
.B(n_513),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2375),
.B(n_76),
.Y(n_2763)
);

AND2x2_ASAP7_75t_L g2764 ( 
.A(n_2328),
.B(n_514),
.Y(n_2764)
);

INVxp67_ASAP7_75t_SL g2765 ( 
.A(n_2320),
.Y(n_2765)
);

INVx3_ASAP7_75t_L g2766 ( 
.A(n_2414),
.Y(n_2766)
);

INVx1_ASAP7_75t_SL g2767 ( 
.A(n_2338),
.Y(n_2767)
);

OAI21xp33_ASAP7_75t_L g2768 ( 
.A1(n_2396),
.A2(n_1110),
.B(n_1111),
.Y(n_2768)
);

NOR2xp33_ASAP7_75t_L g2769 ( 
.A(n_2357),
.B(n_2381),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2399),
.B(n_2295),
.Y(n_2770)
);

CKINVDCx5p33_ASAP7_75t_R g2771 ( 
.A(n_2410),
.Y(n_2771)
);

INVxp67_ASAP7_75t_L g2772 ( 
.A(n_2416),
.Y(n_2772)
);

NAND2x1p5_ASAP7_75t_L g2773 ( 
.A(n_2436),
.B(n_1110),
.Y(n_2773)
);

OAI21x1_ASAP7_75t_L g2774 ( 
.A1(n_2499),
.A2(n_1111),
.B(n_1110),
.Y(n_2774)
);

OAI21x1_ASAP7_75t_L g2775 ( 
.A1(n_2499),
.A2(n_2492),
.B(n_2491),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2380),
.B(n_78),
.Y(n_2776)
);

OR2x2_ASAP7_75t_L g2777 ( 
.A(n_2408),
.B(n_78),
.Y(n_2777)
);

AOI22xp5_ASAP7_75t_L g2778 ( 
.A1(n_2515),
.A2(n_1111),
.B1(n_1060),
.B2(n_1098),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2357),
.B(n_79),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2395),
.Y(n_2780)
);

NOR2xp33_ASAP7_75t_SL g2781 ( 
.A(n_2378),
.B(n_80),
.Y(n_2781)
);

NOR2xp67_ASAP7_75t_L g2782 ( 
.A(n_2296),
.B(n_80),
.Y(n_2782)
);

BUFx6f_ASAP7_75t_L g2783 ( 
.A(n_2414),
.Y(n_2783)
);

OAI22xp5_ASAP7_75t_L g2784 ( 
.A1(n_2434),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_2784)
);

OAI21x1_ASAP7_75t_L g2785 ( 
.A1(n_2428),
.A2(n_1111),
.B(n_1060),
.Y(n_2785)
);

NOR2xp67_ASAP7_75t_SL g2786 ( 
.A(n_2497),
.B(n_1111),
.Y(n_2786)
);

AO32x2_ASAP7_75t_L g2787 ( 
.A1(n_2430),
.A2(n_85),
.A3(n_81),
.B1(n_84),
.B2(n_86),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2397),
.B(n_2320),
.Y(n_2788)
);

INVx1_ASAP7_75t_SL g2789 ( 
.A(n_2488),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2412),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2435),
.Y(n_2791)
);

HB1xp67_ASAP7_75t_L g2792 ( 
.A(n_2478),
.Y(n_2792)
);

BUFx3_ASAP7_75t_L g2793 ( 
.A(n_2513),
.Y(n_2793)
);

AOI21xp5_ASAP7_75t_L g2794 ( 
.A1(n_2397),
.A2(n_2347),
.B(n_2535),
.Y(n_2794)
);

AOI22xp5_ASAP7_75t_L g2795 ( 
.A1(n_2467),
.A2(n_1111),
.B1(n_1060),
.B2(n_1098),
.Y(n_2795)
);

OAI22xp5_ASAP7_75t_L g2796 ( 
.A1(n_2448),
.A2(n_90),
.B1(n_84),
.B2(n_87),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2452),
.Y(n_2797)
);

A2O1A1Ixp33_ASAP7_75t_L g2798 ( 
.A1(n_2282),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_2798)
);

AND2x4_ASAP7_75t_L g2799 ( 
.A(n_2372),
.B(n_92),
.Y(n_2799)
);

BUFx6f_ASAP7_75t_L g2800 ( 
.A(n_2414),
.Y(n_2800)
);

NOR2xp33_ASAP7_75t_SL g2801 ( 
.A(n_2448),
.B(n_94),
.Y(n_2801)
);

OA21x2_ASAP7_75t_L g2802 ( 
.A1(n_2543),
.A2(n_2474),
.B(n_2520),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2725),
.B(n_2417),
.Y(n_2803)
);

NOR2xp33_ASAP7_75t_SL g2804 ( 
.A(n_2614),
.B(n_2296),
.Y(n_2804)
);

NOR2xp33_ASAP7_75t_L g2805 ( 
.A(n_2682),
.B(n_2294),
.Y(n_2805)
);

INVx4_ASAP7_75t_L g2806 ( 
.A(n_2556),
.Y(n_2806)
);

INVx3_ASAP7_75t_L g2807 ( 
.A(n_2775),
.Y(n_2807)
);

OAI21x1_ASAP7_75t_L g2808 ( 
.A1(n_2576),
.A2(n_2428),
.B(n_2372),
.Y(n_2808)
);

OA21x2_ASAP7_75t_L g2809 ( 
.A1(n_2544),
.A2(n_2511),
.B(n_2490),
.Y(n_2809)
);

AND2x2_ASAP7_75t_L g2810 ( 
.A(n_2640),
.B(n_2406),
.Y(n_2810)
);

OAI21x1_ASAP7_75t_L g2811 ( 
.A1(n_2605),
.A2(n_2542),
.B(n_2629),
.Y(n_2811)
);

NAND3xp33_ASAP7_75t_L g2812 ( 
.A(n_2703),
.B(n_2490),
.C(n_2537),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2650),
.Y(n_2813)
);

OAI21x1_ASAP7_75t_L g2814 ( 
.A1(n_2661),
.A2(n_2324),
.B(n_2406),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2546),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2552),
.Y(n_2816)
);

OA21x2_ASAP7_75t_L g2817 ( 
.A1(n_2675),
.A2(n_2479),
.B(n_2462),
.Y(n_2817)
);

BUFx3_ASAP7_75t_L g2818 ( 
.A(n_2626),
.Y(n_2818)
);

OA21x2_ASAP7_75t_L g2819 ( 
.A1(n_2699),
.A2(n_2446),
.B(n_2347),
.Y(n_2819)
);

OA21x2_ASAP7_75t_L g2820 ( 
.A1(n_2684),
.A2(n_2535),
.B(n_2441),
.Y(n_2820)
);

NOR2x1_ASAP7_75t_SL g2821 ( 
.A(n_2556),
.B(n_2613),
.Y(n_2821)
);

AOI21xp5_ASAP7_75t_L g2822 ( 
.A1(n_2592),
.A2(n_2522),
.B(n_2482),
.Y(n_2822)
);

OA21x2_ASAP7_75t_L g2823 ( 
.A1(n_2643),
.A2(n_2460),
.B(n_2457),
.Y(n_2823)
);

OAI21x1_ASAP7_75t_L g2824 ( 
.A1(n_2632),
.A2(n_2440),
.B(n_2461),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2561),
.Y(n_2825)
);

AO31x2_ASAP7_75t_L g2826 ( 
.A1(n_2663),
.A2(n_2482),
.A3(n_2436),
.B(n_2376),
.Y(n_2826)
);

INVx3_ASAP7_75t_L g2827 ( 
.A(n_2555),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2573),
.Y(n_2828)
);

OA21x2_ASAP7_75t_L g2829 ( 
.A1(n_2560),
.A2(n_2381),
.B(n_2424),
.Y(n_2829)
);

CKINVDCx5p33_ASAP7_75t_R g2830 ( 
.A(n_2651),
.Y(n_2830)
);

AND2x4_ASAP7_75t_L g2831 ( 
.A(n_2582),
.B(n_2495),
.Y(n_2831)
);

OR2x6_ASAP7_75t_L g2832 ( 
.A(n_2567),
.B(n_2522),
.Y(n_2832)
);

OR2x6_ASAP7_75t_L g2833 ( 
.A(n_2794),
.B(n_2522),
.Y(n_2833)
);

AO21x1_ASAP7_75t_L g2834 ( 
.A1(n_2662),
.A2(n_2702),
.B(n_2741),
.Y(n_2834)
);

INVx6_ASAP7_75t_L g2835 ( 
.A(n_2627),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2602),
.Y(n_2836)
);

OAI22xp5_ASAP7_75t_L g2837 ( 
.A1(n_2751),
.A2(n_2478),
.B1(n_2329),
.B2(n_2376),
.Y(n_2837)
);

OAI21x1_ASAP7_75t_L g2838 ( 
.A1(n_2633),
.A2(n_2641),
.B(n_2669),
.Y(n_2838)
);

OAI21x1_ASAP7_75t_L g2839 ( 
.A1(n_2666),
.A2(n_2509),
.B(n_2478),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2607),
.Y(n_2840)
);

OAI21x1_ASAP7_75t_L g2841 ( 
.A1(n_2604),
.A2(n_2509),
.B(n_2478),
.Y(n_2841)
);

HB1xp67_ASAP7_75t_L g2842 ( 
.A(n_2748),
.Y(n_2842)
);

AO21x2_ASAP7_75t_L g2843 ( 
.A1(n_2560),
.A2(n_2413),
.B(n_2509),
.Y(n_2843)
);

AOI21xp5_ASAP7_75t_L g2844 ( 
.A1(n_2646),
.A2(n_2664),
.B(n_2708),
.Y(n_2844)
);

AOI21xp5_ASAP7_75t_L g2845 ( 
.A1(n_2646),
.A2(n_2413),
.B(n_2439),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2621),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2652),
.Y(n_2847)
);

OAI21x1_ASAP7_75t_L g2848 ( 
.A1(n_2672),
.A2(n_2439),
.B(n_2427),
.Y(n_2848)
);

OAI21x1_ASAP7_75t_L g2849 ( 
.A1(n_2603),
.A2(n_2678),
.B(n_2749),
.Y(n_2849)
);

INVx6_ASAP7_75t_L g2850 ( 
.A(n_2627),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2668),
.Y(n_2851)
);

AOI22xp5_ASAP7_75t_L g2852 ( 
.A1(n_2801),
.A2(n_2311),
.B1(n_2329),
.B2(n_2439),
.Y(n_2852)
);

OAI21x1_ASAP7_75t_L g2853 ( 
.A1(n_2683),
.A2(n_2439),
.B(n_2427),
.Y(n_2853)
);

BUFx6f_ASAP7_75t_L g2854 ( 
.A(n_2627),
.Y(n_2854)
);

OAI21x1_ASAP7_75t_L g2855 ( 
.A1(n_2677),
.A2(n_2665),
.B(n_2716),
.Y(n_2855)
);

OAI21x1_ASAP7_75t_L g2856 ( 
.A1(n_2559),
.A2(n_2427),
.B(n_94),
.Y(n_2856)
);

OAI21x1_ASAP7_75t_L g2857 ( 
.A1(n_2745),
.A2(n_2427),
.B(n_95),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2673),
.Y(n_2858)
);

OAI21x1_ASAP7_75t_SL g2859 ( 
.A1(n_2741),
.A2(n_95),
.B(n_96),
.Y(n_2859)
);

OAI21x1_ASAP7_75t_L g2860 ( 
.A1(n_2557),
.A2(n_97),
.B(n_98),
.Y(n_2860)
);

A2O1A1Ixp33_ASAP7_75t_L g2861 ( 
.A1(n_2733),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2674),
.Y(n_2862)
);

AND2x2_ASAP7_75t_L g2863 ( 
.A(n_2679),
.B(n_2688),
.Y(n_2863)
);

CKINVDCx8_ASAP7_75t_R g2864 ( 
.A(n_2771),
.Y(n_2864)
);

OAI21x1_ASAP7_75t_L g2865 ( 
.A1(n_2562),
.A2(n_100),
.B(n_101),
.Y(n_2865)
);

A2O1A1Ixp33_ASAP7_75t_L g2866 ( 
.A1(n_2733),
.A2(n_102),
.B(n_100),
.C(n_101),
.Y(n_2866)
);

NOR2xp33_ASAP7_75t_L g2867 ( 
.A(n_2772),
.B(n_102),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2692),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2593),
.Y(n_2869)
);

OAI21xp5_ASAP7_75t_L g2870 ( 
.A1(n_2664),
.A2(n_103),
.B(n_104),
.Y(n_2870)
);

OAI21x1_ASAP7_75t_L g2871 ( 
.A1(n_2774),
.A2(n_103),
.B(n_105),
.Y(n_2871)
);

HB1xp67_ASAP7_75t_L g2872 ( 
.A(n_2680),
.Y(n_2872)
);

AO21x2_ASAP7_75t_L g2873 ( 
.A1(n_2591),
.A2(n_105),
.B(n_106),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2647),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2570),
.Y(n_2875)
);

BUFx3_ASAP7_75t_L g2876 ( 
.A(n_2723),
.Y(n_2876)
);

AND2x2_ASAP7_75t_L g2877 ( 
.A(n_2695),
.B(n_107),
.Y(n_2877)
);

OR2x2_ASAP7_75t_L g2878 ( 
.A(n_2725),
.B(n_108),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2713),
.Y(n_2879)
);

OAI21x1_ASAP7_75t_L g2880 ( 
.A1(n_2585),
.A2(n_109),
.B(n_110),
.Y(n_2880)
);

HB1xp67_ASAP7_75t_L g2881 ( 
.A(n_2767),
.Y(n_2881)
);

OAI21x1_ASAP7_75t_L g2882 ( 
.A1(n_2611),
.A2(n_109),
.B(n_112),
.Y(n_2882)
);

OAI22xp5_ASAP7_75t_L g2883 ( 
.A1(n_2583),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_2883)
);

OAI21x1_ASAP7_75t_L g2884 ( 
.A1(n_2761),
.A2(n_114),
.B(n_115),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2714),
.Y(n_2885)
);

AO32x2_ASAP7_75t_L g2886 ( 
.A1(n_2662),
.A2(n_120),
.A3(n_116),
.B1(n_118),
.B2(n_121),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2726),
.Y(n_2887)
);

OAI21x1_ASAP7_75t_L g2888 ( 
.A1(n_2547),
.A2(n_116),
.B(n_118),
.Y(n_2888)
);

OAI21xp5_ASAP7_75t_L g2889 ( 
.A1(n_2708),
.A2(n_122),
.B(n_123),
.Y(n_2889)
);

A2O1A1Ixp33_ASAP7_75t_L g2890 ( 
.A1(n_2801),
.A2(n_124),
.B(n_122),
.C(n_123),
.Y(n_2890)
);

OAI21x1_ASAP7_75t_L g2891 ( 
.A1(n_2545),
.A2(n_124),
.B(n_125),
.Y(n_2891)
);

AOI221xp5_ASAP7_75t_L g2892 ( 
.A1(n_2724),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.C(n_129),
.Y(n_2892)
);

OAI21x1_ASAP7_75t_L g2893 ( 
.A1(n_2785),
.A2(n_126),
.B(n_127),
.Y(n_2893)
);

INVx1_ASAP7_75t_SL g2894 ( 
.A(n_2729),
.Y(n_2894)
);

OAI21x1_ASAP7_75t_L g2895 ( 
.A1(n_2717),
.A2(n_130),
.B(n_131),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2765),
.B(n_130),
.Y(n_2896)
);

BUFx3_ASAP7_75t_L g2897 ( 
.A(n_2701),
.Y(n_2897)
);

BUFx6f_ASAP7_75t_L g2898 ( 
.A(n_2642),
.Y(n_2898)
);

INVx2_ASAP7_75t_L g2899 ( 
.A(n_2790),
.Y(n_2899)
);

AOI22xp33_ASAP7_75t_L g2900 ( 
.A1(n_2724),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_2900)
);

O2A1O1Ixp33_ASAP7_75t_L g2901 ( 
.A1(n_2654),
.A2(n_134),
.B(n_132),
.C(n_133),
.Y(n_2901)
);

AND2x4_ASAP7_75t_L g2902 ( 
.A(n_2556),
.B(n_134),
.Y(n_2902)
);

HB1xp67_ASAP7_75t_L g2903 ( 
.A(n_2767),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2797),
.Y(n_2904)
);

OAI21x1_ASAP7_75t_L g2905 ( 
.A1(n_2558),
.A2(n_136),
.B(n_139),
.Y(n_2905)
);

AOI21xp5_ASAP7_75t_L g2906 ( 
.A1(n_2727),
.A2(n_136),
.B(n_139),
.Y(n_2906)
);

NOR2xp67_ASAP7_75t_L g2907 ( 
.A(n_2553),
.B(n_140),
.Y(n_2907)
);

BUFx3_ASAP7_75t_L g2908 ( 
.A(n_2701),
.Y(n_2908)
);

CKINVDCx20_ASAP7_75t_R g2909 ( 
.A(n_2756),
.Y(n_2909)
);

OAI21xp5_ASAP7_75t_L g2910 ( 
.A1(n_2798),
.A2(n_140),
.B(n_142),
.Y(n_2910)
);

OAI21x1_ASAP7_75t_L g2911 ( 
.A1(n_2554),
.A2(n_143),
.B(n_144),
.Y(n_2911)
);

OAI21x1_ASAP7_75t_L g2912 ( 
.A1(n_2554),
.A2(n_145),
.B(n_146),
.Y(n_2912)
);

AOI22xp33_ASAP7_75t_L g2913 ( 
.A1(n_2615),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_2913)
);

AO31x2_ASAP7_75t_L g2914 ( 
.A1(n_2702),
.A2(n_150),
.A3(n_148),
.B(n_149),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2571),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2788),
.B(n_150),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2625),
.Y(n_2917)
);

INVx2_ASAP7_75t_L g2918 ( 
.A(n_2759),
.Y(n_2918)
);

OAI21xp33_ASAP7_75t_L g2919 ( 
.A1(n_2730),
.A2(n_152),
.B(n_153),
.Y(n_2919)
);

OAI21x1_ASAP7_75t_L g2920 ( 
.A1(n_2693),
.A2(n_152),
.B(n_153),
.Y(n_2920)
);

OR2x6_ASAP7_75t_L g2921 ( 
.A(n_2575),
.B(n_1027),
.Y(n_2921)
);

OA21x2_ASAP7_75t_L g2922 ( 
.A1(n_2599),
.A2(n_154),
.B(n_155),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2788),
.B(n_2653),
.Y(n_2923)
);

AND2x4_ASAP7_75t_L g2924 ( 
.A(n_2613),
.B(n_154),
.Y(n_2924)
);

BUFx8_ASAP7_75t_L g2925 ( 
.A(n_2642),
.Y(n_2925)
);

OAI21x1_ASAP7_75t_L g2926 ( 
.A1(n_2590),
.A2(n_156),
.B(n_157),
.Y(n_2926)
);

OA21x2_ASAP7_75t_L g2927 ( 
.A1(n_2712),
.A2(n_156),
.B(n_157),
.Y(n_2927)
);

NAND3xp33_ASAP7_75t_L g2928 ( 
.A(n_2712),
.B(n_158),
.C(n_159),
.Y(n_2928)
);

NAND2x1p5_ASAP7_75t_L g2929 ( 
.A(n_2613),
.B(n_158),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2780),
.Y(n_2930)
);

INVx2_ASAP7_75t_SL g2931 ( 
.A(n_2792),
.Y(n_2931)
);

OAI21x1_ASAP7_75t_L g2932 ( 
.A1(n_2584),
.A2(n_160),
.B(n_161),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2791),
.Y(n_2933)
);

OAI21x1_ASAP7_75t_L g2934 ( 
.A1(n_2564),
.A2(n_160),
.B(n_161),
.Y(n_2934)
);

AND2x2_ASAP7_75t_L g2935 ( 
.A(n_2548),
.B(n_2586),
.Y(n_2935)
);

OAI21x1_ASAP7_75t_L g2936 ( 
.A1(n_2568),
.A2(n_163),
.B(n_164),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2586),
.Y(n_2937)
);

OAI21x1_ASAP7_75t_L g2938 ( 
.A1(n_2736),
.A2(n_165),
.B(n_166),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2686),
.Y(n_2939)
);

INVx3_ASAP7_75t_L g2940 ( 
.A(n_2738),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2686),
.Y(n_2941)
);

AND2x4_ASAP7_75t_L g2942 ( 
.A(n_2738),
.B(n_165),
.Y(n_2942)
);

OA21x2_ASAP7_75t_L g2943 ( 
.A1(n_2690),
.A2(n_166),
.B(n_168),
.Y(n_2943)
);

BUFx3_ASAP7_75t_L g2944 ( 
.A(n_2701),
.Y(n_2944)
);

OA21x2_ASAP7_75t_L g2945 ( 
.A1(n_2670),
.A2(n_168),
.B(n_169),
.Y(n_2945)
);

OAI22xp33_ASAP7_75t_L g2946 ( 
.A1(n_2609),
.A2(n_172),
.B1(n_169),
.B2(n_171),
.Y(n_2946)
);

AND2x4_ASAP7_75t_L g2947 ( 
.A(n_2738),
.B(n_172),
.Y(n_2947)
);

BUFx4f_ASAP7_75t_L g2948 ( 
.A(n_2642),
.Y(n_2948)
);

OAI21x1_ASAP7_75t_L g2949 ( 
.A1(n_2740),
.A2(n_173),
.B(n_174),
.Y(n_2949)
);

INVx2_ASAP7_75t_SL g2950 ( 
.A(n_2600),
.Y(n_2950)
);

AND2x2_ASAP7_75t_L g2951 ( 
.A(n_2586),
.B(n_176),
.Y(n_2951)
);

OAI21xp5_ASAP7_75t_L g2952 ( 
.A1(n_2704),
.A2(n_177),
.B(n_179),
.Y(n_2952)
);

INVxp67_ASAP7_75t_SL g2953 ( 
.A(n_2579),
.Y(n_2953)
);

INVx2_ASAP7_75t_SL g2954 ( 
.A(n_2789),
.Y(n_2954)
);

AND2x2_ASAP7_75t_L g2955 ( 
.A(n_2580),
.B(n_181),
.Y(n_2955)
);

OAI21x1_ASAP7_75t_L g2956 ( 
.A1(n_2718),
.A2(n_182),
.B(n_184),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2698),
.Y(n_2957)
);

OAI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_2707),
.A2(n_185),
.B(n_186),
.Y(n_2958)
);

HB1xp67_ASAP7_75t_L g2959 ( 
.A(n_2789),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2770),
.B(n_186),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2698),
.Y(n_2961)
);

CKINVDCx8_ASAP7_75t_R g2962 ( 
.A(n_2754),
.Y(n_2962)
);

AND2x4_ASAP7_75t_L g2963 ( 
.A(n_2655),
.B(n_187),
.Y(n_2963)
);

OAI21x1_ASAP7_75t_L g2964 ( 
.A1(n_2608),
.A2(n_187),
.B(n_188),
.Y(n_2964)
);

A2O1A1Ixp33_ASAP7_75t_L g2965 ( 
.A1(n_2781),
.A2(n_191),
.B(n_189),
.C(n_190),
.Y(n_2965)
);

HB1xp67_ASAP7_75t_L g2966 ( 
.A(n_2580),
.Y(n_2966)
);

BUFx3_ASAP7_75t_L g2967 ( 
.A(n_2754),
.Y(n_2967)
);

INVx2_ASAP7_75t_L g2968 ( 
.A(n_2623),
.Y(n_2968)
);

OAI21x1_ASAP7_75t_L g2969 ( 
.A1(n_2601),
.A2(n_2719),
.B(n_2689),
.Y(n_2969)
);

INVx2_ASAP7_75t_SL g2970 ( 
.A(n_2754),
.Y(n_2970)
);

BUFx2_ASAP7_75t_L g2971 ( 
.A(n_2580),
.Y(n_2971)
);

OAI22xp5_ASAP7_75t_L g2972 ( 
.A1(n_2644),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_2972)
);

AO21x2_ASAP7_75t_L g2973 ( 
.A1(n_2591),
.A2(n_192),
.B(n_193),
.Y(n_2973)
);

BUFx2_ASAP7_75t_R g2974 ( 
.A(n_2793),
.Y(n_2974)
);

AOI21xp33_ASAP7_75t_L g2975 ( 
.A1(n_2635),
.A2(n_2746),
.B(n_2747),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2700),
.Y(n_2976)
);

OAI21x1_ASAP7_75t_L g2977 ( 
.A1(n_2689),
.A2(n_194),
.B(n_195),
.Y(n_2977)
);

NOR2xp33_ASAP7_75t_L g2978 ( 
.A(n_2769),
.B(n_194),
.Y(n_2978)
);

NOR2xp33_ASAP7_75t_L g2979 ( 
.A(n_2636),
.B(n_2696),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2700),
.Y(n_2980)
);

AND2x4_ASAP7_75t_L g2981 ( 
.A(n_2655),
.B(n_195),
.Y(n_2981)
);

OAI21x1_ASAP7_75t_L g2982 ( 
.A1(n_2719),
.A2(n_196),
.B(n_197),
.Y(n_2982)
);

OAI21x1_ASAP7_75t_L g2983 ( 
.A1(n_2694),
.A2(n_2691),
.B(n_2589),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2623),
.Y(n_2984)
);

AOI22xp33_ASAP7_75t_L g2985 ( 
.A1(n_2615),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_2985)
);

OAI21x1_ASAP7_75t_L g2986 ( 
.A1(n_2694),
.A2(n_200),
.B(n_201),
.Y(n_2986)
);

OA21x2_ASAP7_75t_L g2987 ( 
.A1(n_2737),
.A2(n_200),
.B(n_202),
.Y(n_2987)
);

AND2x4_ASAP7_75t_L g2988 ( 
.A(n_2711),
.B(n_202),
.Y(n_2988)
);

O2A1O1Ixp33_ASAP7_75t_L g2989 ( 
.A1(n_2671),
.A2(n_2595),
.B(n_2796),
.C(n_2637),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_2566),
.B(n_203),
.Y(n_2990)
);

AO31x2_ASAP7_75t_L g2991 ( 
.A1(n_2644),
.A2(n_205),
.A3(n_203),
.B(n_204),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2705),
.Y(n_2992)
);

OAI21xp33_ASAP7_75t_SL g2993 ( 
.A1(n_2649),
.A2(n_206),
.B(n_207),
.Y(n_2993)
);

O2A1O1Ixp33_ASAP7_75t_L g2994 ( 
.A1(n_2796),
.A2(n_208),
.B(n_206),
.C(n_207),
.Y(n_2994)
);

BUFx6f_ASAP7_75t_L g2995 ( 
.A(n_2783),
.Y(n_2995)
);

OAI21xp5_ASAP7_75t_L g2996 ( 
.A1(n_2550),
.A2(n_208),
.B(n_209),
.Y(n_2996)
);

OAI21x1_ASAP7_75t_L g2997 ( 
.A1(n_2691),
.A2(n_210),
.B(n_211),
.Y(n_2997)
);

AO21x2_ASAP7_75t_L g2998 ( 
.A1(n_2648),
.A2(n_210),
.B(n_211),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2623),
.Y(n_2999)
);

OAI22xp33_ASAP7_75t_L g3000 ( 
.A1(n_2609),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_3000)
);

OAI21xp5_ASAP7_75t_L g3001 ( 
.A1(n_2735),
.A2(n_212),
.B(n_213),
.Y(n_3001)
);

AOI22xp33_ASAP7_75t_L g3002 ( 
.A1(n_2637),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.Y(n_3002)
);

AND2x2_ASAP7_75t_L g3003 ( 
.A(n_2705),
.B(n_215),
.Y(n_3003)
);

AND2x2_ASAP7_75t_L g3004 ( 
.A(n_2706),
.B(n_217),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2606),
.Y(n_3005)
);

A2O1A1Ixp33_ASAP7_75t_SL g3006 ( 
.A1(n_2784),
.A2(n_2786),
.B(n_2598),
.C(n_2757),
.Y(n_3006)
);

OAI21x1_ASAP7_75t_L g3007 ( 
.A1(n_2773),
.A2(n_217),
.B(n_218),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2587),
.Y(n_3008)
);

INVxp67_ASAP7_75t_L g3009 ( 
.A(n_2549),
.Y(n_3009)
);

HB1xp67_ASAP7_75t_L g3010 ( 
.A(n_2711),
.Y(n_3010)
);

AOI21xp33_ASAP7_75t_L g3011 ( 
.A1(n_2746),
.A2(n_219),
.B(n_220),
.Y(n_3011)
);

BUFx6f_ASAP7_75t_L g3012 ( 
.A(n_2783),
.Y(n_3012)
);

NAND2x1p5_ASAP7_75t_L g3013 ( 
.A(n_2620),
.B(n_219),
.Y(n_3013)
);

AOI21x1_ASAP7_75t_L g3014 ( 
.A1(n_2681),
.A2(n_222),
.B(n_223),
.Y(n_3014)
);

OAI22xp5_ASAP7_75t_SL g3015 ( 
.A1(n_2739),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_3015)
);

OAI21x1_ASAP7_75t_L g3016 ( 
.A1(n_2773),
.A2(n_224),
.B(n_225),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2587),
.Y(n_3017)
);

BUFx2_ASAP7_75t_SL g3018 ( 
.A(n_2800),
.Y(n_3018)
);

INVx2_ASAP7_75t_L g3019 ( 
.A(n_2606),
.Y(n_3019)
);

OAI21x1_ASAP7_75t_L g3020 ( 
.A1(n_2766),
.A2(n_226),
.B(n_227),
.Y(n_3020)
);

OAI21x1_ASAP7_75t_L g3021 ( 
.A1(n_2766),
.A2(n_228),
.B(n_229),
.Y(n_3021)
);

INVxp67_ASAP7_75t_L g3022 ( 
.A(n_2645),
.Y(n_3022)
);

OAI21x1_ASAP7_75t_L g3023 ( 
.A1(n_2732),
.A2(n_228),
.B(n_229),
.Y(n_3023)
);

OAI21x1_ASAP7_75t_L g3024 ( 
.A1(n_2732),
.A2(n_230),
.B(n_231),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2606),
.Y(n_3025)
);

BUFx2_ASAP7_75t_L g3026 ( 
.A(n_2876),
.Y(n_3026)
);

AOI22xp33_ASAP7_75t_L g3027 ( 
.A1(n_2870),
.A2(n_2594),
.B1(n_2577),
.B2(n_2572),
.Y(n_3027)
);

CKINVDCx11_ASAP7_75t_R g3028 ( 
.A(n_2864),
.Y(n_3028)
);

INVx3_ASAP7_75t_L g3029 ( 
.A(n_2807),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2813),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_2813),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2881),
.B(n_2657),
.Y(n_3032)
);

CKINVDCx20_ASAP7_75t_R g3033 ( 
.A(n_2909),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2847),
.Y(n_3034)
);

INVx2_ASAP7_75t_SL g3035 ( 
.A(n_2876),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2847),
.Y(n_3036)
);

OAI21x1_ASAP7_75t_L g3037 ( 
.A1(n_2811),
.A2(n_2743),
.B(n_2734),
.Y(n_3037)
);

AOI21x1_ASAP7_75t_L g3038 ( 
.A1(n_2837),
.A2(n_2742),
.B(n_2722),
.Y(n_3038)
);

BUFx8_ASAP7_75t_L g3039 ( 
.A(n_2902),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2858),
.Y(n_3040)
);

NAND2x1p5_ASAP7_75t_L g3041 ( 
.A(n_2829),
.B(n_2620),
.Y(n_3041)
);

OR2x2_ASAP7_75t_L g3042 ( 
.A(n_2903),
.B(n_2581),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2858),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2862),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2862),
.Y(n_3045)
);

OAI22xp33_ASAP7_75t_L g3046 ( 
.A1(n_2812),
.A2(n_2781),
.B1(n_2577),
.B2(n_2572),
.Y(n_3046)
);

OAI21x1_ASAP7_75t_L g3047 ( 
.A1(n_2811),
.A2(n_2743),
.B(n_2734),
.Y(n_3047)
);

INVx3_ASAP7_75t_L g3048 ( 
.A(n_2807),
.Y(n_3048)
);

OAI21x1_ASAP7_75t_L g3049 ( 
.A1(n_2855),
.A2(n_2728),
.B(n_2660),
.Y(n_3049)
);

AOI22xp33_ASAP7_75t_L g3050 ( 
.A1(n_2834),
.A2(n_2784),
.B1(n_2742),
.B2(n_2721),
.Y(n_3050)
);

INVx2_ASAP7_75t_L g3051 ( 
.A(n_2879),
.Y(n_3051)
);

AOI22xp33_ASAP7_75t_L g3052 ( 
.A1(n_2834),
.A2(n_2721),
.B1(n_2722),
.B2(n_2720),
.Y(n_3052)
);

OA21x2_ASAP7_75t_L g3053 ( 
.A1(n_2975),
.A2(n_2731),
.B(n_2752),
.Y(n_3053)
);

AOI222xp33_ASAP7_75t_L g3054 ( 
.A1(n_2958),
.A2(n_2753),
.B1(n_2763),
.B2(n_2720),
.C1(n_2622),
.C2(n_2634),
.Y(n_3054)
);

CKINVDCx5p33_ASAP7_75t_R g3055 ( 
.A(n_2830),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_2842),
.B(n_2715),
.Y(n_3056)
);

OR2x2_ASAP7_75t_L g3057 ( 
.A(n_2872),
.B(n_2709),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2851),
.Y(n_3058)
);

BUFx2_ASAP7_75t_L g3059 ( 
.A(n_2959),
.Y(n_3059)
);

CKINVDCx20_ASAP7_75t_R g3060 ( 
.A(n_2909),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2868),
.Y(n_3061)
);

INVx3_ASAP7_75t_L g3062 ( 
.A(n_2807),
.Y(n_3062)
);

INVx1_ASAP7_75t_SL g3063 ( 
.A(n_2818),
.Y(n_3063)
);

OAI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_2900),
.A2(n_2758),
.B1(n_2618),
.B2(n_2731),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2879),
.Y(n_3065)
);

AOI22xp33_ASAP7_75t_L g3066 ( 
.A1(n_2892),
.A2(n_2776),
.B1(n_2752),
.B2(n_2777),
.Y(n_3066)
);

OAI22xp5_ASAP7_75t_L g3067 ( 
.A1(n_2861),
.A2(n_2776),
.B1(n_2685),
.B2(n_2697),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2863),
.Y(n_3068)
);

OAI22xp5_ASAP7_75t_L g3069 ( 
.A1(n_2861),
.A2(n_2685),
.B1(n_2782),
.B2(n_2597),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2863),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2815),
.Y(n_3071)
);

HB1xp67_ASAP7_75t_L g3072 ( 
.A(n_2954),
.Y(n_3072)
);

AOI22xp33_ASAP7_75t_SL g3073 ( 
.A1(n_3001),
.A2(n_2910),
.B1(n_2844),
.B2(n_2859),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2816),
.Y(n_3074)
);

CKINVDCx16_ASAP7_75t_R g3075 ( 
.A(n_2804),
.Y(n_3075)
);

BUFx2_ASAP7_75t_L g3076 ( 
.A(n_2950),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2887),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2825),
.Y(n_3078)
);

OAI22xp33_ASAP7_75t_L g3079 ( 
.A1(n_2928),
.A2(n_2778),
.B1(n_2676),
.B2(n_2659),
.Y(n_3079)
);

AND2x2_ASAP7_75t_L g3080 ( 
.A(n_2950),
.B(n_2630),
.Y(n_3080)
);

BUFx2_ASAP7_75t_R g3081 ( 
.A(n_2864),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2828),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2887),
.Y(n_3083)
);

BUFx12f_ASAP7_75t_L g3084 ( 
.A(n_2830),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2899),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2899),
.Y(n_3086)
);

INVx3_ASAP7_75t_L g3087 ( 
.A(n_2827),
.Y(n_3087)
);

AOI22xp5_ASAP7_75t_L g3088 ( 
.A1(n_2919),
.A2(n_2638),
.B1(n_2779),
.B2(n_2616),
.Y(n_3088)
);

AO21x1_ASAP7_75t_L g3089 ( 
.A1(n_3011),
.A2(n_2787),
.B(n_2755),
.Y(n_3089)
);

BUFx6f_ASAP7_75t_L g3090 ( 
.A(n_2854),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2904),
.Y(n_3091)
);

CKINVDCx5p33_ASAP7_75t_R g3092 ( 
.A(n_2974),
.Y(n_3092)
);

BUFx6f_ASAP7_75t_L g3093 ( 
.A(n_2854),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2904),
.Y(n_3094)
);

AOI21x1_ASAP7_75t_L g3095 ( 
.A1(n_3014),
.A2(n_2676),
.B(n_2658),
.Y(n_3095)
);

INVx3_ASAP7_75t_L g3096 ( 
.A(n_2827),
.Y(n_3096)
);

BUFx6f_ASAP7_75t_L g3097 ( 
.A(n_2854),
.Y(n_3097)
);

INVx2_ASAP7_75t_L g3098 ( 
.A(n_2875),
.Y(n_3098)
);

AOI22xp33_ASAP7_75t_SL g3099 ( 
.A1(n_2996),
.A2(n_2639),
.B1(n_2597),
.B2(n_2762),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2836),
.Y(n_3100)
);

OAI22xp33_ASAP7_75t_L g3101 ( 
.A1(n_2889),
.A2(n_2737),
.B1(n_2744),
.B2(n_2795),
.Y(n_3101)
);

CKINVDCx11_ASAP7_75t_R g3102 ( 
.A(n_2894),
.Y(n_3102)
);

CKINVDCx14_ASAP7_75t_R g3103 ( 
.A(n_3015),
.Y(n_3103)
);

AOI22xp33_ASAP7_75t_SL g3104 ( 
.A1(n_2952),
.A2(n_2639),
.B1(n_2764),
.B2(n_2624),
.Y(n_3104)
);

OAI22xp5_ASAP7_75t_L g3105 ( 
.A1(n_2866),
.A2(n_2799),
.B1(n_2687),
.B2(n_2596),
.Y(n_3105)
);

AND2x2_ASAP7_75t_L g3106 ( 
.A(n_2818),
.B(n_2799),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2840),
.Y(n_3107)
);

HB1xp67_ASAP7_75t_L g3108 ( 
.A(n_2954),
.Y(n_3108)
);

AND2x2_ASAP7_75t_L g3109 ( 
.A(n_2931),
.B(n_2612),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2846),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2885),
.Y(n_3111)
);

AOI22xp33_ASAP7_75t_L g3112 ( 
.A1(n_2972),
.A2(n_2563),
.B1(n_2551),
.B2(n_2768),
.Y(n_3112)
);

INVx1_ASAP7_75t_SL g3113 ( 
.A(n_2923),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2957),
.B(n_2565),
.Y(n_3114)
);

AOI22xp33_ASAP7_75t_SL g3115 ( 
.A1(n_2883),
.A2(n_2787),
.B1(n_2755),
.B2(n_2563),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2875),
.Y(n_3116)
);

AOI22xp33_ASAP7_75t_L g3117 ( 
.A1(n_2913),
.A2(n_2569),
.B1(n_2588),
.B2(n_2578),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2869),
.Y(n_3118)
);

BUFx6f_ASAP7_75t_L g3119 ( 
.A(n_2854),
.Y(n_3119)
);

BUFx2_ASAP7_75t_R g3120 ( 
.A(n_2962),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2827),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2874),
.Y(n_3122)
);

OAI21x1_ASAP7_75t_L g3123 ( 
.A1(n_2855),
.A2(n_2574),
.B(n_2578),
.Y(n_3123)
);

BUFx2_ASAP7_75t_R g3124 ( 
.A(n_2962),
.Y(n_3124)
);

INVx1_ASAP7_75t_SL g3125 ( 
.A(n_2835),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2917),
.Y(n_3126)
);

INVxp67_ASAP7_75t_L g3127 ( 
.A(n_2805),
.Y(n_3127)
);

AOI22xp33_ASAP7_75t_L g3128 ( 
.A1(n_2985),
.A2(n_2628),
.B1(n_2760),
.B2(n_2574),
.Y(n_3128)
);

BUFx4_ASAP7_75t_R g3129 ( 
.A(n_2821),
.Y(n_3129)
);

AND2x2_ASAP7_75t_L g3130 ( 
.A(n_2931),
.B(n_2783),
.Y(n_3130)
);

INVx3_ASAP7_75t_L g3131 ( 
.A(n_2806),
.Y(n_3131)
);

HB1xp67_ASAP7_75t_L g3132 ( 
.A(n_3010),
.Y(n_3132)
);

AO21x1_ASAP7_75t_L g3133 ( 
.A1(n_2989),
.A2(n_2787),
.B(n_2755),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2917),
.Y(n_3134)
);

OA21x2_ASAP7_75t_L g3135 ( 
.A1(n_2997),
.A2(n_2750),
.B(n_2656),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2918),
.Y(n_3136)
);

AOI22xp33_ASAP7_75t_L g3137 ( 
.A1(n_3002),
.A2(n_2760),
.B1(n_2628),
.B2(n_2750),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_2918),
.Y(n_3138)
);

INVxp67_ASAP7_75t_SL g3139 ( 
.A(n_2953),
.Y(n_3139)
);

OR2x2_ASAP7_75t_L g3140 ( 
.A(n_2961),
.B(n_2617),
.Y(n_3140)
);

AOI22xp33_ASAP7_75t_SL g3141 ( 
.A1(n_2945),
.A2(n_2750),
.B1(n_2631),
.B2(n_2619),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2933),
.Y(n_3142)
);

OR2x2_ASAP7_75t_L g3143 ( 
.A(n_2976),
.B(n_2617),
.Y(n_3143)
);

OR2x6_ASAP7_75t_L g3144 ( 
.A(n_2833),
.B(n_2800),
.Y(n_3144)
);

AOI21x1_ASAP7_75t_L g3145 ( 
.A1(n_2822),
.A2(n_2710),
.B(n_2617),
.Y(n_3145)
);

AO21x1_ASAP7_75t_L g3146 ( 
.A1(n_2980),
.A2(n_2610),
.B(n_2710),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2933),
.Y(n_3147)
);

CKINVDCx11_ASAP7_75t_R g3148 ( 
.A(n_2898),
.Y(n_3148)
);

AOI22xp33_ASAP7_75t_SL g3149 ( 
.A1(n_2945),
.A2(n_2800),
.B1(n_2667),
.B2(n_2710),
.Y(n_3149)
);

AOI22xp33_ASAP7_75t_L g3150 ( 
.A1(n_2946),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_3150)
);

OAI21x1_ASAP7_75t_L g3151 ( 
.A1(n_2838),
.A2(n_2983),
.B(n_2849),
.Y(n_3151)
);

AOI21x1_ASAP7_75t_L g3152 ( 
.A1(n_2945),
.A2(n_2667),
.B(n_234),
.Y(n_3152)
);

OAI21xp5_ASAP7_75t_SL g3153 ( 
.A1(n_2994),
.A2(n_2901),
.B(n_2890),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2930),
.Y(n_3154)
);

AOI22xp33_ASAP7_75t_SL g3155 ( 
.A1(n_2993),
.A2(n_2667),
.B1(n_235),
.B2(n_236),
.Y(n_3155)
);

BUFx8_ASAP7_75t_L g3156 ( 
.A(n_2902),
.Y(n_3156)
);

AND2x4_ASAP7_75t_L g3157 ( 
.A(n_2940),
.B(n_234),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2937),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_2810),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2992),
.B(n_235),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2810),
.Y(n_3161)
);

OA21x2_ASAP7_75t_L g3162 ( 
.A1(n_2997),
.A2(n_237),
.B(n_238),
.Y(n_3162)
);

AOI22xp33_ASAP7_75t_L g3163 ( 
.A1(n_3000),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2915),
.Y(n_3164)
);

CKINVDCx6p67_ASAP7_75t_R g3165 ( 
.A(n_2902),
.Y(n_3165)
);

AND2x2_ASAP7_75t_L g3166 ( 
.A(n_2831),
.B(n_239),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2937),
.Y(n_3167)
);

AOI21x1_ASAP7_75t_L g3168 ( 
.A1(n_2955),
.A2(n_241),
.B(n_242),
.Y(n_3168)
);

HB1xp67_ASAP7_75t_SL g3169 ( 
.A(n_2925),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_3008),
.Y(n_3170)
);

AND2x2_ASAP7_75t_L g3171 ( 
.A(n_2831),
.B(n_241),
.Y(n_3171)
);

AND2x4_ASAP7_75t_L g3172 ( 
.A(n_2940),
.B(n_242),
.Y(n_3172)
);

OAI22xp5_ASAP7_75t_L g3173 ( 
.A1(n_2866),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_2968),
.Y(n_3174)
);

AO21x1_ASAP7_75t_L g3175 ( 
.A1(n_2955),
.A2(n_244),
.B(n_246),
.Y(n_3175)
);

INVxp67_ASAP7_75t_L g3176 ( 
.A(n_2979),
.Y(n_3176)
);

BUFx4f_ASAP7_75t_SL g3177 ( 
.A(n_2925),
.Y(n_3177)
);

AOI22xp33_ASAP7_75t_L g3178 ( 
.A1(n_2867),
.A2(n_3003),
.B1(n_2907),
.B2(n_2803),
.Y(n_3178)
);

OAI21x1_ASAP7_75t_L g3179 ( 
.A1(n_2838),
.A2(n_246),
.B(n_247),
.Y(n_3179)
);

INVx3_ASAP7_75t_L g3180 ( 
.A(n_2806),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_3017),
.Y(n_3181)
);

INVx2_ASAP7_75t_SL g3182 ( 
.A(n_2831),
.Y(n_3182)
);

HB1xp67_ASAP7_75t_L g3183 ( 
.A(n_2935),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2966),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2939),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2941),
.Y(n_3186)
);

OAI22xp33_ASAP7_75t_L g3187 ( 
.A1(n_2833),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2971),
.Y(n_3188)
);

AOI21x1_ASAP7_75t_L g3189 ( 
.A1(n_2951),
.A2(n_250),
.B(n_251),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2971),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2968),
.Y(n_3191)
);

OAI22xp33_ASAP7_75t_L g3192 ( 
.A1(n_2833),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_3192)
);

INVx2_ASAP7_75t_SL g3193 ( 
.A(n_2940),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2927),
.Y(n_3194)
);

BUFx2_ASAP7_75t_R g3195 ( 
.A(n_3018),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2927),
.Y(n_3196)
);

INVx3_ASAP7_75t_L g3197 ( 
.A(n_2806),
.Y(n_3197)
);

AOI22xp33_ASAP7_75t_L g3198 ( 
.A1(n_3003),
.A2(n_252),
.B1(n_255),
.B2(n_256),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2927),
.Y(n_3199)
);

OA21x2_ASAP7_75t_L g3200 ( 
.A1(n_3005),
.A2(n_256),
.B(n_257),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2935),
.Y(n_3201)
);

BUFx12f_ASAP7_75t_L g3202 ( 
.A(n_2878),
.Y(n_3202)
);

INVx2_ASAP7_75t_L g3203 ( 
.A(n_2984),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_3005),
.Y(n_3204)
);

OA21x2_ASAP7_75t_L g3205 ( 
.A1(n_3019),
.A2(n_258),
.B(n_261),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_2984),
.Y(n_3206)
);

BUFx2_ASAP7_75t_L g3207 ( 
.A(n_2897),
.Y(n_3207)
);

AOI22xp33_ASAP7_75t_L g3208 ( 
.A1(n_2998),
.A2(n_258),
.B1(n_261),
.B2(n_262),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_3009),
.B(n_262),
.Y(n_3209)
);

INVx1_ASAP7_75t_SL g3210 ( 
.A(n_2835),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_3019),
.Y(n_3211)
);

INVx1_ASAP7_75t_SL g3212 ( 
.A(n_2835),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3025),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3025),
.Y(n_3214)
);

AOI22xp33_ASAP7_75t_L g3215 ( 
.A1(n_2998),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_3215)
);

INVx2_ASAP7_75t_L g3216 ( 
.A(n_2999),
.Y(n_3216)
);

AND2x2_ASAP7_75t_L g3217 ( 
.A(n_3022),
.B(n_264),
.Y(n_3217)
);

AO21x1_ASAP7_75t_L g3218 ( 
.A1(n_2929),
.A2(n_265),
.B(n_266),
.Y(n_3218)
);

NAND2x1p5_ASAP7_75t_L g3219 ( 
.A(n_2829),
.B(n_2853),
.Y(n_3219)
);

INVx3_ASAP7_75t_L g3220 ( 
.A(n_2853),
.Y(n_3220)
);

AOI22xp33_ASAP7_75t_L g3221 ( 
.A1(n_3073),
.A2(n_2833),
.B1(n_2998),
.B2(n_2809),
.Y(n_3221)
);

AOI22xp33_ASAP7_75t_L g3222 ( 
.A1(n_3050),
.A2(n_2809),
.B1(n_2942),
.B2(n_2924),
.Y(n_3222)
);

AOI22xp33_ASAP7_75t_SL g3223 ( 
.A1(n_3103),
.A2(n_2929),
.B1(n_2951),
.B2(n_2943),
.Y(n_3223)
);

BUFx2_ASAP7_75t_L g3224 ( 
.A(n_3131),
.Y(n_3224)
);

AOI22xp33_ASAP7_75t_L g3225 ( 
.A1(n_3050),
.A2(n_2809),
.B1(n_2942),
.B2(n_2924),
.Y(n_3225)
);

OAI222xp33_ASAP7_75t_L g3226 ( 
.A1(n_3052),
.A2(n_2878),
.B1(n_2832),
.B2(n_3013),
.C1(n_2942),
.C2(n_2947),
.Y(n_3226)
);

AOI22xp33_ASAP7_75t_SL g3227 ( 
.A1(n_3103),
.A2(n_2943),
.B1(n_2987),
.B2(n_2973),
.Y(n_3227)
);

AOI22xp33_ASAP7_75t_L g3228 ( 
.A1(n_3046),
.A2(n_2924),
.B1(n_2947),
.B2(n_2832),
.Y(n_3228)
);

AOI22xp33_ASAP7_75t_L g3229 ( 
.A1(n_3133),
.A2(n_2947),
.B1(n_2832),
.B2(n_2843),
.Y(n_3229)
);

AOI222xp33_ASAP7_75t_L g3230 ( 
.A1(n_3153),
.A2(n_3027),
.B1(n_3173),
.B2(n_3052),
.C1(n_3067),
.C2(n_3064),
.Y(n_3230)
);

AOI22xp33_ASAP7_75t_SL g3231 ( 
.A1(n_3105),
.A2(n_2943),
.B1(n_2987),
.B2(n_2973),
.Y(n_3231)
);

OAI22xp5_ASAP7_75t_L g3232 ( 
.A1(n_3027),
.A2(n_2965),
.B1(n_2890),
.B2(n_2852),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_3113),
.B(n_2896),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_3139),
.B(n_2916),
.Y(n_3234)
);

OAI21xp33_ASAP7_75t_L g3235 ( 
.A1(n_3208),
.A2(n_2965),
.B(n_3023),
.Y(n_3235)
);

INVx5_ASAP7_75t_SL g3236 ( 
.A(n_3144),
.Y(n_3236)
);

OR2x2_ASAP7_75t_L g3237 ( 
.A(n_3183),
.B(n_2999),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_3031),
.Y(n_3238)
);

AOI22xp33_ASAP7_75t_L g3239 ( 
.A1(n_3054),
.A2(n_2832),
.B1(n_2843),
.B2(n_2817),
.Y(n_3239)
);

INVx3_ASAP7_75t_L g3240 ( 
.A(n_3029),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_3030),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_3034),
.Y(n_3242)
);

AOI22xp33_ASAP7_75t_L g3243 ( 
.A1(n_3175),
.A2(n_2843),
.B1(n_2817),
.B2(n_2845),
.Y(n_3243)
);

OAI22xp5_ASAP7_75t_L g3244 ( 
.A1(n_3137),
.A2(n_3013),
.B1(n_2948),
.B2(n_2981),
.Y(n_3244)
);

AOI22xp33_ASAP7_75t_L g3245 ( 
.A1(n_3089),
.A2(n_2817),
.B1(n_2978),
.B2(n_2973),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_3059),
.B(n_3004),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3031),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_3036),
.Y(n_3248)
);

AOI22xp33_ASAP7_75t_L g3249 ( 
.A1(n_3115),
.A2(n_2873),
.B1(n_2802),
.B2(n_2823),
.Y(n_3249)
);

AOI22xp33_ASAP7_75t_L g3250 ( 
.A1(n_3208),
.A2(n_2873),
.B1(n_2802),
.B2(n_2823),
.Y(n_3250)
);

OAI22xp5_ASAP7_75t_SL g3251 ( 
.A1(n_3075),
.A2(n_2960),
.B1(n_2987),
.B2(n_2981),
.Y(n_3251)
);

NOR2xp33_ASAP7_75t_L g3252 ( 
.A(n_3176),
.B(n_3004),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3118),
.B(n_2990),
.Y(n_3253)
);

CKINVDCx11_ASAP7_75t_R g3254 ( 
.A(n_3084),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3043),
.Y(n_3255)
);

HB1xp67_ASAP7_75t_L g3256 ( 
.A(n_3132),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_3044),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_3122),
.B(n_2990),
.Y(n_3258)
);

AOI22xp33_ASAP7_75t_L g3259 ( 
.A1(n_3215),
.A2(n_2873),
.B1(n_2802),
.B2(n_2823),
.Y(n_3259)
);

NAND3xp33_ASAP7_75t_L g3260 ( 
.A(n_3053),
.B(n_2906),
.C(n_3006),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3045),
.Y(n_3261)
);

OAI22xp5_ASAP7_75t_L g3262 ( 
.A1(n_3137),
.A2(n_2948),
.B1(n_2981),
.B2(n_2963),
.Y(n_3262)
);

INVxp67_ASAP7_75t_L g3263 ( 
.A(n_3072),
.Y(n_3263)
);

OAI22x1_ASAP7_75t_L g3264 ( 
.A1(n_3076),
.A2(n_2988),
.B1(n_2963),
.B2(n_2829),
.Y(n_3264)
);

AND2x2_ASAP7_75t_L g3265 ( 
.A(n_3159),
.B(n_2808),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3083),
.Y(n_3266)
);

OAI22xp5_ASAP7_75t_L g3267 ( 
.A1(n_3215),
.A2(n_2948),
.B1(n_2988),
.B2(n_2963),
.Y(n_3267)
);

NOR2xp33_ASAP7_75t_L g3268 ( 
.A(n_3055),
.B(n_2988),
.Y(n_3268)
);

AOI22xp33_ASAP7_75t_SL g3269 ( 
.A1(n_3069),
.A2(n_3023),
.B1(n_3024),
.B2(n_2922),
.Y(n_3269)
);

AOI22xp33_ASAP7_75t_SL g3270 ( 
.A1(n_3202),
.A2(n_3039),
.B1(n_3156),
.B2(n_3053),
.Y(n_3270)
);

AOI22xp33_ASAP7_75t_L g3271 ( 
.A1(n_3202),
.A2(n_2922),
.B1(n_3024),
.B2(n_2824),
.Y(n_3271)
);

AOI22xp33_ASAP7_75t_L g3272 ( 
.A1(n_3104),
.A2(n_2922),
.B1(n_2824),
.B2(n_2891),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3036),
.Y(n_3273)
);

AOI22xp33_ASAP7_75t_L g3274 ( 
.A1(n_3099),
.A2(n_2891),
.B1(n_2814),
.B2(n_2956),
.Y(n_3274)
);

BUFx4f_ASAP7_75t_SL g3275 ( 
.A(n_3084),
.Y(n_3275)
);

OAI21xp5_ASAP7_75t_SL g3276 ( 
.A1(n_3088),
.A2(n_3198),
.B(n_3066),
.Y(n_3276)
);

AOI22xp33_ASAP7_75t_L g3277 ( 
.A1(n_3150),
.A2(n_2814),
.B1(n_2956),
.B2(n_2949),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_3042),
.B(n_2877),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_3040),
.Y(n_3279)
);

AOI22xp33_ASAP7_75t_L g3280 ( 
.A1(n_3150),
.A2(n_2949),
.B1(n_2938),
.B2(n_2895),
.Y(n_3280)
);

AOI22xp33_ASAP7_75t_L g3281 ( 
.A1(n_3163),
.A2(n_3155),
.B1(n_3218),
.B2(n_3066),
.Y(n_3281)
);

AOI22xp33_ASAP7_75t_L g3282 ( 
.A1(n_3163),
.A2(n_2938),
.B1(n_2895),
.B2(n_2964),
.Y(n_3282)
);

INVx3_ASAP7_75t_L g3283 ( 
.A(n_3029),
.Y(n_3283)
);

CKINVDCx5p33_ASAP7_75t_R g3284 ( 
.A(n_3033),
.Y(n_3284)
);

AOI22xp5_ASAP7_75t_L g3285 ( 
.A1(n_3187),
.A2(n_2835),
.B1(n_2850),
.B2(n_2877),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3085),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3108),
.B(n_2914),
.Y(n_3287)
);

AND2x2_ASAP7_75t_L g3288 ( 
.A(n_3161),
.B(n_2808),
.Y(n_3288)
);

AOI22xp33_ASAP7_75t_SL g3289 ( 
.A1(n_3039),
.A2(n_2964),
.B1(n_2886),
.B2(n_3020),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_3040),
.Y(n_3290)
);

AOI22xp33_ASAP7_75t_SL g3291 ( 
.A1(n_3039),
.A2(n_2886),
.B1(n_3021),
.B2(n_3020),
.Y(n_3291)
);

AND2x2_ASAP7_75t_L g3292 ( 
.A(n_3201),
.B(n_2897),
.Y(n_3292)
);

AOI22xp33_ASAP7_75t_L g3293 ( 
.A1(n_3198),
.A2(n_3178),
.B1(n_3112),
.B2(n_3192),
.Y(n_3293)
);

AOI22xp33_ASAP7_75t_L g3294 ( 
.A1(n_3178),
.A2(n_2819),
.B1(n_2820),
.B2(n_3021),
.Y(n_3294)
);

OAI22xp5_ASAP7_75t_L g3295 ( 
.A1(n_3128),
.A2(n_2850),
.B1(n_2898),
.B2(n_2908),
.Y(n_3295)
);

OAI222xp33_ASAP7_75t_L g3296 ( 
.A1(n_3038),
.A2(n_2886),
.B1(n_2991),
.B2(n_2914),
.C1(n_3006),
.C2(n_2921),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_3051),
.Y(n_3297)
);

OAI22xp5_ASAP7_75t_L g3298 ( 
.A1(n_3128),
.A2(n_3112),
.B1(n_3117),
.B2(n_3141),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_3170),
.B(n_2914),
.Y(n_3299)
);

OAI21xp5_ASAP7_75t_SL g3300 ( 
.A1(n_3079),
.A2(n_2886),
.B(n_2991),
.Y(n_3300)
);

AOI22xp33_ASAP7_75t_SL g3301 ( 
.A1(n_3156),
.A2(n_2886),
.B1(n_2986),
.B2(n_2882),
.Y(n_3301)
);

AOI22xp33_ASAP7_75t_SL g3302 ( 
.A1(n_3156),
.A2(n_2986),
.B1(n_2882),
.B2(n_2920),
.Y(n_3302)
);

AOI22xp33_ASAP7_75t_SL g3303 ( 
.A1(n_3053),
.A2(n_2920),
.B1(n_2850),
.B2(n_2977),
.Y(n_3303)
);

AOI22xp5_ASAP7_75t_L g3304 ( 
.A1(n_3101),
.A2(n_2850),
.B1(n_2925),
.B2(n_2820),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_3026),
.B(n_2908),
.Y(n_3305)
);

OAI21xp33_ASAP7_75t_L g3306 ( 
.A1(n_3168),
.A2(n_2982),
.B(n_2977),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_SL g3307 ( 
.A(n_3114),
.B(n_2898),
.Y(n_3307)
);

AOI22xp33_ASAP7_75t_SL g3308 ( 
.A1(n_3200),
.A2(n_2982),
.B1(n_2936),
.B2(n_2934),
.Y(n_3308)
);

AOI22xp33_ASAP7_75t_SL g3309 ( 
.A1(n_3200),
.A2(n_2936),
.B1(n_2934),
.B2(n_2905),
.Y(n_3309)
);

OR2x2_ASAP7_75t_L g3310 ( 
.A(n_3194),
.B(n_2983),
.Y(n_3310)
);

AND2x2_ASAP7_75t_L g3311 ( 
.A(n_3182),
.B(n_2944),
.Y(n_3311)
);

AOI22xp33_ASAP7_75t_L g3312 ( 
.A1(n_3117),
.A2(n_2819),
.B1(n_2820),
.B2(n_2921),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3091),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_3051),
.Y(n_3314)
);

AOI22xp33_ASAP7_75t_L g3315 ( 
.A1(n_3165),
.A2(n_2819),
.B1(n_2921),
.B2(n_2905),
.Y(n_3315)
);

OAI22xp5_ASAP7_75t_L g3316 ( 
.A1(n_3169),
.A2(n_2898),
.B1(n_2944),
.B2(n_2967),
.Y(n_3316)
);

OAI22xp5_ASAP7_75t_L g3317 ( 
.A1(n_3165),
.A2(n_2967),
.B1(n_2970),
.B2(n_2995),
.Y(n_3317)
);

HB1xp67_ASAP7_75t_L g3318 ( 
.A(n_3121),
.Y(n_3318)
);

INVx5_ASAP7_75t_SL g3319 ( 
.A(n_3144),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_3065),
.Y(n_3320)
);

AND2x2_ASAP7_75t_L g3321 ( 
.A(n_3182),
.B(n_2970),
.Y(n_3321)
);

BUFx3_ASAP7_75t_L g3322 ( 
.A(n_3207),
.Y(n_3322)
);

INVx2_ASAP7_75t_SL g3323 ( 
.A(n_3035),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3065),
.Y(n_3324)
);

INVx2_ASAP7_75t_L g3325 ( 
.A(n_3077),
.Y(n_3325)
);

OAI22xp5_ASAP7_75t_L g3326 ( 
.A1(n_3177),
.A2(n_3127),
.B1(n_3124),
.B2(n_3120),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_3077),
.Y(n_3327)
);

AOI22xp33_ASAP7_75t_L g3328 ( 
.A1(n_3157),
.A2(n_2921),
.B1(n_3016),
.B2(n_3007),
.Y(n_3328)
);

AOI22xp33_ASAP7_75t_SL g3329 ( 
.A1(n_3200),
.A2(n_3205),
.B1(n_3162),
.B2(n_3033),
.Y(n_3329)
);

AOI22xp33_ASAP7_75t_L g3330 ( 
.A1(n_3157),
.A2(n_3016),
.B1(n_3007),
.B2(n_2856),
.Y(n_3330)
);

AOI22xp33_ASAP7_75t_L g3331 ( 
.A1(n_3157),
.A2(n_2856),
.B1(n_2926),
.B2(n_2932),
.Y(n_3331)
);

AOI22xp33_ASAP7_75t_L g3332 ( 
.A1(n_3172),
.A2(n_2926),
.B1(n_2932),
.B2(n_2880),
.Y(n_3332)
);

HB1xp67_ASAP7_75t_L g3333 ( 
.A(n_3121),
.Y(n_3333)
);

AOI22xp5_ASAP7_75t_L g3334 ( 
.A1(n_3172),
.A2(n_2880),
.B1(n_2884),
.B2(n_2865),
.Y(n_3334)
);

AOI22xp33_ASAP7_75t_L g3335 ( 
.A1(n_3172),
.A2(n_2884),
.B1(n_2995),
.B2(n_3012),
.Y(n_3335)
);

AOI22xp33_ASAP7_75t_L g3336 ( 
.A1(n_3146),
.A2(n_3032),
.B1(n_3056),
.B2(n_3080),
.Y(n_3336)
);

AND2x2_ASAP7_75t_L g3337 ( 
.A(n_3068),
.B(n_2995),
.Y(n_3337)
);

INVx2_ASAP7_75t_SL g3338 ( 
.A(n_3035),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3094),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3086),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_3086),
.Y(n_3341)
);

NOR2xp33_ASAP7_75t_L g3342 ( 
.A(n_3055),
.B(n_2995),
.Y(n_3342)
);

HB1xp67_ASAP7_75t_L g3343 ( 
.A(n_3188),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3058),
.Y(n_3344)
);

AOI22xp33_ASAP7_75t_SL g3345 ( 
.A1(n_3205),
.A2(n_2991),
.B1(n_2871),
.B2(n_2888),
.Y(n_3345)
);

AOI22xp33_ASAP7_75t_SL g3346 ( 
.A1(n_3205),
.A2(n_2991),
.B1(n_2871),
.B2(n_2888),
.Y(n_3346)
);

OAI22xp5_ASAP7_75t_L g3347 ( 
.A1(n_3177),
.A2(n_3012),
.B1(n_2995),
.B2(n_2991),
.Y(n_3347)
);

OAI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_3037),
.A2(n_2893),
.B(n_2911),
.Y(n_3348)
);

AOI22xp33_ASAP7_75t_L g3349 ( 
.A1(n_3057),
.A2(n_3012),
.B1(n_2865),
.B2(n_2860),
.Y(n_3349)
);

AOI22xp33_ASAP7_75t_L g3350 ( 
.A1(n_3166),
.A2(n_3012),
.B1(n_2860),
.B2(n_2857),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_3098),
.Y(n_3351)
);

INVx2_ASAP7_75t_L g3352 ( 
.A(n_3098),
.Y(n_3352)
);

OAI21xp5_ASAP7_75t_SL g3353 ( 
.A1(n_3189),
.A2(n_2914),
.B(n_3012),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_3181),
.B(n_3185),
.Y(n_3354)
);

OAI21xp33_ASAP7_75t_L g3355 ( 
.A1(n_3196),
.A2(n_3199),
.B(n_3047),
.Y(n_3355)
);

INVx2_ASAP7_75t_L g3356 ( 
.A(n_3116),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3116),
.Y(n_3357)
);

OAI22xp5_ASAP7_75t_L g3358 ( 
.A1(n_3060),
.A2(n_2914),
.B1(n_2826),
.B2(n_2839),
.Y(n_3358)
);

AOI22xp33_ASAP7_75t_L g3359 ( 
.A1(n_3171),
.A2(n_2857),
.B1(n_2893),
.B2(n_2839),
.Y(n_3359)
);

BUFx2_ASAP7_75t_L g3360 ( 
.A(n_3131),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3061),
.Y(n_3361)
);

INVx2_ASAP7_75t_L g3362 ( 
.A(n_3126),
.Y(n_3362)
);

AND2x4_ASAP7_75t_L g3363 ( 
.A(n_3144),
.B(n_2841),
.Y(n_3363)
);

INVxp67_ASAP7_75t_L g3364 ( 
.A(n_3164),
.Y(n_3364)
);

AND2x2_ASAP7_75t_L g3365 ( 
.A(n_3070),
.B(n_2841),
.Y(n_3365)
);

AOI222xp33_ASAP7_75t_L g3366 ( 
.A1(n_3217),
.A2(n_2912),
.B1(n_2911),
.B2(n_268),
.C1(n_270),
.C2(n_271),
.Y(n_3366)
);

BUFx2_ASAP7_75t_L g3367 ( 
.A(n_3131),
.Y(n_3367)
);

BUFx4f_ASAP7_75t_SL g3368 ( 
.A(n_3060),
.Y(n_3368)
);

BUFx12f_ASAP7_75t_L g3369 ( 
.A(n_3028),
.Y(n_3369)
);

AOI22xp33_ASAP7_75t_L g3370 ( 
.A1(n_3144),
.A2(n_2969),
.B1(n_2912),
.B2(n_2848),
.Y(n_3370)
);

AOI22xp33_ASAP7_75t_L g3371 ( 
.A1(n_3162),
.A2(n_2969),
.B1(n_2848),
.B2(n_2849),
.Y(n_3371)
);

BUFx2_ASAP7_75t_L g3372 ( 
.A(n_3180),
.Y(n_3372)
);

CKINVDCx5p33_ASAP7_75t_R g3373 ( 
.A(n_3028),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_3126),
.Y(n_3374)
);

OAI21xp33_ASAP7_75t_L g3375 ( 
.A1(n_3037),
.A2(n_266),
.B(n_267),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3186),
.B(n_2826),
.Y(n_3376)
);

OAI22xp33_ASAP7_75t_L g3377 ( 
.A1(n_3063),
.A2(n_2826),
.B1(n_272),
.B2(n_273),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3136),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3154),
.B(n_2826),
.Y(n_3379)
);

BUFx4f_ASAP7_75t_SL g3380 ( 
.A(n_3125),
.Y(n_3380)
);

XOR2xp5_ASAP7_75t_L g3381 ( 
.A(n_3284),
.B(n_3092),
.Y(n_3381)
);

OR2x6_ASAP7_75t_L g3382 ( 
.A(n_3369),
.B(n_3041),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_3241),
.Y(n_3383)
);

NAND2xp33_ASAP7_75t_SL g3384 ( 
.A(n_3373),
.B(n_3092),
.Y(n_3384)
);

AND2x4_ASAP7_75t_L g3385 ( 
.A(n_3363),
.B(n_3190),
.Y(n_3385)
);

AND2x4_ASAP7_75t_L g3386 ( 
.A(n_3363),
.B(n_3109),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3256),
.B(n_3071),
.Y(n_3387)
);

NAND2xp33_ASAP7_75t_R g3388 ( 
.A(n_3373),
.B(n_3162),
.Y(n_3388)
);

NOR2xp33_ASAP7_75t_R g3389 ( 
.A(n_3254),
.B(n_3369),
.Y(n_3389)
);

NOR2xp33_ASAP7_75t_R g3390 ( 
.A(n_3254),
.B(n_3102),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3234),
.B(n_3074),
.Y(n_3391)
);

AND2x4_ASAP7_75t_L g3392 ( 
.A(n_3363),
.B(n_3193),
.Y(n_3392)
);

XNOR2xp5_ASAP7_75t_L g3393 ( 
.A(n_3284),
.B(n_3106),
.Y(n_3393)
);

INVxp67_ASAP7_75t_L g3394 ( 
.A(n_3252),
.Y(n_3394)
);

NAND2xp33_ASAP7_75t_R g3395 ( 
.A(n_3342),
.B(n_3209),
.Y(n_3395)
);

NAND2xp33_ASAP7_75t_R g3396 ( 
.A(n_3224),
.B(n_3081),
.Y(n_3396)
);

NAND2xp33_ASAP7_75t_R g3397 ( 
.A(n_3224),
.B(n_3180),
.Y(n_3397)
);

AND2x2_ASAP7_75t_L g3398 ( 
.A(n_3305),
.B(n_3130),
.Y(n_3398)
);

NAND2xp33_ASAP7_75t_R g3399 ( 
.A(n_3360),
.B(n_3180),
.Y(n_3399)
);

BUFx3_ASAP7_75t_L g3400 ( 
.A(n_3368),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3242),
.Y(n_3401)
);

NAND2xp33_ASAP7_75t_R g3402 ( 
.A(n_3360),
.B(n_3197),
.Y(n_3402)
);

OR2x6_ASAP7_75t_L g3403 ( 
.A(n_3316),
.B(n_3041),
.Y(n_3403)
);

AND2x4_ASAP7_75t_L g3404 ( 
.A(n_3323),
.B(n_3193),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3255),
.Y(n_3405)
);

AND2x4_ASAP7_75t_L g3406 ( 
.A(n_3323),
.B(n_3197),
.Y(n_3406)
);

AND2x4_ASAP7_75t_L g3407 ( 
.A(n_3338),
.B(n_3197),
.Y(n_3407)
);

NOR2xp33_ASAP7_75t_R g3408 ( 
.A(n_3275),
.B(n_3102),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_3257),
.Y(n_3409)
);

NAND2xp33_ASAP7_75t_R g3410 ( 
.A(n_3367),
.B(n_3129),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_3240),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3261),
.Y(n_3412)
);

NOR2xp33_ASAP7_75t_R g3413 ( 
.A(n_3380),
.B(n_3148),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_3240),
.Y(n_3414)
);

OR2x2_ASAP7_75t_L g3415 ( 
.A(n_3287),
.B(n_3047),
.Y(n_3415)
);

BUFx2_ASAP7_75t_L g3416 ( 
.A(n_3322),
.Y(n_3416)
);

NOR2xp33_ASAP7_75t_R g3417 ( 
.A(n_3268),
.B(n_3148),
.Y(n_3417)
);

AND2x2_ASAP7_75t_L g3418 ( 
.A(n_3305),
.B(n_3210),
.Y(n_3418)
);

NOR2xp33_ASAP7_75t_R g3419 ( 
.A(n_3281),
.B(n_3095),
.Y(n_3419)
);

NAND2xp33_ASAP7_75t_R g3420 ( 
.A(n_3367),
.B(n_3129),
.Y(n_3420)
);

NAND2xp33_ASAP7_75t_R g3421 ( 
.A(n_3372),
.B(n_3160),
.Y(n_3421)
);

AND2x4_ASAP7_75t_L g3422 ( 
.A(n_3338),
.B(n_3184),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_3336),
.B(n_3078),
.Y(n_3423)
);

NAND2xp33_ASAP7_75t_R g3424 ( 
.A(n_3372),
.B(n_3087),
.Y(n_3424)
);

AND2x4_ASAP7_75t_L g3425 ( 
.A(n_3365),
.B(n_3087),
.Y(n_3425)
);

CKINVDCx5p33_ASAP7_75t_R g3426 ( 
.A(n_3326),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_3263),
.B(n_3082),
.Y(n_3427)
);

NOR2xp33_ASAP7_75t_R g3428 ( 
.A(n_3228),
.B(n_3195),
.Y(n_3428)
);

XOR2xp5_ASAP7_75t_L g3429 ( 
.A(n_3298),
.B(n_3262),
.Y(n_3429)
);

CKINVDCx8_ASAP7_75t_R g3430 ( 
.A(n_3270),
.Y(n_3430)
);

AND2x4_ASAP7_75t_L g3431 ( 
.A(n_3365),
.B(n_3087),
.Y(n_3431)
);

AND2x2_ASAP7_75t_L g3432 ( 
.A(n_3322),
.B(n_3212),
.Y(n_3432)
);

OR2x2_ASAP7_75t_L g3433 ( 
.A(n_3246),
.B(n_3140),
.Y(n_3433)
);

AND2x2_ASAP7_75t_L g3434 ( 
.A(n_3311),
.B(n_3136),
.Y(n_3434)
);

NOR2xp33_ASAP7_75t_R g3435 ( 
.A(n_3293),
.B(n_3233),
.Y(n_3435)
);

NOR2xp33_ASAP7_75t_L g3436 ( 
.A(n_3278),
.B(n_3111),
.Y(n_3436)
);

AND2x4_ASAP7_75t_L g3437 ( 
.A(n_3307),
.B(n_3096),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3266),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_3240),
.Y(n_3439)
);

NOR2xp33_ASAP7_75t_R g3440 ( 
.A(n_3222),
.B(n_3090),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3364),
.B(n_3100),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_L g3442 ( 
.A(n_3300),
.B(n_3107),
.Y(n_3442)
);

NOR2xp33_ASAP7_75t_R g3443 ( 
.A(n_3225),
.B(n_3090),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3358),
.B(n_3110),
.Y(n_3444)
);

AND2x4_ASAP7_75t_L g3445 ( 
.A(n_3307),
.B(n_3096),
.Y(n_3445)
);

INVxp67_ASAP7_75t_L g3446 ( 
.A(n_3253),
.Y(n_3446)
);

NOR2xp33_ASAP7_75t_R g3447 ( 
.A(n_3258),
.B(n_3090),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_3311),
.B(n_3138),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_SL g3449 ( 
.A(n_3223),
.B(n_3090),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3286),
.Y(n_3450)
);

NAND2xp33_ASAP7_75t_R g3451 ( 
.A(n_3321),
.B(n_3096),
.Y(n_3451)
);

AND2x4_ASAP7_75t_L g3452 ( 
.A(n_3321),
.B(n_3029),
.Y(n_3452)
);

AND2x4_ASAP7_75t_L g3453 ( 
.A(n_3292),
.B(n_3048),
.Y(n_3453)
);

HB1xp67_ASAP7_75t_L g3454 ( 
.A(n_3343),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_3354),
.B(n_3344),
.Y(n_3455)
);

OR2x6_ASAP7_75t_L g3456 ( 
.A(n_3251),
.B(n_3179),
.Y(n_3456)
);

BUFx10_ASAP7_75t_L g3457 ( 
.A(n_3361),
.Y(n_3457)
);

AND2x4_ASAP7_75t_SL g3458 ( 
.A(n_3285),
.B(n_3093),
.Y(n_3458)
);

INVxp67_ASAP7_75t_L g3459 ( 
.A(n_3337),
.Y(n_3459)
);

XNOR2xp5_ASAP7_75t_L g3460 ( 
.A(n_3244),
.B(n_3232),
.Y(n_3460)
);

NOR2xp33_ASAP7_75t_R g3461 ( 
.A(n_3221),
.B(n_3093),
.Y(n_3461)
);

AND2x2_ASAP7_75t_L g3462 ( 
.A(n_3337),
.B(n_3138),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3245),
.B(n_3134),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3313),
.Y(n_3464)
);

AND2x2_ASAP7_75t_L g3465 ( 
.A(n_3292),
.B(n_3142),
.Y(n_3465)
);

AND2x2_ASAP7_75t_L g3466 ( 
.A(n_3236),
.B(n_3147),
.Y(n_3466)
);

BUFx10_ASAP7_75t_L g3467 ( 
.A(n_3339),
.Y(n_3467)
);

INVxp67_ASAP7_75t_L g3468 ( 
.A(n_3299),
.Y(n_3468)
);

NAND2xp33_ASAP7_75t_R g3469 ( 
.A(n_3310),
.B(n_3135),
.Y(n_3469)
);

NAND2xp33_ASAP7_75t_R g3470 ( 
.A(n_3310),
.B(n_3135),
.Y(n_3470)
);

AND2x2_ASAP7_75t_L g3471 ( 
.A(n_3236),
.B(n_3048),
.Y(n_3471)
);

NAND2xp33_ASAP7_75t_R g3472 ( 
.A(n_3376),
.B(n_3135),
.Y(n_3472)
);

CKINVDCx5p33_ASAP7_75t_R g3473 ( 
.A(n_3317),
.Y(n_3473)
);

NAND2xp33_ASAP7_75t_R g3474 ( 
.A(n_3379),
.B(n_3143),
.Y(n_3474)
);

AND2x2_ASAP7_75t_L g3475 ( 
.A(n_3236),
.B(n_3048),
.Y(n_3475)
);

INVxp67_ASAP7_75t_L g3476 ( 
.A(n_3318),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3353),
.B(n_3149),
.Y(n_3477)
);

NAND2xp33_ASAP7_75t_R g3478 ( 
.A(n_3283),
.B(n_3062),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_SL g3479 ( 
.A(n_3304),
.B(n_3093),
.Y(n_3479)
);

AND2x2_ASAP7_75t_L g3480 ( 
.A(n_3236),
.B(n_3319),
.Y(n_3480)
);

OR2x6_ASAP7_75t_L g3481 ( 
.A(n_3260),
.B(n_3179),
.Y(n_3481)
);

AND2x4_ASAP7_75t_L g3482 ( 
.A(n_3265),
.B(n_3062),
.Y(n_3482)
);

AND2x4_ASAP7_75t_L g3483 ( 
.A(n_3265),
.B(n_3062),
.Y(n_3483)
);

NAND2xp33_ASAP7_75t_R g3484 ( 
.A(n_3283),
.B(n_3220),
.Y(n_3484)
);

AND2x4_ASAP7_75t_L g3485 ( 
.A(n_3288),
.B(n_3220),
.Y(n_3485)
);

BUFx10_ASAP7_75t_L g3486 ( 
.A(n_3340),
.Y(n_3486)
);

NOR2xp67_ASAP7_75t_L g3487 ( 
.A(n_3264),
.B(n_3220),
.Y(n_3487)
);

AND2x4_ASAP7_75t_L g3488 ( 
.A(n_3288),
.B(n_3093),
.Y(n_3488)
);

AND2x2_ASAP7_75t_L g3489 ( 
.A(n_3319),
.B(n_3097),
.Y(n_3489)
);

INVxp67_ASAP7_75t_L g3490 ( 
.A(n_3333),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3247),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3247),
.Y(n_3492)
);

AND2x2_ASAP7_75t_L g3493 ( 
.A(n_3319),
.B(n_3097),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_SL g3494 ( 
.A(n_3230),
.B(n_3097),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3248),
.Y(n_3495)
);

INVx2_ASAP7_75t_L g3496 ( 
.A(n_3283),
.Y(n_3496)
);

NOR2xp33_ASAP7_75t_R g3497 ( 
.A(n_3229),
.B(n_3097),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3355),
.B(n_3119),
.Y(n_3498)
);

INVx2_ASAP7_75t_SL g3499 ( 
.A(n_3238),
.Y(n_3499)
);

INVxp67_ASAP7_75t_L g3500 ( 
.A(n_3264),
.Y(n_3500)
);

NOR2xp33_ASAP7_75t_R g3501 ( 
.A(n_3335),
.B(n_3119),
.Y(n_3501)
);

NAND2xp33_ASAP7_75t_R g3502 ( 
.A(n_3226),
.B(n_268),
.Y(n_3502)
);

INVx2_ASAP7_75t_L g3503 ( 
.A(n_3238),
.Y(n_3503)
);

AND2x4_ASAP7_75t_L g3504 ( 
.A(n_3334),
.B(n_3119),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3249),
.B(n_3119),
.Y(n_3505)
);

INVxp67_ASAP7_75t_L g3506 ( 
.A(n_3347),
.Y(n_3506)
);

NAND2xp33_ASAP7_75t_R g3507 ( 
.A(n_3357),
.B(n_272),
.Y(n_3507)
);

OR2x2_ASAP7_75t_L g3508 ( 
.A(n_3237),
.B(n_3219),
.Y(n_3508)
);

INVxp67_ASAP7_75t_L g3509 ( 
.A(n_3248),
.Y(n_3509)
);

OR2x6_ASAP7_75t_L g3510 ( 
.A(n_3295),
.B(n_3219),
.Y(n_3510)
);

AND2x2_ASAP7_75t_L g3511 ( 
.A(n_3319),
.B(n_3357),
.Y(n_3511)
);

BUFx3_ASAP7_75t_L g3512 ( 
.A(n_3351),
.Y(n_3512)
);

AND2x2_ASAP7_75t_L g3513 ( 
.A(n_3378),
.B(n_3049),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3383),
.Y(n_3514)
);

HB1xp67_ASAP7_75t_L g3515 ( 
.A(n_3454),
.Y(n_3515)
);

INVx2_ASAP7_75t_L g3516 ( 
.A(n_3512),
.Y(n_3516)
);

AND2x2_ASAP7_75t_L g3517 ( 
.A(n_3392),
.B(n_3403),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_3392),
.B(n_3329),
.Y(n_3518)
);

INVxp67_ASAP7_75t_L g3519 ( 
.A(n_3507),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_3467),
.Y(n_3520)
);

INVxp67_ASAP7_75t_L g3521 ( 
.A(n_3494),
.Y(n_3521)
);

INVxp67_ASAP7_75t_R g3522 ( 
.A(n_3480),
.Y(n_3522)
);

AND2x2_ASAP7_75t_L g3523 ( 
.A(n_3403),
.B(n_3279),
.Y(n_3523)
);

AND2x4_ASAP7_75t_L g3524 ( 
.A(n_3382),
.B(n_3348),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3401),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_3467),
.Y(n_3526)
);

OR2x2_ASAP7_75t_L g3527 ( 
.A(n_3442),
.B(n_3468),
.Y(n_3527)
);

BUFx3_ASAP7_75t_L g3528 ( 
.A(n_3416),
.Y(n_3528)
);

INVx2_ASAP7_75t_SL g3529 ( 
.A(n_3457),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3405),
.Y(n_3530)
);

OR2x2_ASAP7_75t_L g3531 ( 
.A(n_3463),
.B(n_3237),
.Y(n_3531)
);

AND2x2_ASAP7_75t_L g3532 ( 
.A(n_3386),
.B(n_3279),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3409),
.Y(n_3533)
);

AND2x4_ASAP7_75t_L g3534 ( 
.A(n_3382),
.B(n_3290),
.Y(n_3534)
);

AND2x2_ASAP7_75t_L g3535 ( 
.A(n_3386),
.B(n_3290),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3412),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3438),
.Y(n_3537)
);

NOR2xp33_ASAP7_75t_L g3538 ( 
.A(n_3426),
.B(n_3276),
.Y(n_3538)
);

INVx2_ASAP7_75t_L g3539 ( 
.A(n_3457),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3450),
.Y(n_3540)
);

NOR2xp33_ASAP7_75t_L g3541 ( 
.A(n_3384),
.B(n_3235),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3464),
.Y(n_3542)
);

AO21x2_ASAP7_75t_L g3543 ( 
.A1(n_3449),
.A2(n_3296),
.B(n_3377),
.Y(n_3543)
);

AOI22xp33_ASAP7_75t_L g3544 ( 
.A1(n_3429),
.A2(n_3239),
.B1(n_3375),
.B2(n_3269),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3441),
.Y(n_3545)
);

AND2x2_ASAP7_75t_L g3546 ( 
.A(n_3504),
.B(n_3297),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3491),
.Y(n_3547)
);

INVx2_ASAP7_75t_SL g3548 ( 
.A(n_3486),
.Y(n_3548)
);

INVx3_ASAP7_75t_L g3549 ( 
.A(n_3486),
.Y(n_3549)
);

HB1xp67_ASAP7_75t_L g3550 ( 
.A(n_3481),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3446),
.B(n_3291),
.Y(n_3551)
);

AND2x2_ASAP7_75t_L g3552 ( 
.A(n_3504),
.B(n_3297),
.Y(n_3552)
);

AND2x2_ASAP7_75t_L g3553 ( 
.A(n_3488),
.B(n_3314),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3436),
.B(n_3289),
.Y(n_3554)
);

INVx1_ASAP7_75t_SL g3555 ( 
.A(n_3390),
.Y(n_3555)
);

AND2x2_ASAP7_75t_L g3556 ( 
.A(n_3488),
.B(n_3500),
.Y(n_3556)
);

OA21x2_ASAP7_75t_L g3557 ( 
.A1(n_3477),
.A2(n_3151),
.B(n_3371),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3492),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3444),
.B(n_3394),
.Y(n_3559)
);

AND2x2_ASAP7_75t_L g3560 ( 
.A(n_3471),
.B(n_3314),
.Y(n_3560)
);

BUFx2_ASAP7_75t_L g3561 ( 
.A(n_3389),
.Y(n_3561)
);

AND2x2_ASAP7_75t_L g3562 ( 
.A(n_3475),
.B(n_3320),
.Y(n_3562)
);

AND2x4_ASAP7_75t_SL g3563 ( 
.A(n_3432),
.B(n_3330),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3391),
.B(n_3301),
.Y(n_3564)
);

INVxp67_ASAP7_75t_L g3565 ( 
.A(n_3421),
.Y(n_3565)
);

BUFx3_ASAP7_75t_L g3566 ( 
.A(n_3400),
.Y(n_3566)
);

AO21x2_ASAP7_75t_L g3567 ( 
.A1(n_3461),
.A2(n_3152),
.B(n_3306),
.Y(n_3567)
);

OAI322xp33_ASAP7_75t_L g3568 ( 
.A1(n_3502),
.A2(n_3267),
.A3(n_3273),
.B1(n_3324),
.B2(n_3378),
.C1(n_3341),
.C2(n_3325),
.Y(n_3568)
);

INVx3_ASAP7_75t_L g3569 ( 
.A(n_3406),
.Y(n_3569)
);

BUFx2_ASAP7_75t_L g3570 ( 
.A(n_3413),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3495),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3509),
.Y(n_3572)
);

INVx2_ASAP7_75t_L g3573 ( 
.A(n_3513),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_3503),
.Y(n_3574)
);

AND2x2_ASAP7_75t_L g3575 ( 
.A(n_3510),
.B(n_3320),
.Y(n_3575)
);

BUFx3_ASAP7_75t_L g3576 ( 
.A(n_3430),
.Y(n_3576)
);

AND2x2_ASAP7_75t_L g3577 ( 
.A(n_3510),
.B(n_3325),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_3499),
.Y(n_3578)
);

BUFx2_ASAP7_75t_L g3579 ( 
.A(n_3501),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3427),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3387),
.Y(n_3581)
);

OAI211xp5_ASAP7_75t_L g3582 ( 
.A1(n_3419),
.A2(n_3243),
.B(n_3231),
.C(n_3227),
.Y(n_3582)
);

AOI22xp33_ASAP7_75t_SL g3583 ( 
.A1(n_3497),
.A2(n_3366),
.B1(n_3049),
.B2(n_3259),
.Y(n_3583)
);

AND2x2_ASAP7_75t_L g3584 ( 
.A(n_3452),
.B(n_3327),
.Y(n_3584)
);

AOI21xp33_ASAP7_75t_SL g3585 ( 
.A1(n_3460),
.A2(n_3250),
.B(n_3272),
.Y(n_3585)
);

INVx2_ASAP7_75t_L g3586 ( 
.A(n_3411),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3423),
.B(n_3271),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3455),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_3414),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_3439),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3476),
.Y(n_3591)
);

OR2x2_ASAP7_75t_L g3592 ( 
.A(n_3415),
.B(n_3273),
.Y(n_3592)
);

OR2x2_ASAP7_75t_L g3593 ( 
.A(n_3481),
.B(n_3324),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3490),
.Y(n_3594)
);

OAI221xp5_ASAP7_75t_L g3595 ( 
.A1(n_3388),
.A2(n_3303),
.B1(n_3274),
.B2(n_3302),
.C(n_3294),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_3422),
.Y(n_3596)
);

INVx2_ASAP7_75t_L g3597 ( 
.A(n_3496),
.Y(n_3597)
);

INVx2_ASAP7_75t_L g3598 ( 
.A(n_3462),
.Y(n_3598)
);

AOI22xp5_ASAP7_75t_L g3599 ( 
.A1(n_3456),
.A2(n_3346),
.B1(n_3345),
.B2(n_3282),
.Y(n_3599)
);

INVx2_ASAP7_75t_L g3600 ( 
.A(n_3422),
.Y(n_3600)
);

BUFx2_ASAP7_75t_L g3601 ( 
.A(n_3447),
.Y(n_3601)
);

INVxp67_ASAP7_75t_SL g3602 ( 
.A(n_3487),
.Y(n_3602)
);

HB1xp67_ASAP7_75t_L g3603 ( 
.A(n_3459),
.Y(n_3603)
);

BUFx2_ASAP7_75t_L g3604 ( 
.A(n_3456),
.Y(n_3604)
);

AND2x2_ASAP7_75t_L g3605 ( 
.A(n_3452),
.B(n_3327),
.Y(n_3605)
);

AND2x2_ASAP7_75t_L g3606 ( 
.A(n_3511),
.B(n_3341),
.Y(n_3606)
);

HB1xp67_ASAP7_75t_L g3607 ( 
.A(n_3433),
.Y(n_3607)
);

OR2x2_ASAP7_75t_L g3608 ( 
.A(n_3506),
.B(n_3351),
.Y(n_3608)
);

AND2x2_ASAP7_75t_L g3609 ( 
.A(n_3453),
.B(n_3352),
.Y(n_3609)
);

INVx3_ASAP7_75t_L g3610 ( 
.A(n_3406),
.Y(n_3610)
);

HB1xp67_ASAP7_75t_L g3611 ( 
.A(n_3469),
.Y(n_3611)
);

NAND4xp25_ASAP7_75t_L g3612 ( 
.A(n_3505),
.B(n_3479),
.C(n_3395),
.D(n_3396),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3465),
.Y(n_3613)
);

BUFx2_ASAP7_75t_L g3614 ( 
.A(n_3408),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3434),
.Y(n_3615)
);

AND2x2_ASAP7_75t_L g3616 ( 
.A(n_3453),
.B(n_3352),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3448),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3385),
.B(n_3374),
.Y(n_3618)
);

NAND3xp33_ASAP7_75t_L g3619 ( 
.A(n_3472),
.B(n_3359),
.C(n_3277),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3498),
.Y(n_3620)
);

OR2x2_ASAP7_75t_L g3621 ( 
.A(n_3508),
.B(n_3356),
.Y(n_3621)
);

INVx2_ASAP7_75t_L g3622 ( 
.A(n_3425),
.Y(n_3622)
);

AO22x2_ASAP7_75t_L g3623 ( 
.A1(n_3385),
.A2(n_3374),
.B1(n_3362),
.B2(n_3356),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_L g3624 ( 
.A(n_3435),
.B(n_3350),
.Y(n_3624)
);

OAI221xp5_ASAP7_75t_L g3625 ( 
.A1(n_3410),
.A2(n_3420),
.B1(n_3474),
.B2(n_3473),
.C(n_3399),
.Y(n_3625)
);

AND2x2_ASAP7_75t_L g3626 ( 
.A(n_3425),
.B(n_3362),
.Y(n_3626)
);

AND2x2_ASAP7_75t_L g3627 ( 
.A(n_3431),
.B(n_3370),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3437),
.Y(n_3628)
);

NOR2x1_ASAP7_75t_L g3629 ( 
.A(n_3381),
.B(n_3204),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3458),
.B(n_3280),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_3466),
.B(n_3418),
.Y(n_3631)
);

INVx2_ASAP7_75t_L g3632 ( 
.A(n_3431),
.Y(n_3632)
);

HB1xp67_ASAP7_75t_L g3633 ( 
.A(n_3470),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3489),
.B(n_3308),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3437),
.Y(n_3635)
);

INVx1_ASAP7_75t_SL g3636 ( 
.A(n_3417),
.Y(n_3636)
);

AND2x2_ASAP7_75t_L g3637 ( 
.A(n_3493),
.B(n_3312),
.Y(n_3637)
);

INVx3_ASAP7_75t_L g3638 ( 
.A(n_3407),
.Y(n_3638)
);

OR2x2_ASAP7_75t_L g3639 ( 
.A(n_3485),
.B(n_3349),
.Y(n_3639)
);

OR2x2_ASAP7_75t_L g3640 ( 
.A(n_3485),
.B(n_3332),
.Y(n_3640)
);

AND2x2_ASAP7_75t_L g3641 ( 
.A(n_3522),
.B(n_3482),
.Y(n_3641)
);

INVx2_ASAP7_75t_L g3642 ( 
.A(n_3528),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3514),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3514),
.Y(n_3644)
);

AND2x4_ASAP7_75t_L g3645 ( 
.A(n_3556),
.B(n_3482),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_3521),
.B(n_3445),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_3519),
.B(n_3445),
.Y(n_3647)
);

AND2x2_ASAP7_75t_L g3648 ( 
.A(n_3522),
.B(n_3483),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_3528),
.Y(n_3649)
);

HB1xp67_ASAP7_75t_L g3650 ( 
.A(n_3515),
.Y(n_3650)
);

OR2x2_ASAP7_75t_L g3651 ( 
.A(n_3608),
.B(n_3483),
.Y(n_3651)
);

OR2x2_ASAP7_75t_L g3652 ( 
.A(n_3608),
.B(n_3398),
.Y(n_3652)
);

INVx2_ASAP7_75t_L g3653 ( 
.A(n_3623),
.Y(n_3653)
);

NOR2xp33_ASAP7_75t_L g3654 ( 
.A(n_3555),
.B(n_3393),
.Y(n_3654)
);

AND2x2_ASAP7_75t_L g3655 ( 
.A(n_3601),
.B(n_3407),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3547),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3601),
.B(n_3579),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3585),
.B(n_3440),
.Y(n_3658)
);

AND2x2_ASAP7_75t_L g3659 ( 
.A(n_3579),
.B(n_3404),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_3623),
.Y(n_3660)
);

OAI22xp5_ASAP7_75t_L g3661 ( 
.A1(n_3565),
.A2(n_3328),
.B1(n_3309),
.B2(n_3315),
.Y(n_3661)
);

AND2x4_ASAP7_75t_L g3662 ( 
.A(n_3556),
.B(n_3404),
.Y(n_3662)
);

AND2x2_ASAP7_75t_L g3663 ( 
.A(n_3602),
.B(n_3443),
.Y(n_3663)
);

INVx3_ASAP7_75t_L g3664 ( 
.A(n_3569),
.Y(n_3664)
);

NOR2xp33_ASAP7_75t_L g3665 ( 
.A(n_3561),
.B(n_273),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_SL g3666 ( 
.A(n_3629),
.B(n_3428),
.Y(n_3666)
);

NOR2xp33_ASAP7_75t_L g3667 ( 
.A(n_3561),
.B(n_3614),
.Y(n_3667)
);

OR2x2_ASAP7_75t_L g3668 ( 
.A(n_3527),
.B(n_3331),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3623),
.Y(n_3669)
);

BUFx3_ASAP7_75t_L g3670 ( 
.A(n_3614),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3547),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3558),
.Y(n_3672)
);

AND2x2_ASAP7_75t_L g3673 ( 
.A(n_3518),
.B(n_3604),
.Y(n_3673)
);

AND2x4_ASAP7_75t_L g3674 ( 
.A(n_3569),
.B(n_3174),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3558),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3571),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3544),
.B(n_3211),
.Y(n_3677)
);

AND2x4_ASAP7_75t_SL g3678 ( 
.A(n_3517),
.B(n_3397),
.Y(n_3678)
);

AND2x4_ASAP7_75t_SL g3679 ( 
.A(n_3517),
.B(n_3402),
.Y(n_3679)
);

AND2x2_ASAP7_75t_L g3680 ( 
.A(n_3518),
.B(n_3424),
.Y(n_3680)
);

INVx4_ASAP7_75t_R g3681 ( 
.A(n_3576),
.Y(n_3681)
);

HB1xp67_ASAP7_75t_L g3682 ( 
.A(n_3603),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3591),
.B(n_3213),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3571),
.Y(n_3684)
);

INVx2_ASAP7_75t_L g3685 ( 
.A(n_3623),
.Y(n_3685)
);

AND2x2_ASAP7_75t_L g3686 ( 
.A(n_3604),
.B(n_3569),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3591),
.B(n_3214),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3530),
.Y(n_3688)
);

AND2x4_ASAP7_75t_L g3689 ( 
.A(n_3610),
.B(n_3174),
.Y(n_3689)
);

HB1xp67_ASAP7_75t_L g3690 ( 
.A(n_3607),
.Y(n_3690)
);

AND2x2_ASAP7_75t_L g3691 ( 
.A(n_3610),
.B(n_3145),
.Y(n_3691)
);

AND2x2_ASAP7_75t_L g3692 ( 
.A(n_3610),
.B(n_3451),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3530),
.Y(n_3693)
);

BUFx6f_ASAP7_75t_L g3694 ( 
.A(n_3570),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3533),
.Y(n_3695)
);

AND2x2_ASAP7_75t_L g3696 ( 
.A(n_3638),
.B(n_3478),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3533),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3536),
.Y(n_3698)
);

INVxp67_ASAP7_75t_SL g3699 ( 
.A(n_3576),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3594),
.B(n_3191),
.Y(n_3700)
);

INVxp33_ASAP7_75t_L g3701 ( 
.A(n_3570),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3593),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3594),
.B(n_3191),
.Y(n_3703)
);

HB1xp67_ASAP7_75t_L g3704 ( 
.A(n_3578),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3536),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_3559),
.B(n_3203),
.Y(n_3706)
);

INVxp67_ASAP7_75t_SL g3707 ( 
.A(n_3611),
.Y(n_3707)
);

INVx3_ASAP7_75t_L g3708 ( 
.A(n_3638),
.Y(n_3708)
);

AND2x2_ASAP7_75t_L g3709 ( 
.A(n_3638),
.B(n_3203),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3540),
.Y(n_3710)
);

BUFx2_ASAP7_75t_L g3711 ( 
.A(n_3543),
.Y(n_3711)
);

AND2x2_ASAP7_75t_L g3712 ( 
.A(n_3634),
.B(n_3206),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3540),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3525),
.Y(n_3714)
);

INVx2_ASAP7_75t_L g3715 ( 
.A(n_3593),
.Y(n_3715)
);

AND2x2_ASAP7_75t_L g3716 ( 
.A(n_3634),
.B(n_3206),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3587),
.B(n_3216),
.Y(n_3717)
);

OR2x2_ASAP7_75t_L g3718 ( 
.A(n_3527),
.B(n_3216),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3637),
.B(n_3484),
.Y(n_3719)
);

INVx2_ASAP7_75t_L g3720 ( 
.A(n_3618),
.Y(n_3720)
);

INVxp67_ASAP7_75t_SL g3721 ( 
.A(n_3633),
.Y(n_3721)
);

BUFx6f_ASAP7_75t_L g3722 ( 
.A(n_3566),
.Y(n_3722)
);

AND2x6_ASAP7_75t_L g3723 ( 
.A(n_3636),
.B(n_3158),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3537),
.Y(n_3724)
);

AND2x4_ASAP7_75t_L g3725 ( 
.A(n_3600),
.B(n_3596),
.Y(n_3725)
);

OR2x2_ASAP7_75t_L g3726 ( 
.A(n_3531),
.B(n_3572),
.Y(n_3726)
);

OR2x2_ASAP7_75t_L g3727 ( 
.A(n_3531),
.B(n_3158),
.Y(n_3727)
);

AND2x4_ASAP7_75t_L g3728 ( 
.A(n_3600),
.B(n_3151),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3542),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3618),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_3626),
.Y(n_3731)
);

INVxp67_ASAP7_75t_L g3732 ( 
.A(n_3541),
.Y(n_3732)
);

HB1xp67_ASAP7_75t_L g3733 ( 
.A(n_3578),
.Y(n_3733)
);

INVx2_ASAP7_75t_L g3734 ( 
.A(n_3626),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3637),
.B(n_3167),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3580),
.B(n_3167),
.Y(n_3736)
);

INVxp67_ASAP7_75t_L g3737 ( 
.A(n_3538),
.Y(n_3737)
);

AND2x2_ASAP7_75t_L g3738 ( 
.A(n_3546),
.B(n_2826),
.Y(n_3738)
);

HB1xp67_ASAP7_75t_L g3739 ( 
.A(n_3516),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3553),
.Y(n_3740)
);

AND2x2_ASAP7_75t_L g3741 ( 
.A(n_3546),
.B(n_3123),
.Y(n_3741)
);

HB1xp67_ASAP7_75t_L g3742 ( 
.A(n_3516),
.Y(n_3742)
);

CKINVDCx5p33_ASAP7_75t_R g3743 ( 
.A(n_3566),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3545),
.B(n_3123),
.Y(n_3744)
);

OR2x2_ASAP7_75t_L g3745 ( 
.A(n_3572),
.B(n_274),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3553),
.Y(n_3746)
);

AND2x2_ASAP7_75t_L g3747 ( 
.A(n_3552),
.B(n_275),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3574),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3574),
.Y(n_3749)
);

AND2x4_ASAP7_75t_L g3750 ( 
.A(n_3596),
.B(n_275),
.Y(n_3750)
);

HB1xp67_ASAP7_75t_L g3751 ( 
.A(n_3529),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3613),
.Y(n_3752)
);

INVx3_ASAP7_75t_L g3753 ( 
.A(n_3549),
.Y(n_3753)
);

AND2x2_ASAP7_75t_L g3754 ( 
.A(n_3552),
.B(n_276),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_3609),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3690),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3656),
.Y(n_3757)
);

AND2x2_ASAP7_75t_L g3758 ( 
.A(n_3657),
.B(n_3663),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3656),
.Y(n_3759)
);

NOR2xp33_ASAP7_75t_L g3760 ( 
.A(n_3701),
.B(n_3612),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3671),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3671),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_3699),
.B(n_3624),
.Y(n_3763)
);

AND2x4_ASAP7_75t_L g3764 ( 
.A(n_3670),
.B(n_3628),
.Y(n_3764)
);

AND2x2_ASAP7_75t_L g3765 ( 
.A(n_3657),
.B(n_3563),
.Y(n_3765)
);

AND2x4_ASAP7_75t_SL g3766 ( 
.A(n_3722),
.B(n_3694),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3673),
.B(n_3670),
.Y(n_3767)
);

AND2x2_ASAP7_75t_L g3768 ( 
.A(n_3663),
.B(n_3563),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3682),
.Y(n_3769)
);

INVx2_ASAP7_75t_SL g3770 ( 
.A(n_3722),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_3673),
.B(n_3628),
.Y(n_3771)
);

AND2x2_ASAP7_75t_L g3772 ( 
.A(n_3678),
.B(n_3635),
.Y(n_3772)
);

INVx2_ASAP7_75t_L g3773 ( 
.A(n_3694),
.Y(n_3773)
);

AND2x2_ASAP7_75t_L g3774 ( 
.A(n_3678),
.B(n_3635),
.Y(n_3774)
);

BUFx2_ASAP7_75t_L g3775 ( 
.A(n_3694),
.Y(n_3775)
);

AND2x2_ASAP7_75t_L g3776 ( 
.A(n_3679),
.B(n_3659),
.Y(n_3776)
);

AOI21xp5_ASAP7_75t_L g3777 ( 
.A1(n_3666),
.A2(n_3582),
.B(n_3595),
.Y(n_3777)
);

INVx3_ASAP7_75t_L g3778 ( 
.A(n_3694),
.Y(n_3778)
);

OAI221xp5_ASAP7_75t_SL g3779 ( 
.A1(n_3658),
.A2(n_3599),
.B1(n_3583),
.B2(n_3619),
.C(n_3625),
.Y(n_3779)
);

INVx2_ASAP7_75t_L g3780 ( 
.A(n_3694),
.Y(n_3780)
);

AND2x4_ASAP7_75t_L g3781 ( 
.A(n_3662),
.B(n_3529),
.Y(n_3781)
);

NAND2xp5_ASAP7_75t_L g3782 ( 
.A(n_3642),
.B(n_3543),
.Y(n_3782)
);

AND2x2_ASAP7_75t_L g3783 ( 
.A(n_3679),
.B(n_3622),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3672),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3659),
.B(n_3655),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3672),
.Y(n_3786)
);

AND2x2_ASAP7_75t_L g3787 ( 
.A(n_3655),
.B(n_3680),
.Y(n_3787)
);

BUFx3_ASAP7_75t_L g3788 ( 
.A(n_3722),
.Y(n_3788)
);

INVxp67_ASAP7_75t_SL g3789 ( 
.A(n_3667),
.Y(n_3789)
);

NAND2x1_ASAP7_75t_L g3790 ( 
.A(n_3711),
.B(n_3549),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3680),
.B(n_3622),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3675),
.Y(n_3792)
);

AND2x4_ASAP7_75t_L g3793 ( 
.A(n_3662),
.B(n_3549),
.Y(n_3793)
);

AND2x2_ASAP7_75t_L g3794 ( 
.A(n_3686),
.B(n_3641),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3675),
.Y(n_3795)
);

OR2x2_ASAP7_75t_L g3796 ( 
.A(n_3707),
.B(n_3543),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3676),
.Y(n_3797)
);

BUFx3_ASAP7_75t_L g3798 ( 
.A(n_3722),
.Y(n_3798)
);

AND2x2_ASAP7_75t_L g3799 ( 
.A(n_3686),
.B(n_3641),
.Y(n_3799)
);

AND2x2_ASAP7_75t_L g3800 ( 
.A(n_3648),
.B(n_3632),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3676),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3684),
.Y(n_3802)
);

NAND3xp33_ASAP7_75t_L g3803 ( 
.A(n_3711),
.B(n_3550),
.C(n_3554),
.Y(n_3803)
);

INVx2_ASAP7_75t_L g3804 ( 
.A(n_3722),
.Y(n_3804)
);

NAND2x1p5_ASAP7_75t_L g3805 ( 
.A(n_3747),
.B(n_3548),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3684),
.Y(n_3806)
);

AND2x4_ASAP7_75t_L g3807 ( 
.A(n_3662),
.B(n_3520),
.Y(n_3807)
);

NOR2xp33_ASAP7_75t_R g3808 ( 
.A(n_3743),
.B(n_3548),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_L g3809 ( 
.A(n_3642),
.B(n_3588),
.Y(n_3809)
);

AND2x2_ASAP7_75t_L g3810 ( 
.A(n_3648),
.B(n_3632),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3649),
.B(n_3581),
.Y(n_3811)
);

AND2x2_ASAP7_75t_L g3812 ( 
.A(n_3649),
.B(n_3627),
.Y(n_3812)
);

AND2x2_ASAP7_75t_L g3813 ( 
.A(n_3719),
.B(n_3627),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3650),
.B(n_3620),
.Y(n_3814)
);

AND2x2_ASAP7_75t_L g3815 ( 
.A(n_3719),
.B(n_3520),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3698),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_SL g3817 ( 
.A(n_3743),
.B(n_3732),
.Y(n_3817)
);

AND2x2_ASAP7_75t_L g3818 ( 
.A(n_3721),
.B(n_3526),
.Y(n_3818)
);

BUFx2_ASAP7_75t_L g3819 ( 
.A(n_3753),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3747),
.B(n_3620),
.Y(n_3820)
);

AND2x4_ASAP7_75t_L g3821 ( 
.A(n_3645),
.B(n_3526),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3698),
.Y(n_3822)
);

AND2x2_ASAP7_75t_L g3823 ( 
.A(n_3645),
.B(n_3539),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3754),
.B(n_3564),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3705),
.Y(n_3825)
);

AND2x2_ASAP7_75t_L g3826 ( 
.A(n_3645),
.B(n_3539),
.Y(n_3826)
);

OR2x2_ASAP7_75t_L g3827 ( 
.A(n_3726),
.B(n_3551),
.Y(n_3827)
);

INVx2_ASAP7_75t_L g3828 ( 
.A(n_3664),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3705),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3710),
.Y(n_3830)
);

NAND2x1p5_ASAP7_75t_L g3831 ( 
.A(n_3754),
.B(n_3753),
.Y(n_3831)
);

AND2x2_ASAP7_75t_L g3832 ( 
.A(n_3696),
.B(n_3523),
.Y(n_3832)
);

INVxp67_ASAP7_75t_SL g3833 ( 
.A(n_3654),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3710),
.Y(n_3834)
);

AND2x2_ASAP7_75t_L g3835 ( 
.A(n_3696),
.B(n_3523),
.Y(n_3835)
);

AND2x4_ASAP7_75t_L g3836 ( 
.A(n_3753),
.B(n_3664),
.Y(n_3836)
);

OR2x2_ASAP7_75t_L g3837 ( 
.A(n_3726),
.B(n_3613),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3750),
.B(n_3615),
.Y(n_3838)
);

AND2x2_ASAP7_75t_L g3839 ( 
.A(n_3692),
.B(n_3567),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_L g3840 ( 
.A(n_3750),
.B(n_3615),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_3750),
.B(n_3617),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_3739),
.B(n_3617),
.Y(n_3842)
);

AND2x2_ASAP7_75t_L g3843 ( 
.A(n_3692),
.B(n_3567),
.Y(n_3843)
);

INVx2_ASAP7_75t_L g3844 ( 
.A(n_3664),
.Y(n_3844)
);

AND2x2_ASAP7_75t_L g3845 ( 
.A(n_3751),
.B(n_3567),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3708),
.Y(n_3846)
);

AND2x2_ASAP7_75t_L g3847 ( 
.A(n_3708),
.B(n_3575),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3742),
.B(n_3598),
.Y(n_3848)
);

AND2x2_ASAP7_75t_L g3849 ( 
.A(n_3708),
.B(n_3575),
.Y(n_3849)
);

AOI22xp5_ASAP7_75t_L g3850 ( 
.A1(n_3777),
.A2(n_3661),
.B1(n_3737),
.B2(n_3647),
.Y(n_3850)
);

AND2x2_ASAP7_75t_L g3851 ( 
.A(n_3758),
.B(n_3785),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3758),
.B(n_3665),
.Y(n_3852)
);

AND2x2_ASAP7_75t_L g3853 ( 
.A(n_3785),
.B(n_3740),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3778),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_3789),
.B(n_3725),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_3787),
.B(n_3725),
.Y(n_3856)
);

OR2x2_ASAP7_75t_L g3857 ( 
.A(n_3796),
.B(n_3652),
.Y(n_3857)
);

OR2x2_ASAP7_75t_L g3858 ( 
.A(n_3796),
.B(n_3652),
.Y(n_3858)
);

AND2x2_ASAP7_75t_L g3859 ( 
.A(n_3787),
.B(n_3740),
.Y(n_3859)
);

AND2x2_ASAP7_75t_L g3860 ( 
.A(n_3794),
.B(n_3746),
.Y(n_3860)
);

OR2x2_ASAP7_75t_L g3861 ( 
.A(n_3756),
.B(n_3720),
.Y(n_3861)
);

AND2x2_ASAP7_75t_L g3862 ( 
.A(n_3794),
.B(n_3746),
.Y(n_3862)
);

HB1xp67_ASAP7_75t_L g3863 ( 
.A(n_3775),
.Y(n_3863)
);

AND2x2_ASAP7_75t_L g3864 ( 
.A(n_3799),
.B(n_3720),
.Y(n_3864)
);

INVx2_ASAP7_75t_L g3865 ( 
.A(n_3778),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3833),
.B(n_3725),
.Y(n_3866)
);

AND2x2_ASAP7_75t_L g3867 ( 
.A(n_3799),
.B(n_3776),
.Y(n_3867)
);

AND2x2_ASAP7_75t_L g3868 ( 
.A(n_3776),
.B(n_3730),
.Y(n_3868)
);

INVx2_ASAP7_75t_L g3869 ( 
.A(n_3778),
.Y(n_3869)
);

OR2x2_ASAP7_75t_L g3870 ( 
.A(n_3756),
.B(n_3730),
.Y(n_3870)
);

AND2x2_ASAP7_75t_L g3871 ( 
.A(n_3768),
.B(n_3731),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3775),
.Y(n_3872)
);

AND2x2_ASAP7_75t_L g3873 ( 
.A(n_3768),
.B(n_3731),
.Y(n_3873)
);

OR2x2_ASAP7_75t_L g3874 ( 
.A(n_3827),
.B(n_3702),
.Y(n_3874)
);

AND2x2_ASAP7_75t_L g3875 ( 
.A(n_3765),
.B(n_3755),
.Y(n_3875)
);

OR2x2_ASAP7_75t_L g3876 ( 
.A(n_3827),
.B(n_3702),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3819),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_L g3878 ( 
.A(n_3818),
.B(n_3704),
.Y(n_3878)
);

AND2x2_ASAP7_75t_L g3879 ( 
.A(n_3765),
.B(n_3755),
.Y(n_3879)
);

AND2x4_ASAP7_75t_L g3880 ( 
.A(n_3766),
.B(n_3715),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_3818),
.B(n_3733),
.Y(n_3881)
);

AND2x2_ASAP7_75t_L g3882 ( 
.A(n_3813),
.B(n_3734),
.Y(n_3882)
);

AND2x2_ASAP7_75t_L g3883 ( 
.A(n_3813),
.B(n_3734),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3832),
.B(n_3715),
.Y(n_3884)
);

AND2x2_ASAP7_75t_L g3885 ( 
.A(n_3832),
.B(n_3646),
.Y(n_3885)
);

OR2x2_ASAP7_75t_L g3886 ( 
.A(n_3769),
.B(n_3752),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3819),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3757),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3757),
.Y(n_3889)
);

OR2x2_ASAP7_75t_L g3890 ( 
.A(n_3837),
.B(n_3752),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3759),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3759),
.Y(n_3892)
);

AND2x2_ASAP7_75t_L g3893 ( 
.A(n_3835),
.B(n_3712),
.Y(n_3893)
);

NOR2x1_ASAP7_75t_L g3894 ( 
.A(n_3788),
.B(n_3745),
.Y(n_3894)
);

AND2x4_ASAP7_75t_L g3895 ( 
.A(n_3766),
.B(n_3643),
.Y(n_3895)
);

OR2x2_ASAP7_75t_L g3896 ( 
.A(n_3837),
.B(n_3668),
.Y(n_3896)
);

OR2x2_ASAP7_75t_L g3897 ( 
.A(n_3767),
.B(n_3668),
.Y(n_3897)
);

BUFx2_ASAP7_75t_L g3898 ( 
.A(n_3808),
.Y(n_3898)
);

AND2x2_ASAP7_75t_L g3899 ( 
.A(n_3835),
.B(n_3712),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3761),
.Y(n_3900)
);

AND2x2_ASAP7_75t_L g3901 ( 
.A(n_3847),
.B(n_3716),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3761),
.Y(n_3902)
);

INVxp67_ASAP7_75t_SL g3903 ( 
.A(n_3805),
.Y(n_3903)
);

NOR2x1_ASAP7_75t_L g3904 ( 
.A(n_3788),
.B(n_3798),
.Y(n_3904)
);

INVx2_ASAP7_75t_SL g3905 ( 
.A(n_3836),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3836),
.Y(n_3906)
);

AND2x2_ASAP7_75t_L g3907 ( 
.A(n_3847),
.B(n_3716),
.Y(n_3907)
);

AND2x2_ASAP7_75t_L g3908 ( 
.A(n_3849),
.B(n_3735),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3762),
.Y(n_3909)
);

AND2x2_ASAP7_75t_L g3910 ( 
.A(n_3849),
.B(n_3735),
.Y(n_3910)
);

AND2x2_ASAP7_75t_L g3911 ( 
.A(n_3812),
.B(n_3651),
.Y(n_3911)
);

INVxp67_ASAP7_75t_L g3912 ( 
.A(n_3798),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3836),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3771),
.B(n_3745),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3762),
.Y(n_3915)
);

AND2x2_ASAP7_75t_L g3916 ( 
.A(n_3812),
.B(n_3651),
.Y(n_3916)
);

AND2x2_ASAP7_75t_L g3917 ( 
.A(n_3791),
.B(n_3738),
.Y(n_3917)
);

AND2x2_ASAP7_75t_L g3918 ( 
.A(n_3791),
.B(n_3771),
.Y(n_3918)
);

AND2x2_ASAP7_75t_L g3919 ( 
.A(n_3815),
.B(n_3738),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3831),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3764),
.B(n_3815),
.Y(n_3921)
);

AOI22xp5_ASAP7_75t_L g3922 ( 
.A1(n_3760),
.A2(n_3677),
.B1(n_3524),
.B2(n_3630),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3786),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3786),
.Y(n_3924)
);

NAND2xp5_ASAP7_75t_L g3925 ( 
.A(n_3764),
.B(n_3729),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3764),
.B(n_3714),
.Y(n_3926)
);

NOR2xp33_ASAP7_75t_L g3927 ( 
.A(n_3817),
.B(n_3568),
.Y(n_3927)
);

INVx2_ASAP7_75t_L g3928 ( 
.A(n_3831),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3792),
.Y(n_3929)
);

INVx2_ASAP7_75t_L g3930 ( 
.A(n_3831),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3792),
.Y(n_3931)
);

OR2x2_ASAP7_75t_L g3932 ( 
.A(n_3820),
.B(n_3748),
.Y(n_3932)
);

NAND2x1p5_ASAP7_75t_L g3933 ( 
.A(n_3790),
.B(n_3770),
.Y(n_3933)
);

AND2x4_ASAP7_75t_SL g3934 ( 
.A(n_3781),
.B(n_3681),
.Y(n_3934)
);

AND2x2_ASAP7_75t_L g3935 ( 
.A(n_3783),
.B(n_3749),
.Y(n_3935)
);

NAND2x1_ASAP7_75t_L g3936 ( 
.A(n_3793),
.B(n_3723),
.Y(n_3936)
);

OR2x2_ASAP7_75t_L g3937 ( 
.A(n_3773),
.B(n_3714),
.Y(n_3937)
);

INVx2_ASAP7_75t_L g3938 ( 
.A(n_3790),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3805),
.Y(n_3939)
);

INVx3_ASAP7_75t_L g3940 ( 
.A(n_3793),
.Y(n_3940)
);

AND2x4_ASAP7_75t_L g3941 ( 
.A(n_3773),
.B(n_3780),
.Y(n_3941)
);

AND2x2_ASAP7_75t_L g3942 ( 
.A(n_3783),
.B(n_3577),
.Y(n_3942)
);

AND2x2_ASAP7_75t_L g3943 ( 
.A(n_3800),
.B(n_3577),
.Y(n_3943)
);

OAI21xp5_ASAP7_75t_L g3944 ( 
.A1(n_3927),
.A2(n_3779),
.B(n_3803),
.Y(n_3944)
);

OR2x2_ASAP7_75t_L g3945 ( 
.A(n_3878),
.B(n_3763),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3851),
.B(n_3770),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3851),
.B(n_3804),
.Y(n_3947)
);

OR2x2_ASAP7_75t_L g3948 ( 
.A(n_3881),
.B(n_3824),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3863),
.Y(n_3949)
);

AND2x2_ASAP7_75t_L g3950 ( 
.A(n_3867),
.B(n_3800),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3867),
.B(n_3804),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3918),
.B(n_3780),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3933),
.Y(n_3953)
);

NOR2x1_ASAP7_75t_L g3954 ( 
.A(n_3904),
.B(n_3898),
.Y(n_3954)
);

OR2x2_ASAP7_75t_L g3955 ( 
.A(n_3914),
.B(n_3866),
.Y(n_3955)
);

AND2x2_ASAP7_75t_L g3956 ( 
.A(n_3934),
.B(n_3823),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_3918),
.B(n_3805),
.Y(n_3957)
);

NOR2xp33_ASAP7_75t_SL g3958 ( 
.A(n_3898),
.B(n_3781),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_SL g3959 ( 
.A(n_3894),
.B(n_3793),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_L g3960 ( 
.A(n_3871),
.B(n_3823),
.Y(n_3960)
);

AND2x2_ASAP7_75t_L g3961 ( 
.A(n_3934),
.B(n_3810),
.Y(n_3961)
);

INVx2_ASAP7_75t_L g3962 ( 
.A(n_3933),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_L g3963 ( 
.A(n_3871),
.B(n_3826),
.Y(n_3963)
);

AND2x2_ASAP7_75t_L g3964 ( 
.A(n_3942),
.B(n_3810),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3890),
.Y(n_3965)
);

NAND4xp25_ASAP7_75t_L g3966 ( 
.A(n_3850),
.B(n_3782),
.C(n_3774),
.D(n_3772),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3890),
.Y(n_3967)
);

BUFx2_ASAP7_75t_L g3968 ( 
.A(n_3940),
.Y(n_3968)
);

AND2x4_ASAP7_75t_SL g3969 ( 
.A(n_3880),
.B(n_3781),
.Y(n_3969)
);

INVx2_ASAP7_75t_L g3970 ( 
.A(n_3933),
.Y(n_3970)
);

AND2x2_ASAP7_75t_L g3971 ( 
.A(n_3942),
.B(n_3826),
.Y(n_3971)
);

AND2x2_ASAP7_75t_L g3972 ( 
.A(n_3911),
.B(n_3772),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3911),
.B(n_3774),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_3873),
.B(n_3807),
.Y(n_3974)
);

AND2x2_ASAP7_75t_L g3975 ( 
.A(n_3940),
.B(n_3807),
.Y(n_3975)
);

INVx1_ASAP7_75t_L g3976 ( 
.A(n_3884),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3873),
.B(n_3807),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3884),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_3885),
.B(n_3821),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3882),
.Y(n_3980)
);

AND2x2_ASAP7_75t_L g3981 ( 
.A(n_3916),
.B(n_3821),
.Y(n_3981)
);

OAI21xp5_ASAP7_75t_L g3982 ( 
.A1(n_3922),
.A2(n_3843),
.B(n_3839),
.Y(n_3982)
);

INVx2_ASAP7_75t_L g3983 ( 
.A(n_3940),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_3885),
.B(n_3821),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_3880),
.B(n_3838),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3882),
.Y(n_3986)
);

INVx2_ASAP7_75t_L g3987 ( 
.A(n_3880),
.Y(n_3987)
);

INVx1_ASAP7_75t_SL g3988 ( 
.A(n_3896),
.Y(n_3988)
);

AND3x2_ASAP7_75t_L g3989 ( 
.A(n_3903),
.B(n_3845),
.C(n_3844),
.Y(n_3989)
);

INVx3_ASAP7_75t_SL g3990 ( 
.A(n_3895),
.Y(n_3990)
);

OR2x2_ASAP7_75t_L g3991 ( 
.A(n_3852),
.B(n_3840),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3883),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_L g3993 ( 
.A(n_3868),
.B(n_3841),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3868),
.B(n_3809),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3883),
.Y(n_3995)
);

AND2x2_ASAP7_75t_L g3996 ( 
.A(n_3943),
.B(n_3828),
.Y(n_3996)
);

AND2x2_ASAP7_75t_L g3997 ( 
.A(n_3916),
.B(n_3848),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3859),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3859),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3912),
.B(n_3811),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3874),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3875),
.B(n_3814),
.Y(n_4002)
);

INVx1_ASAP7_75t_SL g4003 ( 
.A(n_3896),
.Y(n_4003)
);

INVx2_ASAP7_75t_L g4004 ( 
.A(n_3905),
.Y(n_4004)
);

NOR2xp33_ASAP7_75t_L g4005 ( 
.A(n_3921),
.B(n_3842),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_L g4006 ( 
.A(n_3875),
.B(n_3839),
.Y(n_4006)
);

AND2x4_ASAP7_75t_L g4007 ( 
.A(n_3905),
.B(n_3828),
.Y(n_4007)
);

INVx2_ASAP7_75t_L g4008 ( 
.A(n_3895),
.Y(n_4008)
);

OR2x6_ASAP7_75t_L g4009 ( 
.A(n_3872),
.B(n_3844),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3874),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3876),
.Y(n_4011)
);

NOR2xp33_ASAP7_75t_L g4012 ( 
.A(n_3855),
.B(n_3843),
.Y(n_4012)
);

INVx2_ASAP7_75t_L g4013 ( 
.A(n_3895),
.Y(n_4013)
);

OR2x2_ASAP7_75t_L g4014 ( 
.A(n_3897),
.B(n_3717),
.Y(n_4014)
);

AND2x2_ASAP7_75t_L g4015 ( 
.A(n_3943),
.B(n_3893),
.Y(n_4015)
);

OR2x2_ASAP7_75t_L g4016 ( 
.A(n_3897),
.B(n_3724),
.Y(n_4016)
);

AND2x2_ASAP7_75t_L g4017 ( 
.A(n_3893),
.B(n_3846),
.Y(n_4017)
);

INVx2_ASAP7_75t_L g4018 ( 
.A(n_3938),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3876),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3853),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3853),
.Y(n_4021)
);

NOR2xp33_ASAP7_75t_L g4022 ( 
.A(n_3939),
.B(n_3846),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3877),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3879),
.B(n_3784),
.Y(n_4024)
);

OR2x2_ASAP7_75t_L g4025 ( 
.A(n_3856),
.B(n_3724),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3887),
.Y(n_4026)
);

INVx2_ASAP7_75t_L g4027 ( 
.A(n_3938),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_L g4028 ( 
.A(n_3879),
.B(n_3806),
.Y(n_4028)
);

AND2x2_ASAP7_75t_L g4029 ( 
.A(n_3899),
.B(n_3845),
.Y(n_4029)
);

OR2x2_ASAP7_75t_L g4030 ( 
.A(n_3861),
.B(n_3644),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3935),
.B(n_3906),
.Y(n_4031)
);

AND2x2_ASAP7_75t_L g4032 ( 
.A(n_3860),
.B(n_3532),
.Y(n_4032)
);

AND2x2_ASAP7_75t_L g4033 ( 
.A(n_3899),
.B(n_3688),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3937),
.Y(n_4034)
);

AND2x2_ASAP7_75t_L g4035 ( 
.A(n_3950),
.B(n_3860),
.Y(n_4035)
);

OR2x2_ASAP7_75t_L g4036 ( 
.A(n_3988),
.B(n_4003),
.Y(n_4036)
);

AOI22xp5_ASAP7_75t_L g4037 ( 
.A1(n_3958),
.A2(n_3939),
.B1(n_3935),
.B2(n_3913),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_3968),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3983),
.Y(n_4039)
);

AND2x2_ASAP7_75t_L g4040 ( 
.A(n_3950),
.B(n_3862),
.Y(n_4040)
);

AND2x2_ASAP7_75t_L g4041 ( 
.A(n_3971),
.B(n_3862),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_L g4042 ( 
.A(n_3971),
.B(n_3906),
.Y(n_4042)
);

OR2x2_ASAP7_75t_L g4043 ( 
.A(n_4006),
.B(n_3861),
.Y(n_4043)
);

AOI22xp5_ASAP7_75t_L g4044 ( 
.A1(n_3944),
.A2(n_3913),
.B1(n_3864),
.B2(n_3920),
.Y(n_4044)
);

INVxp67_ASAP7_75t_SL g4045 ( 
.A(n_3954),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3983),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_4015),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_4015),
.Y(n_4048)
);

HB1xp67_ASAP7_75t_L g4049 ( 
.A(n_4009),
.Y(n_4049)
);

OR2x2_ASAP7_75t_L g4050 ( 
.A(n_3951),
.B(n_3870),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_L g4051 ( 
.A(n_3972),
.B(n_3941),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_4004),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_4004),
.Y(n_4053)
);

OR2x2_ASAP7_75t_L g4054 ( 
.A(n_3947),
.B(n_3870),
.Y(n_4054)
);

OR2x2_ASAP7_75t_L g4055 ( 
.A(n_4031),
.B(n_3925),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_4017),
.Y(n_4056)
);

NAND2xp33_ASAP7_75t_L g4057 ( 
.A(n_3990),
.B(n_3857),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_L g4058 ( 
.A(n_3976),
.B(n_3941),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_4017),
.Y(n_4059)
);

NOR3xp33_ASAP7_75t_L g4060 ( 
.A(n_3982),
.B(n_3926),
.C(n_3920),
.Y(n_4060)
);

AND2x2_ASAP7_75t_L g4061 ( 
.A(n_3973),
.B(n_3864),
.Y(n_4061)
);

OR2x2_ASAP7_75t_L g4062 ( 
.A(n_3952),
.B(n_3857),
.Y(n_4062)
);

INVx1_ASAP7_75t_SL g4063 ( 
.A(n_3990),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3978),
.Y(n_4064)
);

NOR2xp33_ASAP7_75t_SL g4065 ( 
.A(n_3987),
.B(n_3928),
.Y(n_4065)
);

AND2x2_ASAP7_75t_L g4066 ( 
.A(n_3964),
.B(n_3901),
.Y(n_4066)
);

AOI22xp33_ASAP7_75t_L g4067 ( 
.A1(n_3966),
.A2(n_3907),
.B1(n_3901),
.B2(n_3908),
.Y(n_4067)
);

NAND2x1_ASAP7_75t_L g4068 ( 
.A(n_3975),
.B(n_3928),
.Y(n_4068)
);

INVx2_ASAP7_75t_L g4069 ( 
.A(n_3969),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3964),
.Y(n_4070)
);

INVx1_ASAP7_75t_SL g4071 ( 
.A(n_3969),
.Y(n_4071)
);

INVx2_ASAP7_75t_L g4072 ( 
.A(n_3975),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_3981),
.B(n_3907),
.Y(n_4073)
);

AND2x4_ASAP7_75t_L g4074 ( 
.A(n_3987),
.B(n_3941),
.Y(n_4074)
);

INVx2_ASAP7_75t_SL g4075 ( 
.A(n_4008),
.Y(n_4075)
);

OR2x2_ASAP7_75t_L g4076 ( 
.A(n_3960),
.B(n_3858),
.Y(n_4076)
);

INVx2_ASAP7_75t_L g4077 ( 
.A(n_4007),
.Y(n_4077)
);

AND2x4_ASAP7_75t_L g4078 ( 
.A(n_4008),
.B(n_3930),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_4034),
.Y(n_4079)
);

OR2x2_ASAP7_75t_L g4080 ( 
.A(n_3963),
.B(n_3858),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_L g4081 ( 
.A(n_3949),
.B(n_3854),
.Y(n_4081)
);

INVx2_ASAP7_75t_L g4082 ( 
.A(n_4007),
.Y(n_4082)
);

AOI22xp33_ASAP7_75t_L g4083 ( 
.A1(n_3961),
.A2(n_3910),
.B1(n_3908),
.B2(n_3919),
.Y(n_4083)
);

OR2x2_ASAP7_75t_L g4084 ( 
.A(n_3993),
.B(n_3932),
.Y(n_4084)
);

NOR5xp2_ASAP7_75t_L g4085 ( 
.A(n_4023),
.B(n_4026),
.C(n_3967),
.D(n_3965),
.E(n_4010),
.Y(n_4085)
);

AOI21xp33_ASAP7_75t_L g4086 ( 
.A1(n_3959),
.A2(n_3930),
.B(n_3865),
.Y(n_4086)
);

NOR2x1_ASAP7_75t_L g4087 ( 
.A(n_3953),
.B(n_3854),
.Y(n_4087)
);

OR2x2_ASAP7_75t_L g4088 ( 
.A(n_3946),
.B(n_3932),
.Y(n_4088)
);

OR2x2_ASAP7_75t_L g4089 ( 
.A(n_3998),
.B(n_3886),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3999),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_4013),
.B(n_3865),
.Y(n_4091)
);

OR2x2_ASAP7_75t_L g4092 ( 
.A(n_4020),
.B(n_3886),
.Y(n_4092)
);

AND2x2_ASAP7_75t_L g4093 ( 
.A(n_3961),
.B(n_3910),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_3956),
.B(n_3919),
.Y(n_4094)
);

AND2x2_ASAP7_75t_L g4095 ( 
.A(n_3997),
.B(n_3917),
.Y(n_4095)
);

INVxp67_ASAP7_75t_L g4096 ( 
.A(n_3959),
.Y(n_4096)
);

OR2x2_ASAP7_75t_L g4097 ( 
.A(n_4021),
.B(n_3869),
.Y(n_4097)
);

INVx1_ASAP7_75t_SL g4098 ( 
.A(n_3989),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_4013),
.B(n_3869),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_3996),
.B(n_3917),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3980),
.Y(n_4101)
);

INVxp67_ASAP7_75t_L g4102 ( 
.A(n_4012),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_3986),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_3996),
.B(n_3992),
.Y(n_4104)
);

AND2x2_ASAP7_75t_L g4105 ( 
.A(n_4032),
.B(n_3937),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_L g4106 ( 
.A(n_3995),
.B(n_3888),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_4007),
.Y(n_4107)
);

INVx1_ASAP7_75t_SL g4108 ( 
.A(n_3989),
.Y(n_4108)
);

INVx2_ASAP7_75t_L g4109 ( 
.A(n_4009),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_4018),
.Y(n_4110)
);

HB1xp67_ASAP7_75t_L g4111 ( 
.A(n_4009),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_4018),
.Y(n_4112)
);

INVx2_ASAP7_75t_L g4113 ( 
.A(n_3953),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_4027),
.Y(n_4114)
);

AOI22xp5_ASAP7_75t_L g4115 ( 
.A1(n_4012),
.A2(n_3891),
.B1(n_3892),
.B2(n_3889),
.Y(n_4115)
);

INVx2_ASAP7_75t_SL g4116 ( 
.A(n_3962),
.Y(n_4116)
);

NAND2x1p5_ASAP7_75t_L g4117 ( 
.A(n_3962),
.B(n_3936),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_4027),
.Y(n_4118)
);

XOR2x2_ASAP7_75t_L g4119 ( 
.A(n_4044),
.B(n_3945),
.Y(n_4119)
);

OAI22xp5_ASAP7_75t_L g4120 ( 
.A1(n_4096),
.A2(n_3984),
.B1(n_3979),
.B2(n_3977),
.Y(n_4120)
);

OAI22xp33_ASAP7_75t_SL g4121 ( 
.A1(n_4098),
.A2(n_4011),
.B1(n_4019),
.B2(n_4001),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_4107),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_4049),
.Y(n_4123)
);

AOI211xp5_ASAP7_75t_SL g4124 ( 
.A1(n_4057),
.A2(n_4022),
.B(n_4000),
.C(n_3985),
.Y(n_4124)
);

OAI22xp5_ASAP7_75t_L g4125 ( 
.A1(n_4045),
.A2(n_3974),
.B1(n_4002),
.B2(n_3957),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_4111),
.Y(n_4126)
);

AOI21xp33_ASAP7_75t_SL g4127 ( 
.A1(n_4036),
.A2(n_4016),
.B(n_3955),
.Y(n_4127)
);

OAI21xp33_ASAP7_75t_SL g4128 ( 
.A1(n_4098),
.A2(n_3970),
.B(n_4029),
.Y(n_4128)
);

AOI22xp5_ASAP7_75t_L g4129 ( 
.A1(n_4108),
.A2(n_4060),
.B1(n_4065),
.B2(n_4044),
.Y(n_4129)
);

AOI22xp5_ASAP7_75t_L g4130 ( 
.A1(n_4108),
.A2(n_4005),
.B1(n_3970),
.B2(n_4022),
.Y(n_4130)
);

XNOR2x1_ASAP7_75t_L g4131 ( 
.A(n_4063),
.B(n_3948),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_4077),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_4082),
.Y(n_4133)
);

OR2x2_ASAP7_75t_L g4134 ( 
.A(n_4063),
.B(n_3994),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_4071),
.B(n_4005),
.Y(n_4135)
);

OAI21xp5_ASAP7_75t_L g4136 ( 
.A1(n_4037),
.A2(n_4028),
.B(n_4024),
.Y(n_4136)
);

AOI21xp33_ASAP7_75t_SL g4137 ( 
.A1(n_4037),
.A2(n_3991),
.B(n_4025),
.Y(n_4137)
);

O2A1O1Ixp33_ASAP7_75t_L g4138 ( 
.A1(n_4086),
.A2(n_3902),
.B(n_3909),
.C(n_3900),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_4074),
.Y(n_4139)
);

OAI21xp5_ASAP7_75t_L g4140 ( 
.A1(n_4102),
.A2(n_4029),
.B(n_4014),
.Y(n_4140)
);

OAI22xp33_ASAP7_75t_SL g4141 ( 
.A1(n_4065),
.A2(n_4030),
.B1(n_3923),
.B2(n_3924),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_4071),
.B(n_4033),
.Y(n_4142)
);

XOR2x2_ASAP7_75t_L g4143 ( 
.A(n_4061),
.B(n_4033),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4074),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_4035),
.Y(n_4145)
);

OAI22xp33_ASAP7_75t_L g4146 ( 
.A1(n_4051),
.A2(n_3653),
.B1(n_3669),
.B2(n_3660),
.Y(n_4146)
);

AOI22xp33_ASAP7_75t_L g4147 ( 
.A1(n_4069),
.A2(n_3557),
.B1(n_3660),
.B2(n_3653),
.Y(n_4147)
);

HB1xp67_ASAP7_75t_L g4148 ( 
.A(n_4068),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_4040),
.Y(n_4149)
);

INVx2_ASAP7_75t_L g4150 ( 
.A(n_4078),
.Y(n_4150)
);

AOI21xp33_ASAP7_75t_SL g4151 ( 
.A1(n_4062),
.A2(n_3931),
.B(n_3929),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_4041),
.Y(n_4152)
);

AND2x4_ASAP7_75t_L g4153 ( 
.A(n_4075),
.B(n_4109),
.Y(n_4153)
);

INVxp33_ASAP7_75t_L g4154 ( 
.A(n_4066),
.Y(n_4154)
);

AOI21xp33_ASAP7_75t_L g4155 ( 
.A1(n_4076),
.A2(n_3915),
.B(n_3822),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_4047),
.Y(n_4156)
);

NAND3xp33_ASAP7_75t_L g4157 ( 
.A(n_4085),
.B(n_3825),
.C(n_3816),
.Y(n_4157)
);

INVx2_ASAP7_75t_SL g4158 ( 
.A(n_4093),
.Y(n_4158)
);

OAI21xp33_ASAP7_75t_L g4159 ( 
.A1(n_4083),
.A2(n_3830),
.B(n_3829),
.Y(n_4159)
);

AOI22xp5_ASAP7_75t_L g4160 ( 
.A1(n_4048),
.A2(n_3795),
.B1(n_3801),
.B2(n_3797),
.Y(n_4160)
);

INVxp67_ASAP7_75t_SL g4161 ( 
.A(n_4087),
.Y(n_4161)
);

OAI21xp33_ASAP7_75t_L g4162 ( 
.A1(n_4067),
.A2(n_3834),
.B(n_3797),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_4078),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_4094),
.B(n_3795),
.Y(n_4164)
);

OAI31xp33_ASAP7_75t_L g4165 ( 
.A1(n_4117),
.A2(n_3802),
.A3(n_3801),
.B(n_3669),
.Y(n_4165)
);

XNOR2x1_ASAP7_75t_L g4166 ( 
.A(n_4073),
.B(n_3524),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_4058),
.Y(n_4167)
);

OAI22xp33_ASAP7_75t_SL g4168 ( 
.A1(n_4117),
.A2(n_3802),
.B1(n_3685),
.B2(n_3713),
.Y(n_4168)
);

OAI21xp33_ASAP7_75t_L g4169 ( 
.A1(n_4095),
.A2(n_3685),
.B(n_3713),
.Y(n_4169)
);

XOR2x2_ASAP7_75t_L g4170 ( 
.A(n_4042),
.B(n_3631),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_4058),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_4072),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4056),
.Y(n_4173)
);

INVx2_ASAP7_75t_L g4174 ( 
.A(n_4059),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_4038),
.B(n_3693),
.Y(n_4175)
);

INVx2_ASAP7_75t_SL g4176 ( 
.A(n_4105),
.Y(n_4176)
);

AO21x1_ASAP7_75t_L g4177 ( 
.A1(n_4086),
.A2(n_3697),
.B(n_3695),
.Y(n_4177)
);

NAND3xp33_ASAP7_75t_SL g4178 ( 
.A(n_4080),
.B(n_3639),
.C(n_3640),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_4070),
.Y(n_4179)
);

AOI21xp5_ASAP7_75t_L g4180 ( 
.A1(n_4104),
.A2(n_3744),
.B(n_3687),
.Y(n_4180)
);

OR2x2_ASAP7_75t_L g4181 ( 
.A(n_4100),
.B(n_3718),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_4091),
.Y(n_4182)
);

O2A1O1Ixp5_ASAP7_75t_L g4183 ( 
.A1(n_4113),
.A2(n_3524),
.B(n_3728),
.C(n_3691),
.Y(n_4183)
);

OAI211xp5_ASAP7_75t_L g4184 ( 
.A1(n_4115),
.A2(n_4099),
.B(n_4081),
.C(n_4053),
.Y(n_4184)
);

AOI21xp33_ASAP7_75t_L g4185 ( 
.A1(n_4050),
.A2(n_3557),
.B(n_3639),
.Y(n_4185)
);

AND2x2_ASAP7_75t_L g4186 ( 
.A(n_4052),
.B(n_3640),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4097),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4163),
.Y(n_4188)
);

INVx2_ASAP7_75t_L g4189 ( 
.A(n_4148),
.Y(n_4189)
);

INVx1_ASAP7_75t_SL g4190 ( 
.A(n_4131),
.Y(n_4190)
);

A2O1A1Ixp33_ASAP7_75t_L g4191 ( 
.A1(n_4129),
.A2(n_4115),
.B(n_4116),
.C(n_4079),
.Y(n_4191)
);

NOR4xp25_ASAP7_75t_L g4192 ( 
.A(n_4128),
.B(n_4046),
.C(n_4039),
.D(n_4110),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4142),
.Y(n_4193)
);

OAI21xp33_ASAP7_75t_L g4194 ( 
.A1(n_4154),
.A2(n_4081),
.B(n_4055),
.Y(n_4194)
);

OR2x2_ASAP7_75t_L g4195 ( 
.A(n_4158),
.B(n_4054),
.Y(n_4195)
);

AND2x2_ASAP7_75t_L g4196 ( 
.A(n_4176),
.B(n_4088),
.Y(n_4196)
);

OAI22xp5_ASAP7_75t_SL g4197 ( 
.A1(n_4161),
.A2(n_4114),
.B1(n_4118),
.B2(n_4112),
.Y(n_4197)
);

AOI222xp33_ASAP7_75t_L g4198 ( 
.A1(n_4119),
.A2(n_4103),
.B1(n_4101),
.B2(n_4090),
.C1(n_4064),
.C2(n_4106),
.Y(n_4198)
);

NAND2xp5_ASAP7_75t_L g4199 ( 
.A(n_4150),
.B(n_4089),
.Y(n_4199)
);

OAI211xp5_ASAP7_75t_SL g4200 ( 
.A1(n_4129),
.A2(n_4084),
.B(n_4043),
.C(n_4106),
.Y(n_4200)
);

OAI22xp5_ASAP7_75t_L g4201 ( 
.A1(n_4157),
.A2(n_4092),
.B1(n_3706),
.B2(n_3683),
.Y(n_4201)
);

A2O1A1Ixp33_ASAP7_75t_L g4202 ( 
.A1(n_4137),
.A2(n_3691),
.B(n_3700),
.C(n_3703),
.Y(n_4202)
);

OAI22xp5_ASAP7_75t_L g4203 ( 
.A1(n_4130),
.A2(n_3718),
.B1(n_3557),
.B2(n_3597),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4139),
.Y(n_4204)
);

NAND2xp33_ASAP7_75t_L g4205 ( 
.A(n_4135),
.B(n_3723),
.Y(n_4205)
);

NOR3xp33_ASAP7_75t_L g4206 ( 
.A(n_4127),
.B(n_3741),
.C(n_3736),
.Y(n_4206)
);

AND2x2_ASAP7_75t_L g4207 ( 
.A(n_4145),
.B(n_3606),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_4153),
.B(n_3723),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_4144),
.Y(n_4209)
);

NOR4xp25_ASAP7_75t_L g4210 ( 
.A(n_4128),
.B(n_3741),
.C(n_3709),
.D(n_3590),
.Y(n_4210)
);

NOR2xp33_ASAP7_75t_L g4211 ( 
.A(n_4134),
.B(n_3723),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4153),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_4177),
.Y(n_4213)
);

AOI22xp5_ASAP7_75t_L g4214 ( 
.A1(n_4149),
.A2(n_4152),
.B1(n_4178),
.B2(n_4120),
.Y(n_4214)
);

OAI21xp5_ASAP7_75t_L g4215 ( 
.A1(n_4121),
.A2(n_3723),
.B(n_3557),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_4123),
.Y(n_4216)
);

OAI221xp5_ASAP7_75t_SL g4217 ( 
.A1(n_4130),
.A2(n_3727),
.B1(n_3573),
.B2(n_3597),
.C(n_3586),
.Y(n_4217)
);

AOI21xp5_ASAP7_75t_L g4218 ( 
.A1(n_4141),
.A2(n_3728),
.B(n_3689),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_L g4219 ( 
.A(n_4124),
.B(n_3723),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4126),
.Y(n_4220)
);

OAI22xp33_ASAP7_75t_SL g4221 ( 
.A1(n_4122),
.A2(n_3728),
.B1(n_3727),
.B2(n_3590),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_4143),
.Y(n_4222)
);

OAI211xp5_ASAP7_75t_SL g4223 ( 
.A1(n_4136),
.A2(n_3589),
.B(n_3586),
.C(n_3573),
.Y(n_4223)
);

NAND3x1_ASAP7_75t_L g4224 ( 
.A(n_4165),
.B(n_4140),
.C(n_4133),
.Y(n_4224)
);

NOR2xp67_ASAP7_75t_L g4225 ( 
.A(n_4184),
.B(n_3589),
.Y(n_4225)
);

OAI22xp5_ASAP7_75t_L g4226 ( 
.A1(n_4166),
.A2(n_3689),
.B1(n_3674),
.B2(n_3534),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_4186),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_4168),
.Y(n_4228)
);

NOR2xp33_ASAP7_75t_L g4229 ( 
.A(n_4125),
.B(n_3674),
.Y(n_4229)
);

INVx1_ASAP7_75t_SL g4230 ( 
.A(n_4187),
.Y(n_4230)
);

OAI321xp33_ASAP7_75t_L g4231 ( 
.A1(n_4146),
.A2(n_3709),
.A3(n_3606),
.B1(n_3592),
.B2(n_3562),
.C(n_3560),
.Y(n_4231)
);

OAI21xp33_ASAP7_75t_L g4232 ( 
.A1(n_4170),
.A2(n_3689),
.B(n_3674),
.Y(n_4232)
);

NOR4xp25_ASAP7_75t_SL g4233 ( 
.A(n_4132),
.B(n_276),
.C(n_277),
.D(n_278),
.Y(n_4233)
);

NAND2x1_ASAP7_75t_L g4234 ( 
.A(n_4160),
.B(n_3584),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_4172),
.B(n_3560),
.Y(n_4235)
);

AND2x2_ASAP7_75t_L g4236 ( 
.A(n_4174),
.B(n_3562),
.Y(n_4236)
);

NOR2xp67_ASAP7_75t_L g4237 ( 
.A(n_4151),
.B(n_278),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_L g4238 ( 
.A(n_4156),
.B(n_4179),
.Y(n_4238)
);

NAND3xp33_ASAP7_75t_SL g4239 ( 
.A(n_4138),
.B(n_4162),
.C(n_4167),
.Y(n_4239)
);

AND2x2_ASAP7_75t_L g4240 ( 
.A(n_4171),
.B(n_3532),
.Y(n_4240)
);

OR2x2_ASAP7_75t_L g4241 ( 
.A(n_4164),
.B(n_3598),
.Y(n_4241)
);

AOI22xp5_ASAP7_75t_L g4242 ( 
.A1(n_4159),
.A2(n_3534),
.B1(n_3535),
.B2(n_3609),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_4160),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_L g4244 ( 
.A(n_4173),
.B(n_3535),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_L g4245 ( 
.A(n_4182),
.B(n_4169),
.Y(n_4245)
);

OR2x2_ASAP7_75t_L g4246 ( 
.A(n_4181),
.B(n_3621),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_SL g4247 ( 
.A(n_4185),
.B(n_3534),
.Y(n_4247)
);

AOI22xp5_ASAP7_75t_L g4248 ( 
.A1(n_4147),
.A2(n_3616),
.B1(n_3605),
.B2(n_3584),
.Y(n_4248)
);

HB1xp67_ASAP7_75t_L g4249 ( 
.A(n_4175),
.Y(n_4249)
);

NOR2xp33_ASAP7_75t_L g4250 ( 
.A(n_4155),
.B(n_3621),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4183),
.Y(n_4251)
);

NOR2xp33_ASAP7_75t_L g4252 ( 
.A(n_4190),
.B(n_4180),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4212),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_4189),
.B(n_4237),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_L g4255 ( 
.A(n_4196),
.B(n_3616),
.Y(n_4255)
);

AOI211xp5_ASAP7_75t_L g4256 ( 
.A1(n_4200),
.A2(n_279),
.B(n_280),
.C(n_281),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_4230),
.B(n_3605),
.Y(n_4257)
);

OAI22x1_ASAP7_75t_L g4258 ( 
.A1(n_4214),
.A2(n_3592),
.B1(n_281),
.B2(n_283),
.Y(n_4258)
);

OR2x2_ASAP7_75t_L g4259 ( 
.A(n_4230),
.B(n_279),
.Y(n_4259)
);

OAI22xp5_ASAP7_75t_L g4260 ( 
.A1(n_4242),
.A2(n_284),
.B1(n_285),
.B2(n_287),
.Y(n_4260)
);

AOI22xp5_ASAP7_75t_L g4261 ( 
.A1(n_4222),
.A2(n_284),
.B1(n_285),
.B2(n_287),
.Y(n_4261)
);

OAI22xp5_ASAP7_75t_L g4262 ( 
.A1(n_4248),
.A2(n_288),
.B1(n_289),
.B2(n_292),
.Y(n_4262)
);

OAI21xp5_ASAP7_75t_L g4263 ( 
.A1(n_4224),
.A2(n_288),
.B(n_292),
.Y(n_4263)
);

AOI221xp5_ASAP7_75t_L g4264 ( 
.A1(n_4239),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.C(n_296),
.Y(n_4264)
);

AOI21xp5_ASAP7_75t_L g4265 ( 
.A1(n_4191),
.A2(n_296),
.B(n_297),
.Y(n_4265)
);

AOI221xp5_ASAP7_75t_L g4266 ( 
.A1(n_4192),
.A2(n_297),
.B1(n_298),
.B2(n_300),
.C(n_301),
.Y(n_4266)
);

OR2x6_ASAP7_75t_L g4267 ( 
.A(n_4195),
.B(n_4199),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4207),
.Y(n_4268)
);

OAI21xp5_ASAP7_75t_SL g4269 ( 
.A1(n_4198),
.A2(n_298),
.B(n_300),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_L g4270 ( 
.A(n_4225),
.B(n_301),
.Y(n_4270)
);

AOI22xp33_ASAP7_75t_L g4271 ( 
.A1(n_4213),
.A2(n_302),
.B1(n_304),
.B2(n_305),
.Y(n_4271)
);

OAI21xp5_ASAP7_75t_L g4272 ( 
.A1(n_4229),
.A2(n_302),
.B(n_304),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4197),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_SL g4274 ( 
.A(n_4210),
.B(n_306),
.Y(n_4274)
);

INVx2_ASAP7_75t_L g4275 ( 
.A(n_4235),
.Y(n_4275)
);

INVx2_ASAP7_75t_L g4276 ( 
.A(n_4234),
.Y(n_4276)
);

AOI22xp5_ASAP7_75t_L g4277 ( 
.A1(n_4227),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_L g4278 ( 
.A(n_4228),
.B(n_307),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4236),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_SL g4280 ( 
.A(n_4210),
.B(n_308),
.Y(n_4280)
);

AOI22xp5_ASAP7_75t_L g4281 ( 
.A1(n_4193),
.A2(n_309),
.B1(n_311),
.B2(n_313),
.Y(n_4281)
);

AND2x2_ASAP7_75t_L g4282 ( 
.A(n_4240),
.B(n_4204),
.Y(n_4282)
);

AND2x2_ASAP7_75t_L g4283 ( 
.A(n_4209),
.B(n_313),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_4188),
.B(n_315),
.Y(n_4284)
);

AOI221xp5_ASAP7_75t_L g4285 ( 
.A1(n_4192),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.C(n_319),
.Y(n_4285)
);

AOI21xp33_ASAP7_75t_L g4286 ( 
.A1(n_4194),
.A2(n_317),
.B(n_320),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_4244),
.Y(n_4287)
);

OAI22xp33_ASAP7_75t_L g4288 ( 
.A1(n_4219),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_4288)
);

AOI221xp5_ASAP7_75t_L g4289 ( 
.A1(n_4201),
.A2(n_322),
.B1(n_326),
.B2(n_327),
.C(n_328),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4216),
.Y(n_4290)
);

OAI31xp33_ASAP7_75t_L g4291 ( 
.A1(n_4243),
.A2(n_326),
.A3(n_328),
.B(n_329),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4220),
.Y(n_4292)
);

INVx3_ASAP7_75t_L g4293 ( 
.A(n_4246),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4238),
.Y(n_4294)
);

NAND2xp33_ASAP7_75t_L g4295 ( 
.A(n_4251),
.B(n_329),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_SL g4296 ( 
.A(n_4215),
.B(n_330),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_4233),
.B(n_330),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4241),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_L g4299 ( 
.A(n_4233),
.B(n_332),
.Y(n_4299)
);

AND2x2_ASAP7_75t_L g4300 ( 
.A(n_4250),
.B(n_334),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4245),
.Y(n_4301)
);

AOI221xp5_ASAP7_75t_L g4302 ( 
.A1(n_4231),
.A2(n_334),
.B1(n_335),
.B2(n_336),
.C(n_340),
.Y(n_4302)
);

NOR2xp33_ASAP7_75t_L g4303 ( 
.A(n_4293),
.B(n_4249),
.Y(n_4303)
);

O2A1O1Ixp33_ASAP7_75t_L g4304 ( 
.A1(n_4256),
.A2(n_4247),
.B(n_4208),
.C(n_4203),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_L g4305 ( 
.A(n_4293),
.B(n_4211),
.Y(n_4305)
);

HB1xp67_ASAP7_75t_L g4306 ( 
.A(n_4267),
.Y(n_4306)
);

NOR2xp33_ASAP7_75t_L g4307 ( 
.A(n_4269),
.B(n_4232),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_L g4308 ( 
.A(n_4256),
.B(n_4218),
.Y(n_4308)
);

OR2x2_ASAP7_75t_L g4309 ( 
.A(n_4267),
.B(n_4202),
.Y(n_4309)
);

NOR2xp33_ASAP7_75t_L g4310 ( 
.A(n_4255),
.B(n_4223),
.Y(n_4310)
);

NOR2xp33_ASAP7_75t_L g4311 ( 
.A(n_4273),
.B(n_4254),
.Y(n_4311)
);

O2A1O1Ixp33_ASAP7_75t_L g4312 ( 
.A1(n_4274),
.A2(n_4205),
.B(n_4221),
.C(n_4206),
.Y(n_4312)
);

HB1xp67_ASAP7_75t_L g4313 ( 
.A(n_4267),
.Y(n_4313)
);

OR2x2_ASAP7_75t_L g4314 ( 
.A(n_4257),
.B(n_4217),
.Y(n_4314)
);

NOR2xp33_ASAP7_75t_L g4315 ( 
.A(n_4268),
.B(n_4226),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4259),
.Y(n_4316)
);

OAI322xp33_ASAP7_75t_L g4317 ( 
.A1(n_4265),
.A2(n_336),
.A3(n_340),
.B1(n_341),
.B2(n_342),
.C1(n_343),
.C2(n_344),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_4276),
.B(n_341),
.Y(n_4318)
);

NOR3x1_ASAP7_75t_L g4319 ( 
.A(n_4263),
.B(n_342),
.C(n_343),
.Y(n_4319)
);

OAI21xp5_ASAP7_75t_L g4320 ( 
.A1(n_4266),
.A2(n_344),
.B(n_345),
.Y(n_4320)
);

OAI21xp5_ASAP7_75t_SL g4321 ( 
.A1(n_4252),
.A2(n_346),
.B(n_348),
.Y(n_4321)
);

NAND4xp25_ASAP7_75t_SL g4322 ( 
.A(n_4302),
.B(n_348),
.C(n_349),
.D(n_350),
.Y(n_4322)
);

AOI21xp5_ASAP7_75t_L g4323 ( 
.A1(n_4280),
.A2(n_350),
.B(n_351),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4283),
.Y(n_4324)
);

NOR3x1_ASAP7_75t_L g4325 ( 
.A(n_4272),
.B(n_352),
.C(n_353),
.Y(n_4325)
);

INVx1_ASAP7_75t_SL g4326 ( 
.A(n_4258),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4282),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4270),
.Y(n_4328)
);

NOR2xp33_ASAP7_75t_L g4329 ( 
.A(n_4253),
.B(n_4297),
.Y(n_4329)
);

AO22x1_ASAP7_75t_L g4330 ( 
.A1(n_4299),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_4330)
);

NOR2xp33_ASAP7_75t_L g4331 ( 
.A(n_4275),
.B(n_354),
.Y(n_4331)
);

NOR2xp33_ASAP7_75t_L g4332 ( 
.A(n_4279),
.B(n_356),
.Y(n_4332)
);

INVxp67_ASAP7_75t_SL g4333 ( 
.A(n_4295),
.Y(n_4333)
);

NAND3xp33_ASAP7_75t_L g4334 ( 
.A(n_4285),
.B(n_356),
.C(n_359),
.Y(n_4334)
);

XNOR2xp5_ASAP7_75t_L g4335 ( 
.A(n_4261),
.B(n_359),
.Y(n_4335)
);

AOI21xp5_ASAP7_75t_L g4336 ( 
.A1(n_4296),
.A2(n_360),
.B(n_361),
.Y(n_4336)
);

NOR3x1_ASAP7_75t_L g4337 ( 
.A(n_4278),
.B(n_4260),
.C(n_4301),
.Y(n_4337)
);

NOR3x1_ASAP7_75t_L g4338 ( 
.A(n_4284),
.B(n_362),
.C(n_363),
.Y(n_4338)
);

NOR2xp33_ASAP7_75t_L g4339 ( 
.A(n_4288),
.B(n_362),
.Y(n_4339)
);

NOR2xp67_ASAP7_75t_SL g4340 ( 
.A(n_4298),
.B(n_363),
.Y(n_4340)
);

NOR2xp33_ASAP7_75t_L g4341 ( 
.A(n_4306),
.B(n_4286),
.Y(n_4341)
);

OAI21xp5_ASAP7_75t_SL g4342 ( 
.A1(n_4326),
.A2(n_4264),
.B(n_4271),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4313),
.Y(n_4343)
);

AOI21xp5_ASAP7_75t_L g4344 ( 
.A1(n_4303),
.A2(n_4262),
.B(n_4289),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_4340),
.Y(n_4345)
);

NAND3xp33_ASAP7_75t_L g4346 ( 
.A(n_4311),
.B(n_4290),
.C(n_4292),
.Y(n_4346)
);

AOI221xp5_ASAP7_75t_L g4347 ( 
.A1(n_4312),
.A2(n_4294),
.B1(n_4287),
.B2(n_4300),
.C(n_4291),
.Y(n_4347)
);

OAI322xp33_ASAP7_75t_L g4348 ( 
.A1(n_4309),
.A2(n_4281),
.A3(n_4277),
.B1(n_4291),
.B2(n_368),
.C1(n_369),
.C2(n_370),
.Y(n_4348)
);

AOI221xp5_ASAP7_75t_L g4349 ( 
.A1(n_4304),
.A2(n_364),
.B1(n_366),
.B2(n_367),
.C(n_369),
.Y(n_4349)
);

OA211x2_ASAP7_75t_L g4350 ( 
.A1(n_4322),
.A2(n_371),
.B(n_372),
.C(n_373),
.Y(n_4350)
);

AOI221xp5_ASAP7_75t_L g4351 ( 
.A1(n_4329),
.A2(n_371),
.B1(n_373),
.B2(n_375),
.C(n_376),
.Y(n_4351)
);

NAND2xp5_ASAP7_75t_L g4352 ( 
.A(n_4330),
.B(n_377),
.Y(n_4352)
);

OAI32xp33_ASAP7_75t_L g4353 ( 
.A1(n_4308),
.A2(n_377),
.A3(n_379),
.B1(n_380),
.B2(n_381),
.Y(n_4353)
);

NOR2xp67_ASAP7_75t_L g4354 ( 
.A(n_4327),
.B(n_379),
.Y(n_4354)
);

A2O1A1Ixp33_ASAP7_75t_L g4355 ( 
.A1(n_4315),
.A2(n_381),
.B(n_382),
.C(n_383),
.Y(n_4355)
);

AOI222xp33_ASAP7_75t_L g4356 ( 
.A1(n_4333),
.A2(n_382),
.B1(n_383),
.B2(n_384),
.C1(n_385),
.C2(n_387),
.Y(n_4356)
);

AOI221xp5_ASAP7_75t_L g4357 ( 
.A1(n_4307),
.A2(n_384),
.B1(n_385),
.B2(n_388),
.C(n_389),
.Y(n_4357)
);

OAI21xp33_ASAP7_75t_SL g4358 ( 
.A1(n_4310),
.A2(n_390),
.B(n_391),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_SL g4359 ( 
.A(n_4323),
.B(n_4316),
.Y(n_4359)
);

AOI211xp5_ASAP7_75t_L g4360 ( 
.A1(n_4320),
.A2(n_390),
.B(n_391),
.C(n_392),
.Y(n_4360)
);

NOR2xp67_ASAP7_75t_L g4361 ( 
.A(n_4336),
.B(n_392),
.Y(n_4361)
);

OAI221xp5_ASAP7_75t_L g4362 ( 
.A1(n_4321),
.A2(n_393),
.B1(n_394),
.B2(n_395),
.C(n_396),
.Y(n_4362)
);

OAI21xp33_ASAP7_75t_L g4363 ( 
.A1(n_4305),
.A2(n_393),
.B(n_395),
.Y(n_4363)
);

NAND2xp5_ASAP7_75t_L g4364 ( 
.A(n_4332),
.B(n_397),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_SL g4365 ( 
.A(n_4354),
.B(n_4320),
.Y(n_4365)
);

O2A1O1Ixp33_ASAP7_75t_SL g4366 ( 
.A1(n_4352),
.A2(n_4318),
.B(n_4314),
.C(n_4324),
.Y(n_4366)
);

AOI222xp33_ASAP7_75t_L g4367 ( 
.A1(n_4343),
.A2(n_4328),
.B1(n_4334),
.B2(n_4339),
.C1(n_4335),
.C2(n_4331),
.Y(n_4367)
);

OAI21xp5_ASAP7_75t_L g4368 ( 
.A1(n_4346),
.A2(n_4358),
.B(n_4344),
.Y(n_4368)
);

AOI21x1_ASAP7_75t_L g4369 ( 
.A1(n_4359),
.A2(n_4338),
.B(n_4319),
.Y(n_4369)
);

O2A1O1Ixp33_ASAP7_75t_L g4370 ( 
.A1(n_4355),
.A2(n_4317),
.B(n_4325),
.C(n_4337),
.Y(n_4370)
);

AOI221xp5_ASAP7_75t_L g4371 ( 
.A1(n_4348),
.A2(n_397),
.B1(n_398),
.B2(n_399),
.C(n_400),
.Y(n_4371)
);

NAND3xp33_ASAP7_75t_L g4372 ( 
.A(n_4349),
.B(n_398),
.C(n_399),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_SL g4373 ( 
.A(n_4356),
.B(n_401),
.Y(n_4373)
);

OAI22xp5_ASAP7_75t_L g4374 ( 
.A1(n_4345),
.A2(n_401),
.B1(n_402),
.B2(n_403),
.Y(n_4374)
);

AOI221xp5_ASAP7_75t_L g4375 ( 
.A1(n_4347),
.A2(n_403),
.B1(n_404),
.B2(n_405),
.C(n_406),
.Y(n_4375)
);

AOI21xp5_ASAP7_75t_L g4376 ( 
.A1(n_4342),
.A2(n_405),
.B(n_406),
.Y(n_4376)
);

NAND2xp5_ASAP7_75t_L g4377 ( 
.A(n_4360),
.B(n_407),
.Y(n_4377)
);

NAND4xp25_ASAP7_75t_SL g4378 ( 
.A(n_4357),
.B(n_408),
.C(n_409),
.D(n_410),
.Y(n_4378)
);

NAND4xp25_ASAP7_75t_L g4379 ( 
.A(n_4341),
.B(n_409),
.C(n_411),
.D(n_412),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4350),
.Y(n_4380)
);

O2A1O1Ixp33_ASAP7_75t_L g4381 ( 
.A1(n_4365),
.A2(n_4353),
.B(n_4362),
.C(n_4364),
.Y(n_4381)
);

NAND4xp25_ASAP7_75t_SL g4382 ( 
.A(n_4371),
.B(n_4351),
.C(n_4361),
.D(n_4363),
.Y(n_4382)
);

NAND4xp25_ASAP7_75t_L g4383 ( 
.A(n_4367),
.B(n_414),
.C(n_415),
.D(n_416),
.Y(n_4383)
);

AOI211xp5_ASAP7_75t_L g4384 ( 
.A1(n_4378),
.A2(n_414),
.B(n_416),
.C(n_417),
.Y(n_4384)
);

NOR4xp25_ASAP7_75t_L g4385 ( 
.A(n_4370),
.B(n_418),
.C(n_419),
.D(n_421),
.Y(n_4385)
);

AOI22xp33_ASAP7_75t_SL g4386 ( 
.A1(n_4380),
.A2(n_419),
.B1(n_421),
.B2(n_422),
.Y(n_4386)
);

OAI221xp5_ASAP7_75t_L g4387 ( 
.A1(n_4368),
.A2(n_422),
.B1(n_423),
.B2(n_424),
.C(n_425),
.Y(n_4387)
);

O2A1O1Ixp33_ASAP7_75t_L g4388 ( 
.A1(n_4373),
.A2(n_424),
.B(n_427),
.C(n_428),
.Y(n_4388)
);

NOR4xp25_ASAP7_75t_L g4389 ( 
.A(n_4366),
.B(n_4375),
.C(n_4372),
.D(n_4377),
.Y(n_4389)
);

O2A1O1Ixp33_ASAP7_75t_L g4390 ( 
.A1(n_4376),
.A2(n_4374),
.B(n_4379),
.C(n_4369),
.Y(n_4390)
);

HB1xp67_ASAP7_75t_L g4391 ( 
.A(n_4369),
.Y(n_4391)
);

OR2x2_ASAP7_75t_L g4392 ( 
.A(n_4385),
.B(n_429),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_4391),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4388),
.Y(n_4394)
);

INVx2_ASAP7_75t_SL g4395 ( 
.A(n_4386),
.Y(n_4395)
);

NAND4xp25_ASAP7_75t_L g4396 ( 
.A(n_4381),
.B(n_430),
.C(n_431),
.D(n_432),
.Y(n_4396)
);

NAND2xp5_ASAP7_75t_L g4397 ( 
.A(n_4384),
.B(n_430),
.Y(n_4397)
);

NAND4xp75_ASAP7_75t_L g4398 ( 
.A(n_4383),
.B(n_431),
.C(n_433),
.D(n_434),
.Y(n_4398)
);

AOI21xp33_ASAP7_75t_SL g4399 ( 
.A1(n_4392),
.A2(n_4387),
.B(n_4390),
.Y(n_4399)
);

NOR2x1_ASAP7_75t_L g4400 ( 
.A(n_4396),
.B(n_4382),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_L g4401 ( 
.A(n_4393),
.B(n_4389),
.Y(n_4401)
);

NOR2xp33_ASAP7_75t_L g4402 ( 
.A(n_4398),
.B(n_434),
.Y(n_4402)
);

NAND4xp75_ASAP7_75t_L g4403 ( 
.A(n_4395),
.B(n_435),
.C(n_437),
.D(n_438),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4397),
.Y(n_4404)
);

NOR3xp33_ASAP7_75t_L g4405 ( 
.A(n_4399),
.B(n_4394),
.C(n_437),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_SL g4406 ( 
.A(n_4401),
.B(n_4402),
.Y(n_4406)
);

XNOR2x1_ASAP7_75t_L g4407 ( 
.A(n_4405),
.B(n_4400),
.Y(n_4407)
);

NOR2xp33_ASAP7_75t_R g4408 ( 
.A(n_4406),
.B(n_4404),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4407),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4409),
.Y(n_4410)
);

INVx2_ASAP7_75t_L g4411 ( 
.A(n_4410),
.Y(n_4411)
);

AND2x2_ASAP7_75t_L g4412 ( 
.A(n_4411),
.B(n_4408),
.Y(n_4412)
);

CKINVDCx14_ASAP7_75t_R g4413 ( 
.A(n_4412),
.Y(n_4413)
);

NAND2xp5_ASAP7_75t_L g4414 ( 
.A(n_4413),
.B(n_4403),
.Y(n_4414)
);

AOI22xp5_ASAP7_75t_L g4415 ( 
.A1(n_4414),
.A2(n_435),
.B1(n_439),
.B2(n_440),
.Y(n_4415)
);

AOI22xp5_ASAP7_75t_L g4416 ( 
.A1(n_4415),
.A2(n_440),
.B1(n_441),
.B2(n_442),
.Y(n_4416)
);

AOI31xp33_ASAP7_75t_L g4417 ( 
.A1(n_4416),
.A2(n_442),
.A3(n_443),
.B(n_444),
.Y(n_4417)
);

AOI322xp5_ASAP7_75t_L g4418 ( 
.A1(n_4417),
.A2(n_443),
.A3(n_445),
.B1(n_446),
.B2(n_450),
.C1(n_451),
.C2(n_452),
.Y(n_4418)
);

AOI221xp5_ASAP7_75t_L g4419 ( 
.A1(n_4418),
.A2(n_450),
.B1(n_452),
.B2(n_453),
.C(n_454),
.Y(n_4419)
);

AOI221xp5_ASAP7_75t_L g4420 ( 
.A1(n_4419),
.A2(n_1027),
.B1(n_1060),
.B2(n_1098),
.C(n_4393),
.Y(n_4420)
);

AOI211xp5_ASAP7_75t_L g4421 ( 
.A1(n_4420),
.A2(n_1098),
.B(n_1027),
.C(n_1060),
.Y(n_4421)
);


endmodule