module fake_jpeg_22491_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_1),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_46),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_22),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_25),
.B1(n_22),
.B2(n_31),
.Y(n_61)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

AO22x1_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_32),
.B1(n_29),
.B2(n_24),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_56),
.A2(n_26),
.B1(n_34),
.B2(n_24),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_59),
.B(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_62),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_61),
.A2(n_34),
.B1(n_26),
.B2(n_23),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_66),
.B(n_64),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_38),
.A2(n_31),
.B1(n_18),
.B2(n_20),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_68),
.A2(n_31),
.B1(n_22),
.B2(n_18),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_40),
.B(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_71),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_117)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_74),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_94),
.B1(n_99),
.B2(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_77),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_82),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_62),
.B(n_59),
.C(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_81),
.B(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_84),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_55),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_87),
.Y(n_128)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_56),
.A2(n_35),
.B(n_32),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_26),
.B(n_34),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_64),
.A2(n_19),
.B1(n_20),
.B2(n_30),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_93),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_54),
.A2(n_19),
.B1(n_30),
.B2(n_23),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_57),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_53),
.Y(n_107)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_101),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_102),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_61),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_24),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_110),
.B1(n_116),
.B2(n_125),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_89),
.Y(n_134)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_118),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_0),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_111),
.B(n_122),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_53),
.B1(n_67),
.B2(n_51),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_1),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_17),
.B(n_28),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_47),
.B(n_40),
.C(n_24),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_2),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_127),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_67),
.B1(n_17),
.B2(n_27),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_47),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_96),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_135),
.B(n_138),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_94),
.B1(n_82),
.B2(n_73),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_137),
.A2(n_117),
.B1(n_120),
.B2(n_115),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_94),
.B(n_89),
.C(n_73),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_139),
.B(n_147),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_117),
.A2(n_94),
.B1(n_76),
.B2(n_90),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_142),
.B(n_144),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_84),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_146),
.Y(n_187)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_94),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_87),
.B(n_28),
.C(n_27),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_156),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_122),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_111),
.Y(n_152)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_110),
.A2(n_116),
.B(n_125),
.C(n_113),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_135),
.B1(n_138),
.B2(n_133),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_113),
.B(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_160),
.Y(n_192)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_109),
.B(n_63),
.Y(n_161)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_110),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_162),
.A2(n_170),
.B(n_171),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_133),
.A2(n_130),
.B(n_126),
.Y(n_163)
);

NAND2xp33_ASAP7_75t_SL g220 ( 
.A(n_163),
.B(n_189),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_179),
.B1(n_184),
.B2(n_188),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_104),
.C(n_142),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_176),
.C(n_154),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_104),
.B(n_119),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_150),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_172),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_174),
.A2(n_190),
.B1(n_28),
.B2(n_27),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_128),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_2),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_115),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_128),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_17),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_140),
.A2(n_90),
.B1(n_112),
.B2(n_97),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_150),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_180),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_111),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_191),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_158),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_183),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_137),
.A2(n_139),
.B1(n_153),
.B2(n_147),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_78),
.B1(n_72),
.B2(n_88),
.Y(n_188)
);

NAND2xp33_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_111),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_149),
.B(n_144),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_134),
.A2(n_122),
.B(n_114),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_189),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_192),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_194),
.Y(n_249)
);

A2O1A1O1Ixp25_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_158),
.B(n_145),
.C(n_122),
.D(n_143),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_204),
.C(n_205),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_183),
.A2(n_157),
.B1(n_160),
.B2(n_156),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_196),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_250)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_221),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_114),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_199),
.B(n_209),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_206),
.A2(n_2),
.B(n_3),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_63),
.B1(n_141),
.B2(n_103),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_188),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_63),
.B1(n_49),
.B2(n_50),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_58),
.B1(n_52),
.B2(n_154),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_52),
.Y(n_212)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_28),
.Y(n_213)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_166),
.C(n_176),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_217),
.C(n_182),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_58),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_216),
.B(n_219),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_58),
.C(n_95),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_218),
.A2(n_180),
.B1(n_165),
.B2(n_173),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_164),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_167),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_178),
.B(n_11),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_222),
.B(n_223),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_178),
.B(n_11),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_198),
.A2(n_168),
.B(n_190),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_227),
.A2(n_229),
.B1(n_235),
.B2(n_241),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_174),
.Y(n_230)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_242),
.C(n_243),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_219),
.B(n_203),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_239),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_SL g235 ( 
.A1(n_203),
.A2(n_162),
.B(n_184),
.C(n_170),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_173),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_240),
.A2(n_247),
.B1(n_248),
.B2(n_197),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_202),
.A2(n_187),
.B1(n_162),
.B2(n_175),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_187),
.C(n_175),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_191),
.C(n_193),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_58),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_246),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_208),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_245),
.A2(n_217),
.B1(n_207),
.B2(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_213),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_205),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_254),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_200),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_267),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_198),
.C(n_204),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_259),
.C(n_260),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_195),
.C(n_202),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_220),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_211),
.B1(n_210),
.B2(n_206),
.Y(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_206),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_263),
.Y(n_281)
);

XNOR2x1_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_27),
.Y(n_264)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_264),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_95),
.B1(n_3),
.B2(n_4),
.Y(n_265)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_15),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_14),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_270),
.C(n_272),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_2),
.C(n_3),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_231),
.B(n_9),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_246),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_9),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_228),
.Y(n_280)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_285),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_234),
.C(n_240),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_288),
.C(n_290),
.Y(n_293)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_264),
.A2(n_233),
.B(n_249),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_279),
.B(n_280),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_248),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_251),
.B(n_247),
.C(n_237),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

OAI221xp5_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_226),
.B1(n_236),
.B2(n_272),
.C(n_261),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_249),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_235),
.Y(n_291)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_291),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_287),
.Y(n_292)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_292),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_250),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_274),
.B(n_260),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_13),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_259),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_296),
.B(n_273),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_276),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_301),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_258),
.C(n_270),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_299),
.C(n_305),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_254),
.C(n_228),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_278),
.A2(n_250),
.B1(n_237),
.B2(n_252),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_14),
.B(n_13),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_275),
.C(n_281),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_291),
.B(n_277),
.CI(n_273),
.CON(n_307),
.SN(n_307)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_5),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_313),
.C(n_317),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_293),
.A2(n_284),
.B(n_238),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_8),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_311),
.B(n_12),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_312),
.A2(n_316),
.B1(n_6),
.B2(n_8),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_302),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_11),
.Y(n_317)
);

AOI21x1_ASAP7_75t_L g318 ( 
.A1(n_292),
.A2(n_296),
.B(n_300),
.Y(n_318)
);

NOR3xp33_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_6),
.C(n_7),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_304),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_322),
.Y(n_329)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_326),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_325),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_314),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_317),
.Y(n_334)
);

AOI31xp67_ASAP7_75t_L g328 ( 
.A1(n_312),
.A2(n_307),
.A3(n_316),
.B(n_311),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_328),
.A2(n_315),
.B(n_306),
.Y(n_335)
);

OA21x2_ASAP7_75t_SL g331 ( 
.A1(n_320),
.A2(n_307),
.B(n_313),
.Y(n_331)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_331),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_325),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_335),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_330),
.Y(n_340)
);

A2O1A1Ixp33_ASAP7_75t_L g338 ( 
.A1(n_332),
.A2(n_321),
.B(n_331),
.C(n_329),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g341 ( 
.A(n_338),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_340),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_336),
.B(n_339),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_341),
.B(n_333),
.Y(n_344)
);


endmodule