module real_jpeg_4440_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_0),
.B(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_0),
.A2(n_43),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_0),
.B(n_136),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_0),
.B(n_322),
.C(n_325),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_L g327 ( 
.A1(n_0),
.A2(n_141),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_0),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_0),
.B(n_226),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_0),
.A2(n_47),
.B1(n_365),
.B2(n_373),
.Y(n_372)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_2),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_2),
.A2(n_57),
.B1(n_189),
.B2(n_192),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_2),
.A2(n_57),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g447 ( 
.A1(n_2),
.A2(n_57),
.B1(n_448),
.B2(n_449),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_3),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_3),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_3),
.A2(n_107),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_3),
.A2(n_107),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_3),
.A2(n_107),
.B1(n_115),
.B2(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_4),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_5),
.A2(n_115),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_5),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_133),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_5),
.A2(n_133),
.B1(n_340),
.B2(n_342),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_5),
.A2(n_133),
.B1(n_354),
.B2(n_355),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_6),
.A2(n_141),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_6),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_6),
.A2(n_48),
.B1(n_164),
.B2(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_6),
.A2(n_37),
.B1(n_164),
.B2(n_228),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_6),
.A2(n_164),
.B1(n_307),
.B2(n_309),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_7),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_66)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_7),
.A2(n_70),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_7),
.A2(n_70),
.B1(n_101),
.B2(n_296),
.Y(n_295)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_8),
.Y(n_180)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_8),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_8),
.Y(n_267)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_10),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_10),
.Y(n_127)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_10),
.Y(n_130)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_12),
.A2(n_96),
.B1(n_100),
.B2(n_101),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_12),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_12),
.A2(n_45),
.B1(n_100),
.B2(n_232),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_12),
.A2(n_49),
.B1(n_100),
.B2(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_12),
.A2(n_100),
.B1(n_203),
.B2(n_405),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_13),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_13),
.Y(n_121)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_13),
.Y(n_124)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_13),
.Y(n_135)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_13),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_13),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_13),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_14),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_14),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_14),
.A2(n_114),
.B1(n_252),
.B2(n_255),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_14),
.A2(n_114),
.B1(n_203),
.B2(n_331),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_14),
.A2(n_114),
.B1(n_366),
.B2(n_368),
.Y(n_365)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_15),
.Y(n_149)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_15),
.Y(n_152)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_15),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_433),
.Y(n_16)
);

OA21x2_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_311),
.B(n_427),
.Y(n_17)
);

NAND3xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_258),
.C(n_288),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_236),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_20),
.A2(n_429),
.B(n_430),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_194),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_21),
.B(n_194),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_138),
.C(n_175),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_22),
.B(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_74),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_23),
.B(n_75),
.C(n_111),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_46),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_24),
.B(n_46),
.Y(n_239)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.A3(n_32),
.B1(n_35),
.B2(n_42),
.Y(n_24)
);

INVx4_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_28),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_28),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g402 ( 
.A(n_28),
.Y(n_402)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_29),
.Y(n_254)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_30),
.Y(n_113)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g448 ( 
.A(n_31),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_34),
.A2(n_102),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp33_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_54),
.B1(n_62),
.B2(n_66),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_47),
.A2(n_66),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_47),
.B(n_182),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_47),
.A2(n_212),
.B(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_47),
.A2(n_210),
.B(n_347),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_47),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_47),
.A2(n_179),
.B1(n_353),
.B2(n_365),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_47),
.A2(n_177),
.B(n_212),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_53),
.Y(n_246)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_53),
.Y(n_377)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_55),
.A2(n_209),
.B(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_59),
.Y(n_348)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_61),
.Y(n_218)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_61),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_69),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_69),
.Y(n_214)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_71),
.Y(n_354)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_72),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_111),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_95),
.B(n_103),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_76),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_76),
.B(n_227),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_76),
.A2(n_226),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_76),
.A2(n_226),
.B1(n_251),
.B2(n_401),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_76),
.A2(n_295),
.B(n_443),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_86),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_77),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_171)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_77),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_77),
.A2(n_172),
.B1(n_173),
.B2(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_77),
.A2(n_275),
.B(n_278),
.Y(n_274)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_83),
.B2(n_85),
.Y(n_77)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_78),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_78),
.Y(n_329)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_79),
.Y(n_163)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_80),
.Y(n_396)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_82),
.Y(n_390)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_83),
.Y(n_202)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_84),
.Y(n_192)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_84),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_84),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_84),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_93),
.Y(n_86)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_90),
.Y(n_276)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI32xp33_ASAP7_75t_L g385 ( 
.A1(n_101),
.A2(n_386),
.A3(n_388),
.B1(n_391),
.B2(n_395),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_102),
.Y(n_229)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_102),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_104),
.A2(n_173),
.B(n_225),
.Y(n_224)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_105),
.Y(n_296)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_117),
.B1(n_131),
.B2(n_136),
.Y(n_111)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_117),
.A2(n_282),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_117),
.B(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_118),
.A2(n_137),
.B1(n_166),
.B2(n_170),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_118),
.A2(n_132),
.B1(n_137),
.B2(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_118),
.A2(n_231),
.B(n_281),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_128),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_129),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_135),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_136),
.B(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_137),
.B(n_306),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_137),
.A2(n_447),
.B(n_450),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_138),
.B(n_175),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_165),
.C(n_171),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g238 ( 
.A(n_139),
.B(n_165),
.CI(n_171),
.CON(n_238),
.SN(n_238)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_145),
.B(n_159),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_140),
.B(n_193),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_140),
.A2(n_145),
.B(n_193),
.Y(n_441)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_147)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_143),
.Y(n_397)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_145),
.A2(n_187),
.B1(n_188),
.B2(n_193),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_145),
.A2(n_159),
.B(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_145),
.B(n_187),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_145),
.A2(n_417),
.B(n_418),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_146),
.A2(n_160),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_146),
.A2(n_160),
.B1(n_327),
.B2(n_330),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_146),
.A2(n_160),
.B1(n_330),
.B2(n_339),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_146),
.A2(n_160),
.B1(n_339),
.B2(n_404),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_153),
.Y(n_146)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_148),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_150),
.B1(n_154),
.B2(n_157),
.Y(n_153)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_154),
.Y(n_325)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_167),
.Y(n_449)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_169),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_186),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_176),
.B(n_186),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

INVx3_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_180),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_189),
.Y(n_405)
);

INVx5_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_191),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_193),
.B(n_328),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_195),
.B(n_197),
.C(n_221),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_221),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_206),
.B2(n_207),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_198),
.B(n_207),
.Y(n_272)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_201),
.Y(n_269)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_219),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_218),
.Y(n_367)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_219),
.Y(n_373)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_235),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_230),
.B2(n_234),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_234),
.C(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_225),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_256),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_237),
.B(n_256),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.C(n_240),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_238),
.B(n_425),
.Y(n_424)
);

BUFx24_ASAP7_75t_SL g457 ( 
.A(n_238),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_239),
.B(n_240),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_247),
.C(n_249),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_241),
.A2(n_242),
.B1(n_247),
.B2(n_248),
.Y(n_412)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_249),
.B(n_412),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

A2O1A1O1Ixp25_ASAP7_75t_L g427 ( 
.A1(n_258),
.A2(n_288),
.B(n_428),
.C(n_431),
.D(n_432),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_287),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_259),
.B(n_287),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_263),
.C(n_286),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_271),
.B1(n_285),
.B2(n_286),
.Y(n_262)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_268),
.B2(n_270),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_264),
.A2(n_265),
.B1(n_304),
.B2(n_310),
.Y(n_303)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_268),
.Y(n_302)
);

AOI21xp33_ASAP7_75t_L g453 ( 
.A1(n_265),
.A2(n_302),
.B(n_304),
.Y(n_453)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_268),
.Y(n_270)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_279),
.C(n_284),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_279),
.B1(n_280),
.B2(n_284),
.Y(n_273)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_289),
.B(n_290),
.Y(n_432)
);

BUFx24_ASAP7_75t_SL g459 ( 
.A(n_290),
.Y(n_459)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_292),
.CI(n_301),
.CON(n_290),
.SN(n_290)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_291),
.B(n_292),
.C(n_301),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_297),
.B(n_300),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_293),
.B(n_297),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_298),
.Y(n_418)
);

FAx1_ASAP7_75t_SL g437 ( 
.A(n_300),
.B(n_438),
.CI(n_453),
.CON(n_437),
.SN(n_437)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_304),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_306),
.Y(n_451)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_422),
.B(n_426),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_313),
.A2(n_407),
.B(n_421),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_381),
.B(n_406),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_315),
.A2(n_349),
.B(n_380),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_334),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_316),
.B(n_334),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_326),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_317),
.B(n_326),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_321),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_328),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_328),
.B(n_392),
.Y(n_391)
);

OAI21xp33_ASAP7_75t_SL g401 ( 
.A1(n_328),
.A2(n_391),
.B(n_402),
.Y(n_401)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_333),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_346),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_338),
.B2(n_345),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_336),
.B(n_345),
.C(n_346),
.Y(n_382)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_338),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_347),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_361),
.B(n_379),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_360),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_351),
.B(n_360),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_352),
.A2(n_356),
.B1(n_357),
.B2(n_358),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_354),
.B(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_362),
.A2(n_371),
.B(n_378),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_363),
.B(n_364),
.Y(n_378)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx4_ASAP7_75t_SL g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_374),
.Y(n_371)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_382),
.B(n_383),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_399),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_384),
.B(n_400),
.C(n_403),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_385),
.B(n_398),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_385),
.B(n_398),
.Y(n_415)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx6_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_403),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_404),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_408),
.B(n_409),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_410),
.A2(n_411),
.B1(n_413),
.B2(n_414),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_410),
.B(n_416),
.C(n_419),
.Y(n_423)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_415),
.A2(n_416),
.B1(n_419),
.B2(n_420),
.Y(n_414)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_415),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_416),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_423),
.B(n_424),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_454),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_435),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_437),
.Y(n_455)
);

BUFx24_ASAP7_75t_SL g458 ( 
.A(n_437),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_439),
.A2(n_440),
.B1(n_446),
.B2(n_452),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_441),
.A2(n_442),
.B1(n_444),
.B2(n_445),
.Y(n_440)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_441),
.Y(n_445)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_442),
.Y(n_444)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_446),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);


endmodule