module fake_jpeg_32008_n_108 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_2),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_19),
.B(n_33),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_2),
.B(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_3),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_54),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_8),
.Y(n_78)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_44),
.B1(n_45),
.B2(n_39),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_75)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_45),
.B1(n_39),
.B2(n_42),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_71),
.B1(n_76),
.B2(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_45),
.B1(n_39),
.B2(n_36),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_74),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_41),
.B1(n_35),
.B2(n_20),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_77),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_23),
.B1(n_31),
.B2(n_9),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_7),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_79),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_8),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_83),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_86),
.Y(n_96)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_10),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_11),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_12),
.C(n_15),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_24),
.B(n_25),
.C(n_27),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_18),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_73),
.B1(n_71),
.B2(n_26),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_85),
.Y(n_100)
);

BUFx24_ASAP7_75t_SL g98 ( 
.A(n_95),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_96),
.B(n_85),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_93),
.C(n_92),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_97),
.B(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_102),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_87),
.Y(n_104)
);

OAI31xp33_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_84),
.A3(n_90),
.B(n_98),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_95),
.B(n_89),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_29),
.B(n_34),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_81),
.Y(n_108)
);


endmodule