module fake_ibex_958_n_2222 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_403, n_423, n_357, n_88, n_412, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_421, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_407, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_199, n_410, n_308, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_385, n_414, n_118, n_378, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_408, n_119, n_361, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_393, n_297, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_2222);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_407;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_410;
input n_308;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_118;
input n_378;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_393;
input n_297;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;

output n_2222;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_452;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_969;
wire n_678;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2151;
wire n_1391;
wire n_884;
wire n_667;
wire n_850;
wire n_1971;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_739;
wire n_853;
wire n_948;
wire n_504;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_641;
wire n_557;
wire n_1937;
wire n_893;
wire n_527;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_2163;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_554;
wire n_553;
wire n_2025;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2189;
wire n_745;
wire n_2112;
wire n_447;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_2203;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_1121;
wire n_693;
wire n_606;
wire n_737;
wire n_1571;
wire n_1980;
wire n_462;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2118;
wire n_2162;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2076;
wire n_974;
wire n_1036;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_1210;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2006;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2146;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1566;
wire n_1464;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_585;
wire n_1982;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_2142;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_2160;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_2094;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_1087;
wire n_757;
wire n_1599;
wire n_712;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_650;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_817;
wire n_2193;
wire n_2095;
wire n_555;
wire n_951;
wire n_2053;
wire n_468;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_2212;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_2170;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_2106;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1845;
wire n_1104;
wire n_1667;
wire n_1011;
wire n_2205;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2064;
wire n_1679;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_2110;
wire n_634;
wire n_961;
wire n_991;
wire n_1331;
wire n_1223;
wire n_1349;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_1353;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_1830;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2210;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2120;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_2108;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_1725;
wire n_2149;
wire n_1135;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_1270;
wire n_834;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_2182;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_1403;
wire n_2181;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_950;
wire n_512;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2078;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_1956;
wire n_681;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_1788;
wire n_2093;
wire n_786;
wire n_505;
wire n_2043;
wire n_1621;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2121;
wire n_1893;
wire n_1570;
wire n_701;
wire n_995;
wire n_1000;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1961;
wire n_1050;
wire n_2218;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_753;
wire n_2126;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_682;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_2131;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_755;
wire n_2091;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2079;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2092;
wire n_566;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_1902;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_SL g425 ( 
.A(n_309),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_287),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_95),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_212),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_41),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_339),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_408),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_18),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_348),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_9),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_390),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_265),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_243),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_420),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_92),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_255),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_84),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_355),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_92),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_27),
.Y(n_444)
);

NOR2xp67_ASAP7_75t_L g445 ( 
.A(n_73),
.B(n_299),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_18),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_47),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_111),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_170),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_377),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_6),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_417),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_402),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_55),
.Y(n_454)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_320),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_274),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_334),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_396),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_180),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_327),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_253),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_342),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_104),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_94),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_146),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_372),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_410),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_398),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_421),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_107),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_292),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_409),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_360),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_215),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_310),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_276),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_288),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_98),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_206),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_379),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_397),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_73),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_394),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_403),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_144),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_232),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_263),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_228),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_328),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_38),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_391),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_415),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_424),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_256),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_164),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_404),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_301),
.Y(n_497)
);

BUFx10_ASAP7_75t_L g498 ( 
.A(n_314),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_72),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_296),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_332),
.Y(n_501)
);

CKINVDCx14_ASAP7_75t_R g502 ( 
.A(n_182),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_165),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_69),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_133),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_78),
.B(n_313),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_87),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_172),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_105),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_54),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_216),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_59),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_381),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_151),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_343),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_290),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_152),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_338),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_225),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_412),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_145),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_113),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_347),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_325),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_285),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_278),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_130),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_388),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_128),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_244),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_201),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_380),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_80),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_60),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_55),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_16),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_61),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_335),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_53),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_89),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_352),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_393),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_366),
.B(n_139),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_392),
.Y(n_544)
);

BUFx5_ASAP7_75t_L g545 ( 
.A(n_341),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_411),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_371),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_87),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_384),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_340),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_228),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_158),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_257),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_96),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_200),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_374),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_272),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_385),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_167),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_172),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_399),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_315),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_368),
.Y(n_563)
);

BUFx5_ASAP7_75t_L g564 ( 
.A(n_229),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_209),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_82),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_103),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_364),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_386),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_R g570 ( 
.A(n_6),
.B(n_318),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_222),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_363),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_175),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_123),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_350),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_7),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_378),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_308),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_161),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_289),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_95),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_387),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_252),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_219),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_175),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_177),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_121),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_233),
.B(n_182),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_3),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_305),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_358),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_101),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_319),
.Y(n_593)
);

BUFx10_ASAP7_75t_L g594 ( 
.A(n_135),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_304),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_158),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_219),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_419),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_53),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_185),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_298),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_149),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_361),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_99),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_231),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_118),
.B(n_235),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_212),
.B(n_306),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_223),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_124),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_183),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_241),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_84),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_136),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_237),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_137),
.Y(n_615)
);

BUFx10_ASAP7_75t_L g616 ( 
.A(n_191),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_142),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_145),
.Y(n_618)
);

BUFx10_ASAP7_75t_L g619 ( 
.A(n_93),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_215),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_58),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_266),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_321),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_344),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_100),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_12),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_149),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_362),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_93),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_232),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_413),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_418),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_62),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_139),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_81),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_96),
.Y(n_636)
);

INVxp67_ASAP7_75t_SL g637 ( 
.A(n_259),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_337),
.B(n_142),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_74),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_354),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_41),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_200),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_204),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_203),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_316),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_382),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_189),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_25),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_191),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_365),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_163),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_65),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_359),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_69),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_357),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_159),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_239),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_423),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_311),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_275),
.Y(n_660)
);

NOR2xp67_ASAP7_75t_L g661 ( 
.A(n_227),
.B(n_356),
.Y(n_661)
);

NOR2xp67_ASAP7_75t_L g662 ( 
.A(n_121),
.B(n_242),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_221),
.Y(n_663)
);

BUFx5_ASAP7_75t_L g664 ( 
.A(n_256),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_414),
.Y(n_665)
);

CKINVDCx14_ASAP7_75t_R g666 ( 
.A(n_401),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_124),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_383),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_43),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_123),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_307),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_331),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_400),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_407),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_161),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_300),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_49),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_376),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_67),
.B(n_405),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_279),
.Y(n_680)
);

CKINVDCx16_ASAP7_75t_R g681 ( 
.A(n_416),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_277),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_43),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_266),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_49),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_3),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_196),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_324),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_260),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_395),
.Y(n_690)
);

BUFx10_ASAP7_75t_L g691 ( 
.A(n_138),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_295),
.Y(n_692)
);

INVxp67_ASAP7_75t_SL g693 ( 
.A(n_189),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_333),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_220),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_83),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_312),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_370),
.Y(n_698)
);

BUFx10_ASAP7_75t_L g699 ( 
.A(n_257),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_14),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_177),
.Y(n_701)
);

BUFx2_ASAP7_75t_L g702 ( 
.A(n_367),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_117),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_58),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_286),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_336),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_136),
.Y(n_707)
);

NOR2xp67_ASAP7_75t_L g708 ( 
.A(n_15),
.B(n_293),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_82),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_373),
.Y(n_710)
);

BUFx2_ASAP7_75t_SL g711 ( 
.A(n_389),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_197),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_70),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_406),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_101),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_422),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_194),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_79),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_178),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_61),
.B(n_157),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_179),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_375),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_369),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_271),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_230),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_450),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_598),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_439),
.B(n_0),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_601),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_435),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_564),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_502),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_502),
.B(n_0),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_SL g734 ( 
.A1(n_459),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_564),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_594),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_598),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_498),
.Y(n_738)
);

INVx4_ASAP7_75t_L g739 ( 
.A(n_498),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_467),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_702),
.B(n_4),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_439),
.B(n_503),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_503),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_566),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_566),
.Y(n_745)
);

BUFx12f_ASAP7_75t_L g746 ( 
.A(n_594),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_698),
.Y(n_747)
);

CKINVDCx6p67_ASAP7_75t_R g748 ( 
.A(n_498),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_698),
.Y(n_749)
);

BUFx12f_ASAP7_75t_L g750 ( 
.A(n_594),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_629),
.B(n_5),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_564),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_446),
.B(n_5),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_546),
.B(n_7),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_698),
.Y(n_755)
);

BUFx12f_ASAP7_75t_L g756 ( 
.A(n_605),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_698),
.Y(n_757)
);

BUFx8_ASAP7_75t_SL g758 ( 
.A(n_459),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_474),
.B(n_8),
.Y(n_759)
);

AOI22x1_ASAP7_75t_SL g760 ( 
.A1(n_478),
.A2(n_485),
.B1(n_488),
.B2(n_482),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_605),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_564),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_564),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_694),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_605),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_564),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_495),
.B(n_8),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_629),
.B(n_9),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_664),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_437),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_634),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_549),
.B(n_10),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_486),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_570),
.Y(n_774)
);

BUFx12f_ASAP7_75t_L g775 ( 
.A(n_616),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_634),
.Y(n_776)
);

BUFx12f_ASAP7_75t_L g777 ( 
.A(n_616),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_517),
.A2(n_13),
.B1(n_10),
.B2(n_11),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_694),
.Y(n_779)
);

OA21x2_ASAP7_75t_L g780 ( 
.A1(n_438),
.A2(n_516),
.B(n_473),
.Y(n_780)
);

AND2x6_ASAP7_75t_L g781 ( 
.A(n_438),
.B(n_282),
.Y(n_781)
);

BUFx12f_ASAP7_75t_L g782 ( 
.A(n_616),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_572),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_664),
.Y(n_784)
);

INVx5_ASAP7_75t_L g785 ( 
.A(n_582),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_508),
.B(n_11),
.Y(n_786)
);

INVx5_ASAP7_75t_L g787 ( 
.A(n_473),
.Y(n_787)
);

INVx5_ASAP7_75t_L g788 ( 
.A(n_516),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_675),
.B(n_13),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_510),
.B(n_14),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_576),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_675),
.B(n_15),
.Y(n_792)
);

INVx6_ASAP7_75t_L g793 ( 
.A(n_619),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_437),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_437),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_476),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_641),
.B(n_700),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_437),
.Y(n_798)
);

BUFx12f_ASAP7_75t_L g799 ( 
.A(n_619),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_707),
.B(n_16),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_531),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_696),
.Y(n_802)
);

BUFx8_ASAP7_75t_SL g803 ( 
.A(n_478),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_664),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_458),
.A2(n_20),
.B1(n_17),
.B2(n_19),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_SL g806 ( 
.A1(n_482),
.A2(n_488),
.B1(n_555),
.B2(n_485),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_696),
.B(n_17),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_427),
.B(n_19),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_531),
.Y(n_809)
);

BUFx8_ASAP7_75t_SL g810 ( 
.A(n_555),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_583),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_664),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_681),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_499),
.Y(n_814)
);

NOR2x1_ASAP7_75t_L g815 ( 
.A(n_499),
.B(n_283),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_724),
.Y(n_816)
);

OAI22x1_ASAP7_75t_SL g817 ( 
.A1(n_573),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_523),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_514),
.B(n_23),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_619),
.B(n_24),
.Y(n_820)
);

OAI22x1_ASAP7_75t_L g821 ( 
.A1(n_606),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_461),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_461),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_573),
.Y(n_824)
);

INVx5_ASAP7_75t_L g825 ( 
.A(n_523),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_545),
.B(n_26),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_428),
.B(n_27),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_463),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_537),
.Y(n_829)
);

INVx4_ASAP7_75t_L g830 ( 
.A(n_426),
.Y(n_830)
);

OAI22x1_ASAP7_75t_SL g831 ( 
.A1(n_581),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_545),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_587),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_537),
.B(n_28),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_463),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_548),
.Y(n_836)
);

BUFx8_ASAP7_75t_L g837 ( 
.A(n_506),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_769),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_819),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_731),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_735),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_819),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_834),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_SL g844 ( 
.A(n_733),
.B(n_458),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_728),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_728),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_752),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_751),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_762),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_751),
.Y(n_850)
);

OR2x6_ASAP7_75t_L g851 ( 
.A(n_746),
.B(n_662),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_763),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_766),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_738),
.B(n_558),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_832),
.B(n_580),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_784),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_793),
.Y(n_857)
);

OAI22xp33_ASAP7_75t_SL g858 ( 
.A1(n_805),
.A2(n_465),
.B1(n_579),
.B2(n_464),
.Y(n_858)
);

AND2x2_ASAP7_75t_SL g859 ( 
.A(n_768),
.B(n_543),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_730),
.B(n_464),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_804),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_768),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_812),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_739),
.B(n_645),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_780),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_730),
.B(n_732),
.Y(n_866)
);

INVxp67_ASAP7_75t_L g867 ( 
.A(n_823),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_732),
.B(n_465),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_780),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_793),
.Y(n_870)
);

INVx6_ASAP7_75t_L g871 ( 
.A(n_742),
.Y(n_871)
);

NAND2xp33_ASAP7_75t_SL g872 ( 
.A(n_739),
.B(n_471),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_787),
.B(n_674),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_796),
.B(n_811),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_789),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_789),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_793),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_822),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_758),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_740),
.B(n_783),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_792),
.Y(n_881)
);

CKINVDCx8_ASAP7_75t_R g882 ( 
.A(n_774),
.Y(n_882)
);

CKINVDCx16_ASAP7_75t_R g883 ( 
.A(n_750),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_726),
.Y(n_884)
);

OR2x2_ASAP7_75t_SL g885 ( 
.A(n_816),
.B(n_588),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_792),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_726),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_830),
.B(n_579),
.Y(n_888)
);

AOI21x1_ASAP7_75t_L g889 ( 
.A1(n_826),
.A2(n_815),
.B(n_433),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_807),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_787),
.B(n_545),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_822),
.Y(n_892)
);

INVxp33_ASAP7_75t_L g893 ( 
.A(n_828),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_758),
.Y(n_894)
);

OR2x6_ASAP7_75t_L g895 ( 
.A(n_756),
.B(n_711),
.Y(n_895)
);

INVxp67_ASAP7_75t_SL g896 ( 
.A(n_816),
.Y(n_896)
);

INVxp33_ASAP7_75t_SL g897 ( 
.A(n_828),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_787),
.B(n_545),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_835),
.Y(n_899)
);

NOR2x1p5_ASAP7_75t_L g900 ( 
.A(n_775),
.B(n_585),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_742),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_736),
.Y(n_902)
);

INVx8_ASAP7_75t_L g903 ( 
.A(n_777),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_807),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_743),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_744),
.Y(n_906)
);

CKINVDCx6p67_ASAP7_75t_R g907 ( 
.A(n_782),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_830),
.B(n_729),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_835),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_824),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_788),
.B(n_545),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_736),
.B(n_585),
.Y(n_912)
);

BUFx10_ASAP7_75t_L g913 ( 
.A(n_741),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_747),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_747),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_749),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_749),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_791),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_761),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_748),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_755),
.Y(n_921)
);

INVxp67_ASAP7_75t_SL g922 ( 
.A(n_773),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_755),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_755),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_761),
.B(n_765),
.Y(n_925)
);

INVx8_ASAP7_75t_L g926 ( 
.A(n_799),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_765),
.B(n_586),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_755),
.Y(n_928)
);

OAI22xp33_ASAP7_75t_SL g929 ( 
.A1(n_805),
.A2(n_701),
.B1(n_703),
.B2(n_586),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_773),
.B(n_455),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_745),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_771),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_757),
.Y(n_933)
);

BUFx10_ASAP7_75t_L g934 ( 
.A(n_741),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_757),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_757),
.Y(n_936)
);

INVx8_ASAP7_75t_L g937 ( 
.A(n_785),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_797),
.B(n_442),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_797),
.B(n_453),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_776),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_785),
.B(n_460),
.Y(n_941)
);

INVx5_ASAP7_75t_L g942 ( 
.A(n_781),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_770),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_802),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_803),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_759),
.Y(n_946)
);

XOR2xp5_ASAP7_75t_L g947 ( 
.A(n_824),
.B(n_471),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_803),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_820),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_770),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_770),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_759),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_767),
.Y(n_953)
);

AOI21x1_ASAP7_75t_L g954 ( 
.A1(n_814),
.A2(n_472),
.B(n_469),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_818),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_794),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_800),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_794),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_794),
.Y(n_959)
);

BUFx6f_ASAP7_75t_SL g960 ( 
.A(n_781),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_800),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_818),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_786),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_794),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_795),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_786),
.Y(n_966)
);

NOR2x1p5_ASAP7_75t_L g967 ( 
.A(n_810),
.B(n_701),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_753),
.Y(n_968)
);

OAI22xp33_ASAP7_75t_SL g969 ( 
.A1(n_813),
.A2(n_704),
.B1(n_703),
.B2(n_720),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_790),
.Y(n_970)
);

AND2x2_ASAP7_75t_SL g971 ( 
.A(n_754),
.B(n_638),
.Y(n_971)
);

NAND3xp33_ASAP7_75t_L g972 ( 
.A(n_790),
.B(n_704),
.C(n_712),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_785),
.B(n_475),
.Y(n_973)
);

INVx8_ASAP7_75t_L g974 ( 
.A(n_781),
.Y(n_974)
);

AO21x2_ASAP7_75t_L g975 ( 
.A1(n_808),
.A2(n_480),
.B(n_477),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_798),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_727),
.B(n_779),
.Y(n_977)
);

NOR2x1_ASAP7_75t_L g978 ( 
.A(n_754),
.B(n_481),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_798),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_798),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_788),
.B(n_493),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_737),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_829),
.B(n_470),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_801),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_836),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_764),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_801),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_788),
.B(n_500),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_825),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_764),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_772),
.B(n_548),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_801),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_801),
.Y(n_993)
);

AO21x2_ASAP7_75t_L g994 ( 
.A1(n_827),
.A2(n_518),
.B(n_501),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_809),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_809),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_810),
.Y(n_997)
);

INVx5_ASAP7_75t_L g998 ( 
.A(n_781),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_825),
.B(n_779),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_827),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_772),
.B(n_520),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_837),
.B(n_524),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_946),
.B(n_837),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_918),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_952),
.B(n_457),
.Y(n_1005)
);

BUFx8_ASAP7_75t_L g1006 ( 
.A(n_948),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_901),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_953),
.B(n_462),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_859),
.A2(n_561),
.B1(n_577),
.B2(n_496),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_1000),
.B(n_957),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_859),
.A2(n_922),
.B1(n_961),
.B2(n_896),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_930),
.B(n_462),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_963),
.B(n_466),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_866),
.B(n_908),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_903),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_878),
.B(n_466),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_892),
.B(n_468),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_966),
.B(n_970),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_903),
.Y(n_1019)
);

INVxp67_ASAP7_75t_SL g1020 ( 
.A(n_897),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_955),
.Y(n_1021)
);

OAI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_893),
.A2(n_778),
.B1(n_584),
.B2(n_608),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_938),
.B(n_655),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_938),
.B(n_655),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_939),
.B(n_692),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_971),
.B(n_692),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_871),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_971),
.B(n_845),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_854),
.B(n_705),
.Y(n_1029)
);

AOI221xp5_ASAP7_75t_L g1030 ( 
.A1(n_858),
.A2(n_821),
.B1(n_806),
.B2(n_831),
.C(n_817),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_871),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_848),
.B(n_430),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_903),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_850),
.A2(n_666),
.B1(n_429),
.B2(n_434),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_862),
.B(n_431),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_871),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_865),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_846),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_SL g1039 ( 
.A(n_895),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_864),
.B(n_452),
.Y(n_1040)
);

INVxp33_ASAP7_75t_L g1041 ( 
.A(n_874),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_SL g1042 ( 
.A(n_895),
.Y(n_1042)
);

NOR2x1p5_ASAP7_75t_L g1043 ( 
.A(n_907),
.B(n_760),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_860),
.B(n_483),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_846),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_962),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_985),
.Y(n_1047)
);

INVx1_ASAP7_75t_SL g1048 ( 
.A(n_899),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_888),
.B(n_484),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_905),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_919),
.B(n_425),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_906),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_919),
.B(n_491),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_978),
.B(n_968),
.Y(n_1054)
);

INVx4_ASAP7_75t_SL g1055 ( 
.A(n_960),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_949),
.A2(n_561),
.B1(n_577),
.B2(n_496),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_931),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_857),
.B(n_515),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_989),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_865),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_932),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_929),
.A2(n_443),
.B(n_448),
.C(n_432),
.Y(n_1062)
);

NOR2xp67_ASAP7_75t_L g1063 ( 
.A(n_867),
.B(n_607),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_885),
.A2(n_628),
.B1(n_653),
.B2(n_591),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_869),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_991),
.B(n_880),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_875),
.B(n_876),
.Y(n_1067)
);

AO221x1_ASAP7_75t_L g1068 ( 
.A1(n_909),
.A2(n_734),
.B1(n_591),
.B2(n_673),
.C(n_653),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_991),
.B(n_880),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_940),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_881),
.B(n_886),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_839),
.A2(n_673),
.B1(n_690),
.B2(n_628),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_944),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_890),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_974),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_904),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_842),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_843),
.A2(n_690),
.B1(n_584),
.B2(n_608),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_972),
.B(n_489),
.Y(n_1079)
);

NOR2xp67_ASAP7_75t_L g1080 ( 
.A(n_912),
.B(n_679),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_975),
.B(n_541),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_975),
.B(n_542),
.Y(n_1082)
);

NOR2x1p5_ASAP7_75t_L g1083 ( 
.A(n_879),
.B(n_894),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_870),
.B(n_578),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_927),
.B(n_492),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_877),
.B(n_650),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_994),
.B(n_544),
.Y(n_1087)
);

BUFx5_ASAP7_75t_L g1088 ( 
.A(n_902),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_868),
.B(n_697),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_925),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_1001),
.B(n_714),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_982),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_926),
.Y(n_1093)
);

AND2x6_ASAP7_75t_L g1094 ( 
.A(n_920),
.B(n_562),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_926),
.Y(n_1095)
);

NOR3xp33_ASAP7_75t_L g1096 ( 
.A(n_969),
.B(n_693),
.C(n_637),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_L g1097 ( 
.A(n_838),
.B(n_568),
.C(n_563),
.Y(n_1097)
);

BUFx5_ASAP7_75t_L g1098 ( 
.A(n_913),
.Y(n_1098)
);

AND2x4_ASAP7_75t_SL g1099 ( 
.A(n_895),
.B(n_691),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_913),
.B(n_497),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_986),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_R g1102 ( 
.A(n_883),
.B(n_581),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_983),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_934),
.B(n_691),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_990),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1002),
.A2(n_725),
.B1(n_721),
.B2(n_440),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_994),
.Y(n_1107)
);

NOR2xp67_ASAP7_75t_L g1108 ( 
.A(n_1002),
.B(n_30),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_934),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_851),
.B(n_716),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_977),
.B(n_513),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_977),
.B(n_525),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_937),
.B(n_528),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_851),
.B(n_532),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_SL g1115 ( 
.A(n_851),
.Y(n_1115)
);

AND3x1_ASAP7_75t_L g1116 ( 
.A(n_872),
.B(n_456),
.C(n_454),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_937),
.B(n_941),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_838),
.B(n_575),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_942),
.B(n_538),
.Y(n_1119)
);

AND2x2_ASAP7_75t_SL g1120 ( 
.A(n_882),
.B(n_633),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_900),
.B(n_699),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_937),
.B(n_547),
.Y(n_1122)
);

XOR2xp5_ASAP7_75t_L g1123 ( 
.A(n_947),
.B(n_627),
.Y(n_1123)
);

NOR3xp33_ASAP7_75t_L g1124 ( 
.A(n_844),
.B(n_617),
.C(n_505),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_967),
.B(n_699),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_840),
.B(n_593),
.Y(n_1126)
);

AO221x1_ASAP7_75t_L g1127 ( 
.A1(n_844),
.A2(n_643),
.B1(n_651),
.B2(n_644),
.C(n_627),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_974),
.B(n_550),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_954),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_889),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_942),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_941),
.B(n_556),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_945),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_973),
.B(n_841),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_942),
.Y(n_1135)
);

OR2x2_ASAP7_75t_L g1136 ( 
.A(n_997),
.B(n_620),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_981),
.B(n_569),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_855),
.A2(n_715),
.B1(n_717),
.B2(n_713),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_910),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_988),
.B(n_590),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_847),
.B(n_595),
.Y(n_1141)
);

OR2x6_ASAP7_75t_L g1142 ( 
.A(n_891),
.B(n_633),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_988),
.B(n_603),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_849),
.B(n_623),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_852),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_960),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_998),
.B(n_624),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_853),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_999),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_998),
.B(n_640),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_856),
.B(n_646),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_958),
.Y(n_1152)
);

BUFx5_ASAP7_75t_L g1153 ( 
.A(n_891),
.Y(n_1153)
);

INVxp33_ASAP7_75t_L g1154 ( 
.A(n_873),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_898),
.B(n_676),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_861),
.B(n_678),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_863),
.B(n_688),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_SL g1158 ( 
.A(n_863),
.B(n_706),
.Y(n_1158)
);

BUFx5_ASAP7_75t_L g1159 ( 
.A(n_911),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_911),
.B(n_710),
.Y(n_1160)
);

AND2x2_ASAP7_75t_SL g1161 ( 
.A(n_943),
.B(n_654),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_950),
.B(n_436),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_951),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_958),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_951),
.A2(n_479),
.B(n_490),
.C(n_487),
.Y(n_1165)
);

INVx8_ASAP7_75t_L g1166 ( 
.A(n_958),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_956),
.A2(n_444),
.B1(n_447),
.B2(n_441),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_956),
.B(n_449),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_959),
.B(n_451),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_884),
.B(n_631),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_884),
.B(n_632),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_964),
.B(n_699),
.Y(n_1172)
);

BUFx12f_ASAP7_75t_SL g1173 ( 
.A(n_984),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_965),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_923),
.B(n_658),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_887),
.B(n_659),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_923),
.B(n_665),
.Y(n_1177)
);

NOR3xp33_ASAP7_75t_L g1178 ( 
.A(n_976),
.B(n_504),
.C(n_494),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_933),
.B(n_668),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_933),
.B(n_671),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_933),
.B(n_672),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_984),
.Y(n_1182)
);

AND2x4_ASAP7_75t_SL g1183 ( 
.A(n_979),
.B(n_643),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_979),
.B(n_511),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_980),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_984),
.Y(n_1186)
);

INVxp33_ASAP7_75t_L g1187 ( 
.A(n_987),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_987),
.B(n_526),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_992),
.Y(n_1189)
);

NOR2xp67_ASAP7_75t_L g1190 ( 
.A(n_993),
.B(n_31),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_995),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1010),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1075),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1004),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1010),
.A2(n_723),
.B(n_722),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1018),
.A2(n_507),
.B(n_512),
.C(n_509),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1038),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1065),
.A2(n_661),
.B(n_445),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1158),
.B(n_534),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1003),
.B(n_644),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1014),
.B(n_536),
.Y(n_1201)
);

AOI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1129),
.A2(n_1107),
.B(n_1082),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1090),
.B(n_551),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1019),
.B(n_519),
.Y(n_1204)
);

NOR3xp33_ASAP7_75t_L g1205 ( 
.A(n_1030),
.B(n_554),
.C(n_552),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1066),
.B(n_557),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1045),
.Y(n_1207)
);

AND2x6_ASAP7_75t_SL g1208 ( 
.A(n_1123),
.B(n_651),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1081),
.A2(n_708),
.B(n_522),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1081),
.A2(n_527),
.B(n_521),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1048),
.B(n_652),
.Y(n_1211)
);

AO21x1_ASAP7_75t_L g1212 ( 
.A1(n_1082),
.A2(n_530),
.B(n_529),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1069),
.B(n_559),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1103),
.B(n_657),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1005),
.B(n_560),
.Y(n_1215)
);

INVx4_ASAP7_75t_L g1216 ( 
.A(n_1019),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1087),
.A2(n_1052),
.B(n_1057),
.C(n_1050),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1008),
.B(n_565),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1023),
.B(n_1024),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_SL g1220 ( 
.A1(n_1087),
.A2(n_535),
.B(n_539),
.C(n_533),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1134),
.A2(n_1071),
.B(n_1067),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1025),
.B(n_567),
.Y(n_1222)
);

BUFx4f_ASAP7_75t_L g1223 ( 
.A(n_1015),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1130),
.A2(n_553),
.B(n_540),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1013),
.B(n_571),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1013),
.B(n_574),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1074),
.B(n_589),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1093),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1076),
.B(n_597),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1012),
.A2(n_915),
.B(n_914),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1047),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1011),
.A2(n_695),
.B1(n_592),
.B2(n_599),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1080),
.B(n_1077),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1098),
.B(n_600),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1037),
.A2(n_917),
.B(n_916),
.Y(n_1235)
);

A2O1A1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1061),
.A2(n_596),
.B(n_615),
.C(n_613),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1028),
.A2(n_622),
.B(n_625),
.C(n_618),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1098),
.B(n_602),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1109),
.B(n_626),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1072),
.B(n_695),
.Y(n_1240)
);

OAI21xp33_ASAP7_75t_L g1241 ( 
.A1(n_1041),
.A2(n_609),
.B(n_604),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1098),
.B(n_610),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1063),
.B(n_1070),
.Y(n_1243)
);

INVxp67_ASAP7_75t_L g1244 ( 
.A(n_1095),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1073),
.B(n_611),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1089),
.B(n_1054),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1091),
.B(n_612),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1059),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1034),
.B(n_614),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1097),
.A2(n_636),
.B(n_630),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1088),
.B(n_1104),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1029),
.B(n_621),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1060),
.A2(n_924),
.B(n_921),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1046),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1009),
.A2(n_647),
.B1(n_649),
.B2(n_642),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1172),
.B(n_635),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1072),
.B(n_639),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1026),
.A2(n_1124),
.B1(n_1096),
.B2(n_1116),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1102),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1056),
.A2(n_667),
.B1(n_669),
.B2(n_663),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1016),
.B(n_648),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1007),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1097),
.A2(n_677),
.B(n_670),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1062),
.A2(n_682),
.B(n_689),
.C(n_680),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1060),
.A2(n_928),
.B(n_924),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1125),
.A2(n_656),
.B1(n_684),
.B2(n_683),
.Y(n_1266)
);

BUFx12f_ASAP7_75t_L g1267 ( 
.A(n_1006),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1027),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1017),
.B(n_685),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1022),
.A2(n_709),
.B(n_996),
.C(n_995),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1118),
.A2(n_936),
.B(n_935),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1044),
.B(n_686),
.Y(n_1272)
);

NOR2x1_ASAP7_75t_R g1273 ( 
.A(n_1133),
.B(n_718),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1078),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1033),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1165),
.A2(n_719),
.B(n_660),
.C(n_687),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1031),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1036),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1131),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1078),
.Y(n_1280)
);

NAND2x1p5_ASAP7_75t_L g1281 ( 
.A(n_1105),
.B(n_587),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1168),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1051),
.B(n_31),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1144),
.A2(n_833),
.B(n_284),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1126),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1053),
.B(n_32),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1064),
.A2(n_1126),
.B(n_1141),
.C(n_1079),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1131),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1021),
.Y(n_1289)
);

CKINVDCx20_ASAP7_75t_R g1290 ( 
.A(n_1139),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1121),
.B(n_34),
.Y(n_1291)
);

O2A1O1Ixp5_ASAP7_75t_L g1292 ( 
.A1(n_1085),
.A2(n_294),
.B(n_297),
.C(n_291),
.Y(n_1292)
);

OR2x2_ASAP7_75t_SL g1293 ( 
.A(n_1043),
.B(n_35),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1161),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1064),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1141),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1099),
.B(n_39),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1040),
.A2(n_44),
.B1(n_40),
.B2(n_42),
.Y(n_1298)
);

AO21x1_ASAP7_75t_L g1299 ( 
.A1(n_1179),
.A2(n_42),
.B(n_44),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1106),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1100),
.B(n_1032),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1035),
.B(n_46),
.Y(n_1302)
);

INVx8_ASAP7_75t_L g1303 ( 
.A(n_1039),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1049),
.B(n_48),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1183),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1146),
.B(n_50),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1156),
.A2(n_303),
.B(n_302),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1108),
.A2(n_54),
.B(n_51),
.C(n_52),
.Y(n_1308)
);

BUFx5_ASAP7_75t_L g1309 ( 
.A(n_1163),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1138),
.B(n_52),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1114),
.B(n_56),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1136),
.B(n_56),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1178),
.A2(n_63),
.B(n_57),
.C(n_62),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1039),
.A2(n_64),
.B1(n_57),
.B2(n_63),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1110),
.B(n_64),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1122),
.B(n_65),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1111),
.A2(n_322),
.B(n_317),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1092),
.B(n_66),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1101),
.B(n_66),
.Y(n_1319)
);

INVx6_ASAP7_75t_L g1320 ( 
.A(n_1083),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1112),
.A2(n_326),
.B(n_323),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1145),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1117),
.A2(n_330),
.B(n_329),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1094),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1170),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1120),
.B(n_68),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1148),
.B(n_71),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1171),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1055),
.B(n_72),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1171),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1176),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1094),
.Y(n_1332)
);

AO21x1_ASAP7_75t_L g1333 ( 
.A1(n_1181),
.A2(n_74),
.B(n_75),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1142),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1173),
.Y(n_1335)
);

AND2x6_ASAP7_75t_L g1336 ( 
.A(n_1055),
.B(n_345),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1154),
.B(n_79),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1068),
.B(n_80),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1055),
.B(n_83),
.Y(n_1339)
);

AND2x2_ASAP7_75t_SL g1340 ( 
.A(n_1042),
.B(n_85),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1128),
.B(n_86),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1167),
.B(n_86),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1160),
.A2(n_349),
.B(n_346),
.Y(n_1343)
);

AOI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1042),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1142),
.B(n_88),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1132),
.A2(n_353),
.B(n_351),
.Y(n_1346)
);

CKINVDCx11_ASAP7_75t_R g1347 ( 
.A(n_1115),
.Y(n_1347)
);

O2A1O1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1149),
.A2(n_94),
.B(n_90),
.C(n_91),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1153),
.B(n_91),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1162),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1058),
.B(n_97),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1084),
.B(n_97),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1169),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_SL g1354 ( 
.A(n_1153),
.B(n_98),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1086),
.B(n_100),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_1113),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1137),
.B(n_1140),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1159),
.B(n_102),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1143),
.B(n_102),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1115),
.B(n_103),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1151),
.B(n_105),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1184),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1188),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1155),
.B(n_106),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1157),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_1365)
);

OAI21xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1127),
.A2(n_108),
.B(n_109),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1135),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1119),
.B(n_1147),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1190),
.B(n_112),
.Y(n_1369)
);

INVx5_ASAP7_75t_L g1370 ( 
.A(n_1135),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1150),
.A2(n_1187),
.B(n_1177),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1135),
.B(n_114),
.Y(n_1372)
);

BUFx12f_ASAP7_75t_L g1373 ( 
.A(n_1164),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1175),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1182),
.B(n_115),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1166),
.B(n_116),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1180),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_1377)
);

AND2x2_ASAP7_75t_SL g1378 ( 
.A(n_1152),
.B(n_120),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1185),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1191),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1174),
.B(n_122),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1189),
.B(n_122),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1186),
.Y(n_1383)
);

O2A1O1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1010),
.A2(n_125),
.B(n_126),
.C(n_127),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1003),
.B(n_127),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1010),
.B(n_128),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1010),
.B(n_129),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1010),
.B(n_129),
.Y(n_1388)
);

NAND2x1p5_ASAP7_75t_L g1389 ( 
.A(n_1216),
.B(n_130),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1296),
.B(n_131),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1370),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1200),
.B(n_132),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1370),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1254),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1240),
.B(n_134),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1194),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1224),
.A2(n_134),
.B(n_135),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1211),
.B(n_138),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1231),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1244),
.Y(n_1400)
);

AO31x2_ASAP7_75t_L g1401 ( 
.A1(n_1212),
.A2(n_140),
.A3(n_141),
.B(n_143),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1224),
.A2(n_144),
.B(n_146),
.Y(n_1402)
);

NOR2xp67_ASAP7_75t_SL g1403 ( 
.A(n_1267),
.B(n_147),
.Y(n_1403)
);

AOI221xp5_ASAP7_75t_L g1404 ( 
.A1(n_1260),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.C(n_152),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1257),
.B(n_1274),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1271),
.A2(n_150),
.B(n_153),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1325),
.A2(n_1330),
.B(n_1328),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1331),
.A2(n_153),
.B(n_154),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1271),
.A2(n_155),
.B(n_156),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1214),
.B(n_157),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1350),
.B(n_159),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1353),
.B(n_160),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1280),
.B(n_162),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1362),
.B(n_163),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1282),
.B(n_1251),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1363),
.B(n_164),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1210),
.B(n_166),
.Y(n_1417)
);

INVx1_ASAP7_75t_SL g1418 ( 
.A(n_1204),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1357),
.A2(n_167),
.B(n_168),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1210),
.B(n_168),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1290),
.Y(n_1421)
);

INVx4_ASAP7_75t_L g1422 ( 
.A(n_1303),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1235),
.A2(n_169),
.B(n_170),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1246),
.B(n_171),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1386),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1370),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_SL g1427 ( 
.A(n_1223),
.B(n_1378),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1258),
.B(n_173),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1279),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1201),
.B(n_174),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1287),
.A2(n_1196),
.B(n_1385),
.C(n_1195),
.Y(n_1431)
);

AO31x2_ASAP7_75t_L g1432 ( 
.A1(n_1333),
.A2(n_176),
.A3(n_178),
.B(n_179),
.Y(n_1432)
);

AOI211x1_ASAP7_75t_L g1433 ( 
.A1(n_1209),
.A2(n_180),
.B(n_181),
.C(n_183),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1221),
.A2(n_1276),
.B(n_1387),
.Y(n_1434)
);

NOR2xp67_ASAP7_75t_L g1435 ( 
.A(n_1305),
.B(n_184),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1388),
.B(n_185),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1279),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1303),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1322),
.Y(n_1439)
);

CKINVDCx14_ASAP7_75t_R g1440 ( 
.A(n_1347),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1237),
.A2(n_186),
.B(n_187),
.C(n_188),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1253),
.A2(n_186),
.B(n_187),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1265),
.A2(n_188),
.B(n_190),
.Y(n_1443)
);

AOI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1255),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1345),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_1445)
);

O2A1O1Ixp5_ASAP7_75t_L g1446 ( 
.A1(n_1209),
.A2(n_195),
.B(n_198),
.C(n_199),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1239),
.B(n_198),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1233),
.A2(n_201),
.B(n_202),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1239),
.B(n_202),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1340),
.B(n_203),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1232),
.B(n_204),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1243),
.A2(n_205),
.B(n_206),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1250),
.A2(n_207),
.B(n_208),
.Y(n_1453)
);

O2A1O1Ixp5_ASAP7_75t_L g1454 ( 
.A1(n_1316),
.A2(n_207),
.B(n_208),
.C(n_210),
.Y(n_1454)
);

OAI22x1_ASAP7_75t_L g1455 ( 
.A1(n_1314),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1197),
.B(n_1207),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1262),
.Y(n_1457)
);

AND3x1_ASAP7_75t_L g1458 ( 
.A(n_1205),
.B(n_211),
.C(n_213),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1275),
.B(n_214),
.Y(n_1459)
);

OAI22x1_ASAP7_75t_L g1460 ( 
.A1(n_1344),
.A2(n_217),
.B1(n_218),
.B2(n_220),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1326),
.B(n_224),
.Y(n_1461)
);

NAND3xp33_ASAP7_75t_SL g1462 ( 
.A(n_1295),
.B(n_225),
.C(n_226),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1223),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1250),
.A2(n_227),
.B(n_229),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1373),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1203),
.B(n_230),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1225),
.A2(n_231),
.B(n_233),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1356),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1264),
.B(n_234),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1226),
.A2(n_236),
.B(n_237),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_1303),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1208),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1263),
.A2(n_238),
.B(n_239),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1263),
.A2(n_238),
.B(n_240),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1236),
.B(n_243),
.Y(n_1475)
);

BUFx12f_ASAP7_75t_L g1476 ( 
.A(n_1293),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1312),
.B(n_244),
.Y(n_1477)
);

BUFx12f_ASAP7_75t_L g1478 ( 
.A(n_1320),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1289),
.B(n_245),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1351),
.B(n_246),
.C(n_247),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1228),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1206),
.B(n_247),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1213),
.B(n_248),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1323),
.A2(n_248),
.B(n_249),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1248),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1291),
.B(n_249),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1245),
.B(n_250),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1335),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1218),
.A2(n_250),
.B(n_251),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1279),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1270),
.B(n_251),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1238),
.A2(n_252),
.B(n_253),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1320),
.B(n_281),
.Y(n_1493)
);

OAI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1317),
.A2(n_1321),
.B(n_1343),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1222),
.B(n_254),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1380),
.Y(n_1496)
);

OAI22x1_ASAP7_75t_L g1497 ( 
.A1(n_1259),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_1497)
);

AO31x2_ASAP7_75t_L g1498 ( 
.A1(n_1308),
.A2(n_261),
.A3(n_262),
.B(n_263),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1242),
.A2(n_264),
.B(n_265),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1304),
.B(n_267),
.Y(n_1500)
);

NAND3xp33_ASAP7_75t_SL g1501 ( 
.A(n_1300),
.B(n_268),
.C(n_269),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1227),
.B(n_270),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1342),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_1503)
);

INVx6_ASAP7_75t_L g1504 ( 
.A(n_1339),
.Y(n_1504)
);

BUFx6f_ASAP7_75t_L g1505 ( 
.A(n_1288),
.Y(n_1505)
);

A2O1A1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1352),
.A2(n_273),
.B(n_274),
.C(n_275),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1229),
.B(n_273),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1266),
.B(n_278),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1272),
.A2(n_279),
.B(n_280),
.Y(n_1509)
);

NOR2x1_ASAP7_75t_SL g1510 ( 
.A(n_1332),
.B(n_1288),
.Y(n_1510)
);

NAND2x1p5_ASAP7_75t_L g1511 ( 
.A(n_1324),
.B(n_1193),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1311),
.B(n_1220),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1341),
.A2(n_1283),
.B1(n_1286),
.B2(n_1359),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1379),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1247),
.B(n_1252),
.Y(n_1515)
);

OAI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1307),
.A2(n_1346),
.B(n_1284),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1256),
.B(n_1301),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1215),
.B(n_1249),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1355),
.A2(n_1337),
.B1(n_1261),
.B2(n_1269),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1234),
.A2(n_1371),
.B(n_1230),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1315),
.B(n_1302),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1360),
.Y(n_1522)
);

OR2x6_ASAP7_75t_L g1523 ( 
.A(n_1281),
.B(n_1329),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1310),
.A2(n_1292),
.B(n_1327),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1318),
.B(n_1319),
.Y(n_1525)
);

BUFx12f_ASAP7_75t_L g1526 ( 
.A(n_1336),
.Y(n_1526)
);

OA22x2_ASAP7_75t_L g1527 ( 
.A1(n_1338),
.A2(n_1306),
.B1(n_1241),
.B2(n_1294),
.Y(n_1527)
);

A2O1A1Ixp33_ASAP7_75t_L g1528 ( 
.A1(n_1348),
.A2(n_1384),
.B(n_1361),
.C(n_1364),
.Y(n_1528)
);

NOR2xp67_ASAP7_75t_L g1529 ( 
.A(n_1366),
.B(n_1297),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1309),
.B(n_1278),
.Y(n_1530)
);

AOI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1349),
.A2(n_1354),
.B(n_1358),
.Y(n_1531)
);

O2A1O1Ixp33_ASAP7_75t_SL g1532 ( 
.A1(n_1381),
.A2(n_1382),
.B(n_1369),
.C(n_1199),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1309),
.B(n_1277),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1268),
.Y(n_1534)
);

AOI21xp33_ASAP7_75t_L g1535 ( 
.A1(n_1375),
.A2(n_1376),
.B(n_1198),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_SL g1536 ( 
.A1(n_1334),
.A2(n_1298),
.B(n_1377),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1365),
.Y(n_1537)
);

OAI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1285),
.A2(n_1374),
.B(n_1372),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_SL g1539 ( 
.A(n_1273),
.B(n_1367),
.Y(n_1539)
);

BUFx12f_ASAP7_75t_L g1540 ( 
.A(n_1368),
.Y(n_1540)
);

INVx8_ASAP7_75t_L g1541 ( 
.A(n_1367),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1542)
);

NAND3xp33_ASAP7_75t_SL g1543 ( 
.A(n_1194),
.B(n_1102),
.C(n_1004),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1223),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1192),
.B(n_1004),
.Y(n_1545)
);

NOR3xp33_ASAP7_75t_L g1546 ( 
.A(n_1366),
.B(n_1200),
.C(n_1020),
.Y(n_1546)
);

OAI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1217),
.A2(n_1107),
.B(n_1202),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1200),
.B(n_1020),
.Y(n_1549)
);

AOI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1192),
.A2(n_1072),
.B1(n_1020),
.B2(n_1004),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1217),
.A2(n_1107),
.B(n_1202),
.Y(n_1553)
);

AO31x2_ASAP7_75t_L g1554 ( 
.A1(n_1212),
.A2(n_1217),
.A3(n_1333),
.B(n_1299),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1555)
);

CKINVDCx16_ASAP7_75t_R g1556 ( 
.A(n_1267),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1557)
);

NAND2x1p5_ASAP7_75t_L g1558 ( 
.A(n_1216),
.B(n_1192),
.Y(n_1558)
);

INVxp67_ASAP7_75t_SL g1559 ( 
.A(n_1192),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1192),
.B(n_1004),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1217),
.A2(n_1107),
.B(n_1202),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1192),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1563)
);

OAI22x1_ASAP7_75t_L g1564 ( 
.A1(n_1240),
.A2(n_947),
.B1(n_1056),
.B2(n_1009),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1192),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1267),
.Y(n_1570)
);

BUFx12f_ASAP7_75t_L g1571 ( 
.A(n_1267),
.Y(n_1571)
);

OAI22x1_ASAP7_75t_L g1572 ( 
.A1(n_1240),
.A2(n_947),
.B1(n_1056),
.B2(n_1009),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1192),
.B(n_1004),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1383),
.Y(n_1574)
);

INVxp67_ASAP7_75t_SL g1575 ( 
.A(n_1192),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1383),
.Y(n_1576)
);

AOI21xp33_ASAP7_75t_L g1577 ( 
.A1(n_1287),
.A2(n_1313),
.B(n_1286),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1192),
.B(n_1004),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1192),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1194),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1584)
);

NAND2x1p5_ASAP7_75t_L g1585 ( 
.A(n_1216),
.B(n_1192),
.Y(n_1585)
);

NOR2x1_ASAP7_75t_SL g1586 ( 
.A(n_1192),
.B(n_1216),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1194),
.Y(n_1587)
);

BUFx12f_ASAP7_75t_L g1588 ( 
.A(n_1267),
.Y(n_1588)
);

OAI22x1_ASAP7_75t_L g1589 ( 
.A1(n_1240),
.A2(n_947),
.B1(n_1056),
.B2(n_1009),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1590)
);

NOR2x1_ASAP7_75t_SL g1591 ( 
.A(n_1192),
.B(n_1216),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1200),
.B(n_1020),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1267),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_1267),
.Y(n_1594)
);

NOR2xp67_ASAP7_75t_L g1595 ( 
.A(n_1267),
.B(n_1019),
.Y(n_1595)
);

AND3x2_ASAP7_75t_L g1596 ( 
.A(n_1240),
.B(n_948),
.C(n_1004),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1192),
.B(n_1004),
.Y(n_1597)
);

OAI22x1_ASAP7_75t_L g1598 ( 
.A1(n_1240),
.A2(n_947),
.B1(n_1056),
.B2(n_1009),
.Y(n_1598)
);

INVx3_ASAP7_75t_SL g1599 ( 
.A(n_1194),
.Y(n_1599)
);

INVx2_ASAP7_75t_SL g1600 ( 
.A(n_1223),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1192),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1192),
.B(n_1004),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1603)
);

AO31x2_ASAP7_75t_L g1604 ( 
.A1(n_1212),
.A2(n_1217),
.A3(n_1333),
.B(n_1299),
.Y(n_1604)
);

AOI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1260),
.A2(n_858),
.B1(n_929),
.B2(n_969),
.C(n_1022),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1606)
);

NAND3xp33_ASAP7_75t_L g1607 ( 
.A(n_1200),
.B(n_837),
.C(n_1002),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1609)
);

NAND2x1p5_ASAP7_75t_L g1610 ( 
.A(n_1216),
.B(n_1192),
.Y(n_1610)
);

OAI21xp33_ASAP7_75t_SL g1611 ( 
.A1(n_1192),
.A2(n_1378),
.B(n_1296),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1192),
.B(n_1010),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1192),
.B(n_1004),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1192),
.B(n_1004),
.Y(n_1614)
);

NOR2xp67_ASAP7_75t_L g1615 ( 
.A(n_1422),
.B(n_1438),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1542),
.A2(n_1551),
.B(n_1548),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1562),
.A2(n_1575),
.B1(n_1559),
.B2(n_1548),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1545),
.B(n_1573),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1578),
.B(n_1597),
.Y(n_1619)
);

AO21x2_ASAP7_75t_L g1620 ( 
.A1(n_1547),
.A2(n_1561),
.B(n_1553),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1557),
.B(n_1569),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1569),
.B(n_1580),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1558),
.Y(n_1623)
);

BUFx10_ASAP7_75t_L g1624 ( 
.A(n_1593),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1599),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1602),
.B(n_1613),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1585),
.Y(n_1627)
);

BUFx12f_ASAP7_75t_L g1628 ( 
.A(n_1571),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1405),
.A2(n_1546),
.B1(n_1581),
.B2(n_1572),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1581),
.B(n_1551),
.Y(n_1630)
);

INVx8_ASAP7_75t_L g1631 ( 
.A(n_1588),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1585),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_L g1633 ( 
.A(n_1433),
.B(n_1519),
.C(n_1607),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1555),
.B(n_1582),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1582),
.Y(n_1635)
);

BUFx2_ASAP7_75t_R g1636 ( 
.A(n_1570),
.Y(n_1636)
);

OAI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1431),
.A2(n_1528),
.B(n_1515),
.Y(n_1637)
);

BUFx2_ASAP7_75t_SL g1638 ( 
.A(n_1595),
.Y(n_1638)
);

INVx3_ASAP7_75t_L g1639 ( 
.A(n_1610),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1584),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1610),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1590),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1391),
.Y(n_1643)
);

CKINVDCx11_ASAP7_75t_R g1644 ( 
.A(n_1556),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1515),
.A2(n_1603),
.B(n_1590),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1603),
.B(n_1606),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1606),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1612),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1612),
.B(n_1552),
.Y(n_1649)
);

NAND2x1p5_ASAP7_75t_L g1650 ( 
.A(n_1562),
.B(n_1422),
.Y(n_1650)
);

BUFx2_ASAP7_75t_SL g1651 ( 
.A(n_1594),
.Y(n_1651)
);

NAND2x1p5_ASAP7_75t_L g1652 ( 
.A(n_1438),
.B(n_1391),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1550),
.B(n_1549),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1393),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1563),
.B(n_1566),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1471),
.Y(n_1656)
);

NAND2x1p5_ASAP7_75t_L g1657 ( 
.A(n_1393),
.B(n_1426),
.Y(n_1657)
);

AO21x2_ASAP7_75t_L g1658 ( 
.A1(n_1577),
.A2(n_1524),
.B(n_1434),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1567),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1568),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1516),
.A2(n_1520),
.B(n_1494),
.Y(n_1661)
);

CKINVDCx16_ASAP7_75t_R g1662 ( 
.A(n_1440),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1608),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1614),
.B(n_1609),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1592),
.B(n_1418),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_L g1666 ( 
.A(n_1454),
.B(n_1446),
.C(n_1480),
.Y(n_1666)
);

NOR2xp67_ASAP7_75t_L g1667 ( 
.A(n_1543),
.B(n_1478),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1394),
.Y(n_1668)
);

BUFx2_ASAP7_75t_SL g1669 ( 
.A(n_1463),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1565),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1407),
.B(n_1586),
.Y(n_1671)
);

BUFx12f_ASAP7_75t_L g1672 ( 
.A(n_1421),
.Y(n_1672)
);

OAI21x1_ASAP7_75t_L g1673 ( 
.A1(n_1531),
.A2(n_1409),
.B(n_1406),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1396),
.Y(n_1674)
);

AO21x2_ASAP7_75t_L g1675 ( 
.A1(n_1535),
.A2(n_1538),
.B(n_1484),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1407),
.B(n_1591),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1601),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_L g1678 ( 
.A(n_1392),
.B(n_1513),
.C(n_1611),
.Y(n_1678)
);

CKINVDCx11_ASAP7_75t_R g1679 ( 
.A(n_1493),
.Y(n_1679)
);

INVxp67_ASAP7_75t_SL g1680 ( 
.A(n_1416),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1418),
.Y(n_1681)
);

INVx5_ASAP7_75t_L g1682 ( 
.A(n_1526),
.Y(n_1682)
);

OAI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1517),
.A2(n_1518),
.B(n_1521),
.Y(n_1683)
);

BUFx12f_ASAP7_75t_L g1684 ( 
.A(n_1465),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1457),
.Y(n_1685)
);

OA21x2_ASAP7_75t_L g1686 ( 
.A1(n_1423),
.A2(n_1443),
.B(n_1442),
.Y(n_1686)
);

OA21x2_ASAP7_75t_L g1687 ( 
.A1(n_1408),
.A2(n_1402),
.B(n_1397),
.Y(n_1687)
);

AO21x2_ASAP7_75t_L g1688 ( 
.A1(n_1512),
.A2(n_1408),
.B(n_1436),
.Y(n_1688)
);

BUFx4f_ASAP7_75t_L g1689 ( 
.A(n_1493),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1579),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1395),
.B(n_1605),
.Y(n_1691)
);

AO21x2_ASAP7_75t_L g1692 ( 
.A1(n_1512),
.A2(n_1436),
.B(n_1402),
.Y(n_1692)
);

OA21x2_ASAP7_75t_L g1693 ( 
.A1(n_1397),
.A2(n_1464),
.B(n_1453),
.Y(n_1693)
);

INVxp67_ASAP7_75t_SL g1694 ( 
.A(n_1416),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1564),
.A2(n_1598),
.B1(n_1589),
.B2(n_1537),
.Y(n_1695)
);

CKINVDCx20_ASAP7_75t_R g1696 ( 
.A(n_1583),
.Y(n_1696)
);

INVx3_ASAP7_75t_SL g1697 ( 
.A(n_1493),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1514),
.Y(n_1698)
);

INVx2_ASAP7_75t_SL g1699 ( 
.A(n_1504),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1456),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1461),
.B(n_1413),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1411),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1504),
.A2(n_1449),
.B1(n_1427),
.B2(n_1424),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1587),
.B(n_1400),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1425),
.B(n_1415),
.Y(n_1705)
);

INVx4_ASAP7_75t_L g1706 ( 
.A(n_1541),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1496),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1411),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1450),
.B(n_1449),
.Y(n_1709)
);

CKINVDCx6p67_ASAP7_75t_R g1710 ( 
.A(n_1476),
.Y(n_1710)
);

AOI22x1_ASAP7_75t_L g1711 ( 
.A1(n_1489),
.A2(n_1509),
.B1(n_1467),
.B2(n_1470),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1412),
.Y(n_1712)
);

AOI22x1_ASAP7_75t_L g1713 ( 
.A1(n_1492),
.A2(n_1499),
.B1(n_1389),
.B2(n_1419),
.Y(n_1713)
);

OA21x2_ASAP7_75t_L g1714 ( 
.A1(n_1453),
.A2(n_1474),
.B(n_1473),
.Y(n_1714)
);

CKINVDCx14_ASAP7_75t_R g1715 ( 
.A(n_1472),
.Y(n_1715)
);

OAI21x1_ASAP7_75t_L g1716 ( 
.A1(n_1530),
.A2(n_1533),
.B(n_1511),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1398),
.B(n_1477),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1560),
.B(n_1410),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1451),
.B(n_1508),
.Y(n_1719)
);

OAI221xp5_ASAP7_75t_SL g1720 ( 
.A1(n_1536),
.A2(n_1468),
.B1(n_1444),
.B2(n_1458),
.C(n_1404),
.Y(n_1720)
);

AO21x2_ASAP7_75t_L g1721 ( 
.A1(n_1417),
.A2(n_1420),
.B(n_1500),
.Y(n_1721)
);

INVx6_ASAP7_75t_L g1722 ( 
.A(n_1541),
.Y(n_1722)
);

OA21x2_ASAP7_75t_L g1723 ( 
.A1(n_1464),
.A2(n_1474),
.B(n_1473),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1412),
.Y(n_1724)
);

NOR2x1_ASAP7_75t_SL g1725 ( 
.A(n_1523),
.B(n_1429),
.Y(n_1725)
);

CKINVDCx20_ASAP7_75t_R g1726 ( 
.A(n_1481),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1439),
.Y(n_1727)
);

BUFx12f_ASAP7_75t_L g1728 ( 
.A(n_1540),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1399),
.B(n_1485),
.Y(n_1729)
);

CKINVDCx16_ASAP7_75t_R g1730 ( 
.A(n_1539),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1488),
.B(n_1414),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1479),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1525),
.A2(n_1532),
.B(n_1430),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1429),
.B(n_1437),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1536),
.B(n_1525),
.Y(n_1735)
);

NAND3xp33_ASAP7_75t_L g1736 ( 
.A(n_1506),
.B(n_1503),
.C(n_1441),
.Y(n_1736)
);

CKINVDCx11_ASAP7_75t_R g1737 ( 
.A(n_1459),
.Y(n_1737)
);

BUFx2_ASAP7_75t_L g1738 ( 
.A(n_1389),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1534),
.Y(n_1739)
);

BUFx8_ASAP7_75t_L g1740 ( 
.A(n_1544),
.Y(n_1740)
);

AO21x2_ASAP7_75t_L g1741 ( 
.A1(n_1491),
.A2(n_1462),
.B(n_1501),
.Y(n_1741)
);

BUFx10_ASAP7_75t_L g1742 ( 
.A(n_1459),
.Y(n_1742)
);

AO31x2_ASAP7_75t_L g1743 ( 
.A1(n_1445),
.A2(n_1475),
.A3(n_1469),
.B(n_1428),
.Y(n_1743)
);

OAI21x1_ASAP7_75t_SL g1744 ( 
.A1(n_1510),
.A2(n_1445),
.B(n_1475),
.Y(n_1744)
);

OAI21x1_ASAP7_75t_L g1745 ( 
.A1(n_1527),
.A2(n_1390),
.B(n_1487),
.Y(n_1745)
);

OAI21x1_ASAP7_75t_L g1746 ( 
.A1(n_1502),
.A2(n_1507),
.B(n_1495),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1466),
.B(n_1529),
.Y(n_1747)
);

OAI21x1_ASAP7_75t_L g1748 ( 
.A1(n_1495),
.A2(n_1483),
.B(n_1482),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1482),
.B(n_1483),
.Y(n_1749)
);

INVx5_ASAP7_75t_L g1750 ( 
.A(n_1490),
.Y(n_1750)
);

BUFx2_ASAP7_75t_SL g1751 ( 
.A(n_1600),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1574),
.Y(n_1752)
);

INVxp33_ASAP7_75t_L g1753 ( 
.A(n_1539),
.Y(n_1753)
);

AOI22x1_ASAP7_75t_L g1754 ( 
.A1(n_1455),
.A2(n_1460),
.B1(n_1452),
.B2(n_1448),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1447),
.Y(n_1755)
);

AO21x2_ASAP7_75t_L g1756 ( 
.A1(n_1486),
.A2(n_1469),
.B(n_1604),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1505),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1576),
.Y(n_1758)
);

NOR2x1_ASAP7_75t_SL g1759 ( 
.A(n_1523),
.B(n_1505),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_1596),
.Y(n_1760)
);

AOI21x1_ASAP7_75t_L g1761 ( 
.A1(n_1523),
.A2(n_1435),
.B(n_1497),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1401),
.Y(n_1762)
);

BUFx8_ASAP7_75t_L g1763 ( 
.A(n_1505),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1522),
.A2(n_1403),
.B1(n_1554),
.B2(n_1498),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1432),
.Y(n_1765)
);

INVx4_ASAP7_75t_L g1766 ( 
.A(n_1571),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1405),
.A2(n_1127),
.B1(n_1280),
.B2(n_1274),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1557),
.B(n_1569),
.Y(n_1768)
);

AOI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1542),
.A2(n_1551),
.B(n_1548),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1550),
.B(n_1274),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1550),
.B(n_1274),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1542),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1550),
.B(n_1274),
.Y(n_1773)
);

OAI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1431),
.A2(n_1528),
.B(n_1219),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1545),
.B(n_1004),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1571),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1599),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_L g1778 ( 
.A(n_1546),
.B(n_1433),
.C(n_1519),
.Y(n_1778)
);

INVx1_ASAP7_75t_SL g1779 ( 
.A(n_1599),
.Y(n_1779)
);

NAND2x1_ASAP7_75t_L g1780 ( 
.A(n_1557),
.B(n_1336),
.Y(n_1780)
);

NAND2x1p5_ASAP7_75t_L g1781 ( 
.A(n_1557),
.B(n_1216),
.Y(n_1781)
);

BUFx2_ASAP7_75t_L g1782 ( 
.A(n_1599),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1670),
.Y(n_1783)
);

OAI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1616),
.A2(n_1769),
.B(n_1678),
.Y(n_1784)
);

INVx2_ASAP7_75t_SL g1785 ( 
.A(n_1631),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1634),
.B(n_1630),
.Y(n_1786)
);

BUFx4f_ASAP7_75t_L g1787 ( 
.A(n_1631),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1681),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1735),
.A2(n_1653),
.B1(n_1634),
.B2(n_1770),
.Y(n_1789)
);

OR2x6_ASAP7_75t_L g1790 ( 
.A(n_1616),
.B(n_1769),
.Y(n_1790)
);

NAND2x1p5_ASAP7_75t_L g1791 ( 
.A(n_1689),
.B(n_1682),
.Y(n_1791)
);

BUFx6f_ASAP7_75t_SL g1792 ( 
.A(n_1766),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1635),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_SL g1794 ( 
.A1(n_1680),
.A2(n_1694),
.B1(n_1689),
.B2(n_1653),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1635),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1677),
.Y(n_1796)
);

INVx4_ASAP7_75t_L g1797 ( 
.A(n_1631),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1668),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1648),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1685),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1739),
.Y(n_1801)
);

AOI21x1_ASAP7_75t_L g1802 ( 
.A1(n_1780),
.A2(n_1765),
.B(n_1762),
.Y(n_1802)
);

BUFx2_ASAP7_75t_L g1803 ( 
.A(n_1726),
.Y(n_1803)
);

CKINVDCx11_ASAP7_75t_R g1804 ( 
.A(n_1628),
.Y(n_1804)
);

OR2x6_ASAP7_75t_L g1805 ( 
.A(n_1781),
.B(n_1650),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1735),
.A2(n_1634),
.B1(n_1771),
.B2(n_1770),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1664),
.Y(n_1807)
);

OAI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1736),
.A2(n_1633),
.B(n_1666),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1618),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1619),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1626),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1659),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_SL g1813 ( 
.A(n_1763),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1661),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1680),
.A2(n_1694),
.B1(n_1630),
.B2(n_1646),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1698),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1698),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1727),
.Y(n_1818)
);

AO21x1_ASAP7_75t_L g1819 ( 
.A1(n_1617),
.A2(n_1676),
.B(n_1671),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1649),
.Y(n_1820)
);

BUFx2_ASAP7_75t_L g1821 ( 
.A(n_1696),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1655),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1707),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1660),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1663),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1681),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1690),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1700),
.Y(n_1828)
);

INVx4_ASAP7_75t_L g1829 ( 
.A(n_1628),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1774),
.A2(n_1749),
.B(n_1733),
.Y(n_1830)
);

OR2x6_ASAP7_75t_SL g1831 ( 
.A(n_1656),
.B(n_1776),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1630),
.B(n_1623),
.Y(n_1832)
);

AOI21xp33_ASAP7_75t_L g1833 ( 
.A1(n_1747),
.A2(n_1637),
.B(n_1749),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1640),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1642),
.Y(n_1835)
);

BUFx3_ASAP7_75t_L g1836 ( 
.A(n_1763),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1686),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1709),
.B(n_1645),
.Y(n_1838)
);

CKINVDCx11_ASAP7_75t_R g1839 ( 
.A(n_1644),
.Y(n_1839)
);

INVx2_ASAP7_75t_SL g1840 ( 
.A(n_1740),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1647),
.Y(n_1841)
);

OAI21x1_ASAP7_75t_SL g1842 ( 
.A1(n_1744),
.A2(n_1759),
.B(n_1725),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1772),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1665),
.A2(n_1621),
.B1(n_1768),
.B2(n_1622),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1775),
.B(n_1704),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1729),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1686),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1716),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1729),
.Y(n_1849)
);

INVx3_ASAP7_75t_L g1850 ( 
.A(n_1632),
.Y(n_1850)
);

CKINVDCx11_ASAP7_75t_R g1851 ( 
.A(n_1644),
.Y(n_1851)
);

INVx3_ASAP7_75t_L g1852 ( 
.A(n_1763),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1658),
.Y(n_1853)
);

AO21x1_ASAP7_75t_L g1854 ( 
.A1(n_1671),
.A2(n_1676),
.B(n_1733),
.Y(n_1854)
);

AND2x4_ASAP7_75t_L g1855 ( 
.A(n_1671),
.B(n_1676),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1781),
.Y(n_1856)
);

BUFx4f_ASAP7_75t_SL g1857 ( 
.A(n_1766),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1771),
.A2(n_1773),
.B1(n_1679),
.B2(n_1695),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1738),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1773),
.A2(n_1679),
.B1(n_1695),
.B2(n_1629),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1731),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1757),
.Y(n_1862)
);

CKINVDCx11_ASAP7_75t_R g1863 ( 
.A(n_1624),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1622),
.Y(n_1864)
);

BUFx2_ASAP7_75t_L g1865 ( 
.A(n_1696),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1768),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1768),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1720),
.B(n_1691),
.Y(n_1868)
);

AOI21x1_ASAP7_75t_L g1869 ( 
.A1(n_1761),
.A2(n_1734),
.B(n_1673),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1719),
.A2(n_1683),
.B(n_1745),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1702),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1665),
.B(n_1767),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1697),
.A2(n_1720),
.B1(n_1629),
.B2(n_1701),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1708),
.Y(n_1874)
);

CKINVDCx11_ASAP7_75t_R g1875 ( 
.A(n_1624),
.Y(n_1875)
);

BUFx12f_ASAP7_75t_L g1876 ( 
.A(n_1776),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1712),
.Y(n_1877)
);

BUFx3_ASAP7_75t_L g1878 ( 
.A(n_1722),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1724),
.Y(n_1879)
);

OAI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1697),
.A2(n_1717),
.B1(n_1718),
.B2(n_1730),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1652),
.Y(n_1881)
);

BUFx3_ASAP7_75t_L g1882 ( 
.A(n_1722),
.Y(n_1882)
);

BUFx3_ASAP7_75t_L g1883 ( 
.A(n_1722),
.Y(n_1883)
);

BUFx3_ASAP7_75t_L g1884 ( 
.A(n_1740),
.Y(n_1884)
);

INVx8_ASAP7_75t_L g1885 ( 
.A(n_1682),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1652),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1705),
.Y(n_1887)
);

BUFx3_ASAP7_75t_L g1888 ( 
.A(n_1740),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1806),
.B(n_1756),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1805),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1812),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1845),
.B(n_1674),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1809),
.B(n_1674),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1810),
.B(n_1737),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1806),
.B(n_1789),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1837),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1789),
.B(n_1756),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1811),
.B(n_1838),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_1804),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1807),
.B(n_1737),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1822),
.B(n_1627),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1861),
.B(n_1639),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1783),
.Y(n_1903)
);

AND2x4_ASAP7_75t_SL g1904 ( 
.A(n_1797),
.B(n_1641),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1796),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1798),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1800),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1820),
.B(n_1641),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1801),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1828),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1790),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1834),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1835),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1841),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1868),
.A2(n_1778),
.B1(n_1754),
.B2(n_1741),
.Y(n_1915)
);

INVx2_ASAP7_75t_SL g1916 ( 
.A(n_1787),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1868),
.B(n_1705),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1786),
.B(n_1742),
.Y(n_1918)
);

INVx1_ASAP7_75t_SL g1919 ( 
.A(n_1813),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1843),
.Y(n_1920)
);

AND2x4_ASAP7_75t_SL g1921 ( 
.A(n_1797),
.B(n_1742),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1871),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1824),
.B(n_1779),
.Y(n_1923)
);

OAI21xp5_ASAP7_75t_SL g1924 ( 
.A1(n_1791),
.A2(n_1753),
.B(n_1760),
.Y(n_1924)
);

AND2x4_ASAP7_75t_L g1925 ( 
.A(n_1855),
.B(n_1682),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1874),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1793),
.B(n_1675),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1860),
.A2(n_1873),
.B1(n_1858),
.B2(n_1872),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1795),
.B(n_1675),
.Y(n_1929)
);

AO31x2_ASAP7_75t_L g1930 ( 
.A1(n_1853),
.A2(n_1732),
.A3(n_1758),
.B(n_1752),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1877),
.Y(n_1931)
);

INVx4_ASAP7_75t_L g1932 ( 
.A(n_1885),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1825),
.B(n_1625),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1799),
.B(n_1782),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1879),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1790),
.Y(n_1936)
);

AND2x4_ASAP7_75t_L g1937 ( 
.A(n_1855),
.B(n_1682),
.Y(n_1937)
);

AOI22xp5_ASAP7_75t_L g1938 ( 
.A1(n_1860),
.A2(n_1703),
.B1(n_1764),
.B2(n_1755),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1799),
.B(n_1743),
.Y(n_1939)
);

INVx4_ASAP7_75t_L g1940 ( 
.A(n_1885),
.Y(n_1940)
);

INVx2_ASAP7_75t_SL g1941 ( 
.A(n_1787),
.Y(n_1941)
);

BUFx2_ASAP7_75t_L g1942 ( 
.A(n_1884),
.Y(n_1942)
);

OAI21xp5_ASAP7_75t_SL g1943 ( 
.A1(n_1791),
.A2(n_1753),
.B(n_1715),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1858),
.A2(n_1741),
.B1(n_1687),
.B2(n_1693),
.Y(n_1944)
);

BUFx2_ASAP7_75t_L g1945 ( 
.A(n_1884),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1847),
.Y(n_1946)
);

INVx2_ASAP7_75t_SL g1947 ( 
.A(n_1888),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_SL g1948 ( 
.A1(n_1815),
.A2(n_1687),
.B1(n_1693),
.B2(n_1714),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_SL g1949 ( 
.A(n_1829),
.B(n_1636),
.Y(n_1949)
);

BUFx2_ASAP7_75t_L g1950 ( 
.A(n_1836),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1880),
.B(n_1715),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1830),
.B(n_1743),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1790),
.Y(n_1953)
);

AND2x4_ASAP7_75t_L g1954 ( 
.A(n_1832),
.B(n_1750),
.Y(n_1954)
);

INVx2_ASAP7_75t_SL g1955 ( 
.A(n_1857),
.Y(n_1955)
);

BUFx2_ASAP7_75t_L g1956 ( 
.A(n_1836),
.Y(n_1956)
);

INVx3_ASAP7_75t_SL g1957 ( 
.A(n_1813),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1803),
.B(n_1657),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1821),
.B(n_1777),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1816),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1817),
.Y(n_1961)
);

OAI22xp5_ASAP7_75t_L g1962 ( 
.A1(n_1794),
.A2(n_1687),
.B1(n_1693),
.B2(n_1714),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1833),
.B(n_1743),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1852),
.B(n_1643),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1794),
.A2(n_1723),
.B1(n_1714),
.B2(n_1711),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1788),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1852),
.B(n_1654),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1856),
.B(n_1859),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1827),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1865),
.B(n_1656),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1898),
.B(n_1862),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1891),
.Y(n_1972)
);

BUFx3_ASAP7_75t_L g1973 ( 
.A(n_1957),
.Y(n_1973)
);

BUFx3_ASAP7_75t_L g1974 ( 
.A(n_1957),
.Y(n_1974)
);

AOI222xp33_ASAP7_75t_L g1975 ( 
.A1(n_1895),
.A2(n_1928),
.B1(n_1951),
.B2(n_1917),
.C1(n_1949),
.C2(n_1943),
.Y(n_1975)
);

NAND2x1_ASAP7_75t_L g1976 ( 
.A(n_1932),
.B(n_1842),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1934),
.B(n_1788),
.Y(n_1977)
);

INVxp67_ASAP7_75t_L g1978 ( 
.A(n_1950),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1968),
.B(n_1826),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1911),
.B(n_1802),
.Y(n_1980)
);

NOR2xp67_ASAP7_75t_L g1981 ( 
.A(n_1932),
.B(n_1840),
.Y(n_1981)
);

AOI22xp33_ASAP7_75t_L g1982 ( 
.A1(n_1928),
.A2(n_1819),
.B1(n_1713),
.B2(n_1864),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1896),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1903),
.Y(n_1984)
);

AOI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1917),
.A2(n_1844),
.B1(n_1887),
.B2(n_1867),
.Y(n_1985)
);

BUFx2_ASAP7_75t_L g1986 ( 
.A(n_1956),
.Y(n_1986)
);

AND2x4_ASAP7_75t_L g1987 ( 
.A(n_1911),
.B(n_1784),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1936),
.B(n_1953),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1936),
.B(n_1620),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1905),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1953),
.B(n_1869),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1906),
.Y(n_1992)
);

NOR3xp33_ASAP7_75t_L g1993 ( 
.A(n_1924),
.B(n_1829),
.C(n_1808),
.Y(n_1993)
);

AOI22xp33_ASAP7_75t_L g1994 ( 
.A1(n_1895),
.A2(n_1866),
.B1(n_1870),
.B2(n_1849),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1907),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_L g1996 ( 
.A(n_1951),
.B(n_1846),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1952),
.B(n_1963),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1909),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1930),
.B(n_1848),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1910),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1912),
.Y(n_2001)
);

AND2x4_ASAP7_75t_L g2002 ( 
.A(n_1930),
.B(n_1814),
.Y(n_2002)
);

AOI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1900),
.A2(n_1894),
.B1(n_1938),
.B2(n_1944),
.Y(n_2003)
);

INVx2_ASAP7_75t_SL g2004 ( 
.A(n_1966),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1913),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1914),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_L g2007 ( 
.A(n_1923),
.B(n_1881),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1920),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1922),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1902),
.B(n_1818),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_L g2011 ( 
.A(n_1933),
.B(n_1886),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1926),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1931),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1935),
.Y(n_2014)
);

AND2x4_ASAP7_75t_SL g2015 ( 
.A(n_1940),
.B(n_1850),
.Y(n_2015)
);

BUFx3_ASAP7_75t_L g2016 ( 
.A(n_1904),
.Y(n_2016)
);

AOI22xp33_ASAP7_75t_L g2017 ( 
.A1(n_1944),
.A2(n_1688),
.B1(n_1721),
.B2(n_1692),
.Y(n_2017)
);

AND2x4_ASAP7_75t_L g2018 ( 
.A(n_1930),
.B(n_1853),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1901),
.B(n_1823),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1997),
.B(n_1948),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_2002),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1983),
.Y(n_2022)
);

OR2x2_ASAP7_75t_L g2023 ( 
.A(n_1997),
.B(n_1952),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_2002),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_2004),
.B(n_1889),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1971),
.B(n_1960),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1989),
.B(n_1948),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1989),
.B(n_1897),
.Y(n_2028)
);

OR2x2_ASAP7_75t_L g2029 ( 
.A(n_2004),
.B(n_1889),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1972),
.Y(n_2030)
);

OR2x6_ASAP7_75t_L g2031 ( 
.A(n_1976),
.B(n_1854),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1987),
.B(n_1897),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1984),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1987),
.B(n_1963),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1979),
.B(n_1961),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1986),
.B(n_2019),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1987),
.B(n_1939),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_2010),
.B(n_1969),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1983),
.Y(n_2039)
);

NOR2x1_ASAP7_75t_L g2040 ( 
.A(n_1973),
.B(n_1940),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1990),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1992),
.B(n_1908),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1988),
.B(n_1927),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1991),
.B(n_1946),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1995),
.B(n_1942),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1998),
.Y(n_2046)
);

NOR2xp33_ASAP7_75t_L g2047 ( 
.A(n_1978),
.B(n_1947),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2000),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_2001),
.B(n_1945),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1988),
.B(n_1929),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2005),
.Y(n_2051)
);

HB1xp67_ASAP7_75t_L g2052 ( 
.A(n_2036),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_2034),
.B(n_1999),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2030),
.Y(n_2054)
);

OAI211xp5_ASAP7_75t_L g2055 ( 
.A1(n_2040),
.A2(n_1975),
.B(n_2003),
.C(n_1993),
.Y(n_2055)
);

NAND4xp75_ASAP7_75t_L g2056 ( 
.A(n_2040),
.B(n_1981),
.C(n_1955),
.D(n_1941),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2051),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_L g2058 ( 
.A(n_2047),
.B(n_1973),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2030),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2051),
.Y(n_2060)
);

NOR2xp67_ASAP7_75t_L g2061 ( 
.A(n_2021),
.B(n_1974),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2034),
.B(n_1999),
.Y(n_2062)
);

INVx2_ASAP7_75t_SL g2063 ( 
.A(n_2044),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_2020),
.B(n_2006),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2033),
.Y(n_2065)
);

INVxp67_ASAP7_75t_SL g2066 ( 
.A(n_2044),
.Y(n_2066)
);

AND2x4_ASAP7_75t_L g2067 ( 
.A(n_2021),
.B(n_1991),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2022),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_2021),
.B(n_2024),
.Y(n_2069)
);

INVx2_ASAP7_75t_SL g2070 ( 
.A(n_2044),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2020),
.B(n_1999),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_2022),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2032),
.B(n_2018),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2032),
.B(n_2018),
.Y(n_2074)
);

AND2x4_ASAP7_75t_L g2075 ( 
.A(n_2024),
.B(n_1980),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2033),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2041),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2041),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2046),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2023),
.B(n_2008),
.Y(n_2080)
);

AND2x4_ASAP7_75t_SL g2081 ( 
.A(n_2031),
.B(n_1925),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_2039),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_2023),
.B(n_1977),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_2037),
.B(n_2018),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2043),
.B(n_2009),
.Y(n_2085)
);

OAI33xp33_ASAP7_75t_L g2086 ( 
.A1(n_2080),
.A2(n_2049),
.A3(n_2045),
.B1(n_1959),
.B2(n_1970),
.B3(n_2035),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2071),
.B(n_2073),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2071),
.B(n_2028),
.Y(n_2088)
);

AOI22xp33_ASAP7_75t_SL g2089 ( 
.A1(n_2055),
.A2(n_2016),
.B1(n_1974),
.B2(n_1890),
.Y(n_2089)
);

AOI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_2052),
.A2(n_1993),
.B1(n_2003),
.B2(n_2027),
.Y(n_2090)
);

OAI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_2061),
.A2(n_2031),
.B1(n_2016),
.B2(n_1919),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2064),
.B(n_2027),
.Y(n_2092)
);

INVx1_ASAP7_75t_SL g2093 ( 
.A(n_2058),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2054),
.Y(n_2094)
);

INVx3_ASAP7_75t_SL g2095 ( 
.A(n_2081),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_2068),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2068),
.Y(n_2097)
);

INVx2_ASAP7_75t_SL g2098 ( 
.A(n_2081),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_2083),
.B(n_2025),
.Y(n_2099)
);

INVx1_ASAP7_75t_SL g2100 ( 
.A(n_2083),
.Y(n_2100)
);

INVx2_ASAP7_75t_SL g2101 ( 
.A(n_2063),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_2072),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2085),
.B(n_2028),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2073),
.B(n_2037),
.Y(n_2104)
);

AOI32xp33_ASAP7_75t_L g2105 ( 
.A1(n_2053),
.A2(n_2015),
.A3(n_1982),
.B1(n_2007),
.B2(n_1996),
.Y(n_2105)
);

OAI21xp33_ASAP7_75t_L g2106 ( 
.A1(n_2053),
.A2(n_2062),
.B(n_2074),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_2075),
.B(n_2031),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_2074),
.B(n_2025),
.Y(n_2108)
);

OAI211xp5_ASAP7_75t_L g2109 ( 
.A1(n_2066),
.A2(n_1851),
.B(n_1839),
.C(n_1982),
.Y(n_2109)
);

INVx1_ASAP7_75t_SL g2110 ( 
.A(n_2056),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2054),
.Y(n_2111)
);

OAI32xp33_ASAP7_75t_L g2112 ( 
.A1(n_2063),
.A2(n_1831),
.A3(n_1662),
.B1(n_2038),
.B2(n_2026),
.Y(n_2112)
);

INVx1_ASAP7_75t_SL g2113 ( 
.A(n_2056),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2057),
.Y(n_2114)
);

HB1xp67_ASAP7_75t_L g2115 ( 
.A(n_2084),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2057),
.B(n_2043),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2062),
.B(n_2050),
.Y(n_2117)
);

AOI21xp5_ASAP7_75t_L g2118 ( 
.A1(n_2086),
.A2(n_2031),
.B(n_2070),
.Y(n_2118)
);

AOI22xp5_ASAP7_75t_L g2119 ( 
.A1(n_2090),
.A2(n_2075),
.B1(n_2070),
.B2(n_2067),
.Y(n_2119)
);

AOI221xp5_ASAP7_75t_L g2120 ( 
.A1(n_2112),
.A2(n_2084),
.B1(n_2048),
.B2(n_2046),
.C(n_2065),
.Y(n_2120)
);

AOI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_2089),
.A2(n_2075),
.B1(n_2067),
.B2(n_1996),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2099),
.Y(n_2122)
);

NAND3xp33_ASAP7_75t_L g2123 ( 
.A(n_2105),
.B(n_1915),
.C(n_2059),
.Y(n_2123)
);

OAI211xp5_ASAP7_75t_L g2124 ( 
.A1(n_2109),
.A2(n_1839),
.B(n_1851),
.C(n_1804),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2100),
.B(n_2059),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_L g2126 ( 
.A(n_2093),
.B(n_1899),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2099),
.Y(n_2127)
);

OR2x2_ASAP7_75t_L g2128 ( 
.A(n_2116),
.B(n_2029),
.Y(n_2128)
);

OA21x2_ASAP7_75t_L g2129 ( 
.A1(n_2110),
.A2(n_2082),
.B(n_2072),
.Y(n_2129)
);

NOR2x1_ASAP7_75t_SL g2130 ( 
.A(n_2098),
.B(n_2031),
.Y(n_2130)
);

OAI31xp33_ASAP7_75t_L g2131 ( 
.A1(n_2113),
.A2(n_2015),
.A3(n_2075),
.B(n_2067),
.Y(n_2131)
);

INVx1_ASAP7_75t_SL g2132 ( 
.A(n_2095),
.Y(n_2132)
);

OAI22xp33_ASAP7_75t_SL g2133 ( 
.A1(n_2095),
.A2(n_2048),
.B1(n_2065),
.B2(n_2060),
.Y(n_2133)
);

OAI22xp5_ASAP7_75t_L g2134 ( 
.A1(n_2098),
.A2(n_2067),
.B1(n_2007),
.B2(n_2011),
.Y(n_2134)
);

AOI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2107),
.A2(n_2050),
.B1(n_2069),
.B2(n_2060),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2094),
.Y(n_2136)
);

OR2x2_ASAP7_75t_L g2137 ( 
.A(n_2122),
.B(n_2103),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_SL g2138 ( 
.A(n_2133),
.B(n_2091),
.Y(n_2138)
);

AOI22xp5_ASAP7_75t_L g2139 ( 
.A1(n_2132),
.A2(n_2107),
.B1(n_2101),
.B2(n_2106),
.Y(n_2139)
);

AOI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_2121),
.A2(n_2107),
.B1(n_2101),
.B2(n_2092),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2127),
.Y(n_2141)
);

AO21x1_ASAP7_75t_L g2142 ( 
.A1(n_2118),
.A2(n_1904),
.B(n_1921),
.Y(n_2142)
);

AOI211xp5_ASAP7_75t_SL g2143 ( 
.A1(n_2124),
.A2(n_1857),
.B(n_1667),
.C(n_1925),
.Y(n_2143)
);

OAI32xp33_ASAP7_75t_L g2144 ( 
.A1(n_2134),
.A2(n_2115),
.A3(n_2108),
.B1(n_2087),
.B2(n_2112),
.Y(n_2144)
);

OAI211xp5_ASAP7_75t_L g2145 ( 
.A1(n_2131),
.A2(n_2120),
.B(n_2119),
.C(n_2126),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2123),
.B(n_2088),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2125),
.Y(n_2147)
);

AOI22xp5_ASAP7_75t_L g2148 ( 
.A1(n_2135),
.A2(n_2088),
.B1(n_2104),
.B2(n_2087),
.Y(n_2148)
);

OAI221xp5_ASAP7_75t_L g2149 ( 
.A1(n_2129),
.A2(n_2108),
.B1(n_1915),
.B2(n_2114),
.C(n_2111),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2136),
.B(n_2117),
.Y(n_2150)
);

AOI221xp5_ASAP7_75t_L g2151 ( 
.A1(n_2128),
.A2(n_2114),
.B1(n_2117),
.B2(n_2042),
.C(n_2076),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2130),
.B(n_2104),
.Y(n_2152)
);

AOI322xp5_ASAP7_75t_L g2153 ( 
.A1(n_2129),
.A2(n_2102),
.A3(n_2097),
.B1(n_2096),
.B2(n_2078),
.C1(n_2077),
.C2(n_2079),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2122),
.B(n_2076),
.Y(n_2154)
);

OAI321xp33_ASAP7_75t_L g2155 ( 
.A1(n_2121),
.A2(n_1994),
.A3(n_1892),
.B1(n_1916),
.B2(n_1893),
.C(n_1965),
.Y(n_2155)
);

CKINVDCx16_ASAP7_75t_R g2156 ( 
.A(n_2132),
.Y(n_2156)
);

OAI221xp5_ASAP7_75t_SL g2157 ( 
.A1(n_2132),
.A2(n_1994),
.B1(n_1985),
.B2(n_2029),
.C(n_1965),
.Y(n_2157)
);

INVx2_ASAP7_75t_SL g2158 ( 
.A(n_2156),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2137),
.Y(n_2159)
);

NOR2x1_ASAP7_75t_SL g2160 ( 
.A(n_2138),
.B(n_2145),
.Y(n_2160)
);

NAND3xp33_ASAP7_75t_SL g2161 ( 
.A(n_2142),
.B(n_2153),
.C(n_2139),
.Y(n_2161)
);

NOR2xp33_ASAP7_75t_SL g2162 ( 
.A(n_2144),
.B(n_1792),
.Y(n_2162)
);

NOR2x1_ASAP7_75t_L g2163 ( 
.A(n_2152),
.B(n_1651),
.Y(n_2163)
);

OAI211xp5_ASAP7_75t_L g2164 ( 
.A1(n_2143),
.A2(n_1875),
.B(n_1863),
.C(n_1885),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2146),
.B(n_2077),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2141),
.Y(n_2166)
);

XNOR2xp5_ASAP7_75t_L g2167 ( 
.A(n_2140),
.B(n_1785),
.Y(n_2167)
);

AOI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_2155),
.A2(n_1921),
.B(n_2096),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2154),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2147),
.Y(n_2170)
);

AOI22xp5_ASAP7_75t_L g2171 ( 
.A1(n_2148),
.A2(n_2069),
.B1(n_1792),
.B2(n_2011),
.Y(n_2171)
);

NAND3xp33_ASAP7_75t_L g2172 ( 
.A(n_2157),
.B(n_1875),
.C(n_1863),
.Y(n_2172)
);

NOR2x1_ASAP7_75t_L g2173 ( 
.A(n_2172),
.B(n_1638),
.Y(n_2173)
);

NOR4xp75_ASAP7_75t_L g2174 ( 
.A(n_2161),
.B(n_2149),
.C(n_2155),
.D(n_2150),
.Y(n_2174)
);

NAND4xp25_ASAP7_75t_L g2175 ( 
.A(n_2172),
.B(n_2151),
.C(n_1615),
.D(n_1937),
.Y(n_2175)
);

NAND5xp2_ASAP7_75t_L g2176 ( 
.A(n_2162),
.B(n_1710),
.C(n_2017),
.D(n_1958),
.E(n_1918),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2160),
.B(n_2078),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2158),
.Y(n_2178)
);

NAND3xp33_ASAP7_75t_L g2179 ( 
.A(n_2170),
.B(n_2168),
.C(n_2166),
.Y(n_2179)
);

NOR2x1_ASAP7_75t_L g2180 ( 
.A(n_2164),
.B(n_1878),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_2159),
.Y(n_2181)
);

AOI211xp5_ASAP7_75t_L g2182 ( 
.A1(n_2167),
.A2(n_1937),
.B(n_1967),
.C(n_1964),
.Y(n_2182)
);

NOR3xp33_ASAP7_75t_L g2183 ( 
.A(n_2163),
.B(n_1699),
.C(n_1706),
.Y(n_2183)
);

OA211x2_ASAP7_75t_L g2184 ( 
.A1(n_2165),
.A2(n_1876),
.B(n_1672),
.C(n_1684),
.Y(n_2184)
);

NOR3xp33_ASAP7_75t_L g2185 ( 
.A(n_2169),
.B(n_1706),
.C(n_1672),
.Y(n_2185)
);

BUFx6f_ASAP7_75t_L g2186 ( 
.A(n_2171),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2178),
.B(n_2097),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_2186),
.B(n_1684),
.Y(n_2188)
);

AO22x2_ASAP7_75t_L g2189 ( 
.A1(n_2181),
.A2(n_1751),
.B1(n_1669),
.B2(n_2012),
.Y(n_2189)
);

NOR3xp33_ASAP7_75t_SL g2190 ( 
.A(n_2179),
.B(n_1728),
.C(n_1962),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2177),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2185),
.B(n_2102),
.Y(n_2192)
);

NOR2x1_ASAP7_75t_L g2193 ( 
.A(n_2173),
.B(n_1878),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_2175),
.B(n_2079),
.Y(n_2194)
);

NOR2x1_ASAP7_75t_L g2195 ( 
.A(n_2180),
.B(n_1882),
.Y(n_2195)
);

NAND3xp33_ASAP7_75t_L g2196 ( 
.A(n_2186),
.B(n_1750),
.C(n_2013),
.Y(n_2196)
);

NOR3xp33_ASAP7_75t_L g2197 ( 
.A(n_2188),
.B(n_2176),
.C(n_2183),
.Y(n_2197)
);

AO22x2_ASAP7_75t_L g2198 ( 
.A1(n_2191),
.A2(n_2174),
.B1(n_2184),
.B2(n_2182),
.Y(n_2198)
);

NAND2x1p5_ASAP7_75t_L g2199 ( 
.A(n_2195),
.B(n_1882),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2187),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2192),
.Y(n_2201)
);

NOR3xp33_ASAP7_75t_L g2202 ( 
.A(n_2196),
.B(n_1728),
.C(n_1883),
.Y(n_2202)
);

NOR2xp33_ASAP7_75t_L g2203 ( 
.A(n_2194),
.B(n_2014),
.Y(n_2203)
);

BUFx3_ASAP7_75t_L g2204 ( 
.A(n_2189),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_2193),
.B(n_2069),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2200),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2204),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_2201),
.B(n_2190),
.Y(n_2208)
);

AND2x4_ASAP7_75t_L g2209 ( 
.A(n_2202),
.B(n_2197),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2198),
.B(n_2189),
.Y(n_2210)
);

INVxp33_ASAP7_75t_SL g2211 ( 
.A(n_2198),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2203),
.Y(n_2212)
);

AO21x2_ASAP7_75t_L g2213 ( 
.A1(n_2210),
.A2(n_2205),
.B(n_2199),
.Y(n_2213)
);

NOR3xp33_ASAP7_75t_L g2214 ( 
.A(n_2207),
.B(n_1883),
.C(n_1850),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2206),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2215),
.Y(n_2216)
);

OAI22xp5_ASAP7_75t_L g2217 ( 
.A1(n_2216),
.A2(n_2211),
.B1(n_2209),
.B2(n_2208),
.Y(n_2217)
);

AOI21xp5_ASAP7_75t_L g2218 ( 
.A1(n_2217),
.A2(n_2209),
.B(n_2213),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2218),
.B(n_2214),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2219),
.B(n_2212),
.Y(n_2220)
);

OR2x6_ASAP7_75t_L g2221 ( 
.A(n_2220),
.B(n_1954),
.Y(n_2221)
);

AOI21xp5_ASAP7_75t_L g2222 ( 
.A1(n_2221),
.A2(n_1748),
.B(n_1746),
.Y(n_2222)
);


endmodule