module fake_jpeg_3351_n_181 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_181);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_43),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_41),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_68),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_66),
.Y(n_72)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_74),
.B(n_77),
.Y(n_81)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

CKINVDCx9p33_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_76),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_67),
.Y(n_88)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_80),
.A2(n_50),
.B1(n_56),
.B2(n_66),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_94),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_62),
.B1(n_51),
.B2(n_68),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_87),
.B1(n_89),
.B2(n_51),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_90),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_67),
.B1(n_61),
.B2(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_61),
.B1(n_50),
.B2(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_58),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_62),
.B(n_58),
.C(n_59),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_71),
.B(n_54),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_95),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_52),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_53),
.C(n_48),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_57),
.C(n_46),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_110),
.B1(n_85),
.B2(n_4),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_105),
.C(n_2),
.Y(n_125)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_91),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_54),
.C(n_45),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_0),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_112),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_0),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_38),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_36),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_115),
.C(n_92),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_2),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_114),
.B(n_32),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_SL g115 ( 
.A(n_83),
.B(n_45),
.C(n_3),
.Y(n_115)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_83),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_118),
.Y(n_138)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_128),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_112),
.A2(n_113),
.B1(n_98),
.B2(n_109),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_144)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_123),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_91),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_132),
.C(n_5),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_3),
.B(n_5),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_10),
.B(n_11),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_129),
.B(n_6),
.Y(n_137)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_31),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_10),
.C(n_11),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_141),
.C(n_142),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_140),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_134),
.B(n_6),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_30),
.C(n_28),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_27),
.C(n_25),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_144),
.B(n_146),
.Y(n_154)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_122),
.B(n_9),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_12),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_130),
.B1(n_117),
.B2(n_123),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_116),
.A2(n_24),
.B(n_23),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_SL g157 ( 
.A1(n_149),
.A2(n_20),
.B(n_22),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_150),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_155),
.Y(n_166)
);

AOI221xp5_ASAP7_75t_L g153 ( 
.A1(n_151),
.A2(n_119),
.B1(n_117),
.B2(n_120),
.C(n_118),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g167 ( 
.A(n_153),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_158),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_139),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_159),
.B(n_161),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_12),
.C(n_13),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_141),
.C(n_142),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_156),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_164),
.B(n_168),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_154),
.A2(n_138),
.B1(n_143),
.B2(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_169),
.B(n_166),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_160),
.C(n_144),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_171),
.C(n_155),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_148),
.C(n_162),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_163),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_172),
.B(n_15),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_14),
.C(n_16),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_14),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_16),
.Y(n_181)
);


endmodule