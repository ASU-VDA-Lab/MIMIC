module real_jpeg_31430_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_0),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_0),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_0),
.Y(n_141)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_0),
.Y(n_280)
);

AND2x4_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_1),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_1),
.B(n_128),
.Y(n_127)
);

AND2x4_ASAP7_75t_L g175 ( 
.A(n_1),
.B(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_1),
.B(n_141),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_2),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_2),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_3),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_4),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_5),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_6),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_6),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_6),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_7),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_7),
.B(n_118),
.Y(n_117)
);

NAND2x1_ASAP7_75t_L g160 ( 
.A(n_7),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_7),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_7),
.B(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_7),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_8),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_8),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_8),
.B(n_126),
.Y(n_125)
);

NAND2x1_ASAP7_75t_SL g158 ( 
.A(n_8),
.B(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_9),
.Y(n_241)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_10),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_11),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_11),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_11),
.B(n_107),
.Y(n_106)
);

NAND2xp33_ASAP7_75t_SL g237 ( 
.A(n_11),
.B(n_238),
.Y(n_237)
);

NAND2x1_ASAP7_75t_L g252 ( 
.A(n_11),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_11),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_11),
.B(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_12),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_13),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_13),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_13),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_13),
.B(n_171),
.Y(n_170)
);

AND2x4_ASAP7_75t_SL g234 ( 
.A(n_13),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_13),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_13),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_13),
.B(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_14),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_14),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_14),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_15),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_15),
.B(n_77),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g184 ( 
.A(n_15),
.B(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_15),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_15),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_15),
.B(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_191),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_190),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_142),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_20),
.B(n_142),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_69),
.C(n_93),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_22),
.A2(n_69),
.B1(n_70),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_22),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_41),
.Y(n_22)
);

OAI21x1_ASAP7_75t_L g187 ( 
.A1(n_23),
.A2(n_188),
.B(n_189),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_26),
.B(n_31),
.C(n_36),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_29),
.Y(n_159)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_39),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_40),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_53),
.B2(n_54),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_42),
.B(n_53),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_42),
.B(n_53),
.Y(n_189)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_44),
.B(n_48),
.Y(n_92)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_52),
.Y(n_154)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_60),
.C(n_65),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_56),
.B1(n_65),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_58),
.Y(n_182)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_58),
.Y(n_235)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_58),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_59),
.Y(n_215)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_63),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_68),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_68),
.Y(n_255)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.C(n_92),
.Y(n_70)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_71),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.C(n_86),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_76),
.B(n_80),
.C(n_86),
.Y(n_199)
);

XNOR2x1_ASAP7_75t_L g297 ( 
.A(n_76),
.B(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2x1_ASAP7_75t_L g298 ( 
.A(n_80),
.B(n_86),
.Y(n_298)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_92),
.B(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_93),
.B(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_123),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_105),
.B1(n_121),
.B2(n_122),
.Y(n_94)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B(n_103),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_100),
.Y(n_104)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_99),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_102),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_103),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_121),
.C(n_123),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_112),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_113),
.C(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_130),
.C(n_137),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_124),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_169),
.B1(n_170),
.B2(n_173),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_125),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_125),
.A2(n_127),
.B1(n_173),
.B2(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_SL g233 ( 
.A(n_126),
.Y(n_233)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_127),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_129),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_130),
.A2(n_131),
.B1(n_137),
.B2(n_138),
.Y(n_202)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_164),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx4f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_160),
.B2(n_163),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_187),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_178),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_174),
.B2(n_175),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_SL g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_183),
.B1(n_184),
.B2(n_186),
.Y(n_179)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_221),
.B(n_308),
.Y(n_193)
);

NOR2xp67_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_218),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_195),
.B(n_218),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.C(n_203),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_196),
.B(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_203),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_210),
.C(n_216),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_204),
.B(n_210),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_206),
.B(n_207),
.Y(n_247)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_216),
.B(n_300),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_302),
.B(n_307),
.Y(n_221)
);

OAI21x1_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_290),
.B(n_301),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_258),
.B(n_289),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_242),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_225),
.B(n_242),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_234),
.C(n_236),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_226),
.A2(n_227),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_231),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_234),
.A2(n_236),
.B1(n_237),
.B2(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_234),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_248),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_244),
.B(n_247),
.C(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_248),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_249),
.B(n_252),
.C(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_256),
.Y(n_251)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_256),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_282),
.B(n_288),
.Y(n_258)
);

AOI21xp33_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_271),
.B(n_281),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_268),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_268),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_265),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_276),
.Y(n_271)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_284),
.Y(n_288)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_293),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_299),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_297),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_297),
.C(n_299),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_306),
.Y(n_307)
);


endmodule