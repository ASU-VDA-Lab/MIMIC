module fake_jpeg_16850_n_158 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_23),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_50),
.B1(n_52),
.B2(n_4),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_0),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_43),
.Y(n_82)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_64),
.B(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_6),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_87),
.B1(n_62),
.B2(n_6),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_1),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_78),
.B(n_3),
.Y(n_96)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_61),
.B1(n_59),
.B2(n_46),
.Y(n_87)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_61),
.B1(n_54),
.B2(n_60),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_98),
.B1(n_102),
.B2(n_106),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_57),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_95),
.B(n_96),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_99),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_55),
.B1(n_43),
.B2(n_53),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_88),
.A2(n_47),
.B1(n_44),
.B2(n_62),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

CKINVDCx10_ASAP7_75t_R g114 ( 
.A(n_103),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_107),
.B1(n_15),
.B2(n_16),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_83),
.B(n_5),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_108),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_7),
.B1(n_8),
.B2(n_14),
.Y(n_115)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_119),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_108),
.A3(n_98),
.B1(n_101),
.B2(n_20),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_104),
.Y(n_121)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_121),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_127),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_109),
.C(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_130),
.B(n_116),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_135),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_125),
.B1(n_111),
.B2(n_90),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_134),
.A2(n_114),
.B1(n_100),
.B2(n_19),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_111),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_91),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_139),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_143),
.B(n_17),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_137),
.C(n_140),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_145),
.C(n_143),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_146),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_141),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_18),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_149),
.B(n_22),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_24),
.C(n_26),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_28),
.C(n_29),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_31),
.Y(n_155)
);

NOR2xp67_ASAP7_75t_SL g156 ( 
.A(n_155),
.B(n_32),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_33),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_35),
.B(n_36),
.Y(n_158)
);


endmodule