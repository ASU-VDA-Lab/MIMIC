module fake_jpeg_4972_n_232 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_232);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_30),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_13),
.B(n_6),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_29),
.B(n_20),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_21),
.B1(n_15),
.B2(n_31),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_27),
.B1(n_18),
.B2(n_16),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_16),
.B1(n_18),
.B2(n_27),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_17),
.B1(n_23),
.B2(n_24),
.Y(n_69)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_54),
.Y(n_95)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AOI32xp33_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_17),
.A3(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_58),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_21),
.B1(n_33),
.B2(n_19),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_64),
.B1(n_68),
.B2(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_22),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_70),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_15),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_SL g89 ( 
.A1(n_61),
.A2(n_73),
.B(n_22),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_33),
.B(n_36),
.C(n_37),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_21),
.B1(n_13),
.B2(n_43),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_25),
.B1(n_51),
.B2(n_35),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_33),
.B1(n_35),
.B2(n_30),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_67),
.A2(n_17),
.B1(n_23),
.B2(n_22),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_49),
.B1(n_44),
.B2(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_22),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_50),
.C(n_41),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_73),
.Y(n_100)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_83),
.Y(n_108)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_85),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_62),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_55),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_92),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_48),
.B1(n_41),
.B2(n_30),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_90),
.B1(n_91),
.B2(n_72),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_72),
.B1(n_25),
.B2(n_37),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_67),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_59),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_96),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_106),
.B(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_99),
.B(n_1),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_109),
.B1(n_77),
.B2(n_80),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_73),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_88),
.Y(n_122)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_61),
.A3(n_66),
.B1(n_67),
.B2(n_54),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_53),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_67),
.B(n_71),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_111),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_115),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_113),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_79),
.A2(n_75),
.B(n_94),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_87),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_28),
.B1(n_51),
.B2(n_63),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_80),
.B1(n_63),
.B2(n_2),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_103),
.A2(n_91),
.B1(n_92),
.B2(n_82),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_82),
.B1(n_76),
.B2(n_78),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_131),
.B1(n_139),
.B2(n_100),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_122),
.B(n_125),
.Y(n_156)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_128),
.C(n_110),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_77),
.C(n_84),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_130),
.Y(n_142)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_0),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_134),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_6),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_135),
.Y(n_145)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_136),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_115),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_99),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_97),
.B(n_1),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_140),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_108),
.B1(n_97),
.B2(n_102),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_148),
.B1(n_159),
.B2(n_122),
.Y(n_169)
);

OAI32xp33_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_102),
.A3(n_106),
.B1(n_100),
.B2(n_101),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_157),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_149),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_117),
.B1(n_109),
.B2(n_105),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_121),
.C(n_129),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_160),
.C(n_134),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_123),
.Y(n_175)
);

NOR2x1_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_120),
.A2(n_111),
.B1(n_105),
.B2(n_113),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_116),
.C(n_3),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_173),
.C(n_149),
.Y(n_179)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_136),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_167),
.Y(n_181)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_133),
.B1(n_143),
.B2(n_153),
.Y(n_186)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_154),
.B(n_127),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_119),
.C(n_128),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_148),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

NAND2x1p5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_185),
.C(n_189),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_170),
.B1(n_168),
.B2(n_165),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_182),
.A2(n_184),
.B1(n_188),
.B2(n_167),
.Y(n_190)
);

XNOR2x1_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_150),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_186),
.B1(n_177),
.B2(n_189),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_150),
.B1(n_152),
.B2(n_144),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_164),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_143),
.B1(n_142),
.B2(n_139),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_137),
.C(n_153),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_178),
.B(n_127),
.Y(n_191)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_125),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_199),
.Y(n_204)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_195),
.A2(n_125),
.B(n_130),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_197),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_180),
.B(n_145),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_154),
.C(n_116),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_162),
.B1(n_131),
.B2(n_135),
.Y(n_200)
);

OAI321xp33_ASAP7_75t_L g203 ( 
.A1(n_200),
.A2(n_188),
.A3(n_184),
.B1(n_140),
.B2(n_147),
.C(n_130),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_185),
.C(n_146),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_200),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_203),
.A2(n_205),
.B1(n_2),
.B2(n_3),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_198),
.C(n_194),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_210),
.A2(n_212),
.B(n_215),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_190),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_211),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_202),
.A2(n_206),
.B1(n_208),
.B2(n_198),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_5),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_2),
.C(n_3),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_9),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_222),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_218),
.A2(n_220),
.B(n_7),
.C(n_10),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_210),
.B1(n_215),
.B2(n_6),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_12),
.C(n_4),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_5),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_224),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_226),
.C(n_218),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_223),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_227),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_12),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_4),
.Y(n_232)
);


endmodule