module real_jpeg_26446_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_139;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_1),
.A2(n_27),
.B1(n_39),
.B2(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_1),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_1),
.A2(n_32),
.B1(n_65),
.B2(n_75),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_1),
.A2(n_57),
.B1(n_58),
.B2(n_65),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_1),
.A2(n_43),
.B1(n_47),
.B2(n_65),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_2),
.A2(n_27),
.B1(n_39),
.B2(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_2),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_2),
.A2(n_68),
.B1(n_75),
.B2(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_2),
.A2(n_57),
.B1(n_58),
.B2(n_68),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_2),
.A2(n_43),
.B1(n_47),
.B2(n_68),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_3),
.A2(n_43),
.B1(n_47),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_3),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_4),
.A2(n_43),
.B1(n_47),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_4),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_5),
.Y(n_97)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_7),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_7),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_7),
.A2(n_27),
.B1(n_39),
.B2(n_73),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_7),
.A2(n_57),
.B1(n_58),
.B2(n_73),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_7),
.A2(n_43),
.B1(n_47),
.B2(n_73),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_9),
.A2(n_57),
.B1(n_58),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_9),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_9),
.A2(n_27),
.B1(n_39),
.B2(n_101),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_9),
.A2(n_43),
.B1(n_47),
.B2(n_101),
.Y(n_158)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_10),
.B(n_77),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_10),
.B(n_58),
.C(n_60),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_10),
.A2(n_27),
.B1(n_31),
.B2(n_39),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_10),
.B(n_69),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_10),
.A2(n_31),
.B1(n_57),
.B2(n_58),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_10),
.B(n_43),
.C(n_96),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_10),
.A2(n_42),
.B(n_205),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_11),
.A2(n_43),
.B1(n_47),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_11),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_14),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_14),
.A2(n_48),
.B1(n_57),
.B2(n_58),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_16),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_16),
.A2(n_41),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_140),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_139),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_114),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_21),
.B(n_114),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_84),
.C(n_103),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_22),
.B(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_53),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_23),
.B(n_54),
.C(n_70),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_151),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_30),
.C(n_34),
.Y(n_25)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_26),
.A2(n_27),
.B1(n_35),
.B2(n_39),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_26),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_83)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_27),
.A2(n_39),
.B1(n_60),
.B2(n_61),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_27),
.B(n_168),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_30),
.A2(n_31),
.B(n_36),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_31),
.B(n_99),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_31),
.B(n_44),
.Y(n_230)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_36),
.C(n_39),
.Y(n_34)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_40),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_45),
.B1(n_49),
.B2(n_51),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_42),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_42),
.A2(n_87),
.B1(n_89),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_42),
.A2(n_46),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_42),
.B(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_42),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_43),
.A2(n_47),
.B1(n_96),
.B2(n_98),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_47),
.B(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_50),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_51),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_70),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_63),
.B(n_66),
.Y(n_54)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_55),
.A2(n_66),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_56),
.A2(n_136),
.B(n_137),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_56),
.A2(n_137),
.B(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_57),
.A2(n_58),
.B1(n_96),
.B2(n_98),
.Y(n_95)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_58),
.B(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_69),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_67),
.B(n_110),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_76),
.B(n_78),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_72),
.A2(n_77),
.B1(n_82),
.B2(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_80),
.Y(n_113)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_84),
.B(n_103),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_92),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_85),
.B(n_92),
.Y(n_138)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_91),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_93),
.A2(n_192),
.B(n_193),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_93),
.A2(n_193),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_94),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_94),
.A2(n_125),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_100),
.B(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_99),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_99),
.A2(n_106),
.B(n_178),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.C(n_111),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_107),
.B(n_125),
.Y(n_193)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_109),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_128),
.B2(n_129),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_122),
.B1(n_126),
.B2(n_127),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_119),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_138),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_249),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_162),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_160),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_144),
.B(n_160),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.C(n_152),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_145),
.A2(n_146),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_152),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.C(n_157),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_187),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_159),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_242),
.B(n_248),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_194),
.B(n_241),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_183),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_165),
.B(n_183),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_176),
.C(n_180),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_166),
.B(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_169),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B(n_174),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_176),
.A2(n_180),
.B1(n_181),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_176),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_188),
.B2(n_189),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_184),
.B(n_190),
.C(n_191),
.Y(n_247)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_235),
.B(n_240),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_214),
.B(n_234),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_208),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_208),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_202),
.C(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_204),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_212),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_222),
.B(n_233),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_220),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_218),
.A2(n_226),
.B(n_227),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_228),
.B(n_232),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_225),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_239),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_247),
.Y(n_248)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);


endmodule