module real_jpeg_6163_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_1),
.Y(n_123)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_1),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_2),
.B(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_2),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_2),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_2),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_2),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_2),
.B(n_215),
.Y(n_413)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_4),
.Y(n_127)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_4),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_4),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_5),
.B(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_5),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_5),
.B(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_5),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_5),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_6),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_6),
.B(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_6),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_6),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_6),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_6),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_6),
.B(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_6),
.B(n_394),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_7),
.Y(n_102)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_7),
.Y(n_145)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_9),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_9),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_9),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_9),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_9),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g235 ( 
.A(n_9),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_9),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_9),
.B(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_10),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_10),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_10),
.Y(n_254)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_10),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_10),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_11),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_11),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_11),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_11),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_11),
.B(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_11),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_11),
.B(n_36),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_11),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_12),
.B(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_12),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_12),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_12),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_12),
.B(n_122),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_12),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_12),
.B(n_182),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_12),
.B(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_13),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_13),
.Y(n_183)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_13),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_14),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_14),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_14),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_14),
.B(n_170),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_14),
.B(n_351),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_15),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_15),
.B(n_82),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_15),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_15),
.B(n_36),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_15),
.B(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_15),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_15),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_15),
.B(n_373),
.Y(n_425)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

A2O1A1O1Ixp25_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_110),
.B(n_350),
.C(n_509),
.D(n_511),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_71),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_20),
.B(n_71),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_56),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_44),
.C(n_48),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_22),
.A2(n_23),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_43),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_26),
.A2(n_27),
.B1(n_63),
.B2(n_67),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_26),
.A2(n_27),
.B1(n_230),
.B2(n_237),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_L g511 ( 
.A(n_26),
.B(n_60),
.C(n_63),
.Y(n_511)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_27),
.B(n_33),
.C(n_39),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_27),
.B(n_317),
.C(n_318),
.Y(n_316)
);

OR2x2_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_29),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_30),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_30),
.Y(n_221)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_31),
.Y(n_131)
);

OR2x2_ASAP7_75t_SL g34 ( 
.A(n_32),
.B(n_35),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_32),
.B(n_105),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_32),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_49),
.C(n_54),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_33),
.A2(n_34),
.B1(n_49),
.B2(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_33),
.A2(n_34),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_34),
.B(n_150),
.C(n_155),
.Y(n_251)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_38),
.Y(n_179)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_38),
.Y(n_200)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_39),
.A2(n_43),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_39),
.B(n_335),
.C(n_339),
.Y(n_484)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_47),
.B(n_61),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_98),
.C(n_103),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_49),
.A2(n_109),
.B1(n_177),
.B2(n_185),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_49),
.B(n_178),
.C(n_181),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_49),
.A2(n_103),
.B1(n_104),
.B2(n_109),
.Y(n_483)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_52),
.Y(n_370)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_52),
.Y(n_387)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_53),
.Y(n_135)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_53),
.Y(n_213)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_53),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g399 ( 
.A(n_53),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_69),
.B2(n_70),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_68),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_59),
.A2(n_60),
.B1(n_476),
.B2(n_477),
.Y(n_475)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_84),
.C(n_88),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_63),
.A2(n_67),
.B1(n_301),
.B2(n_303),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_63),
.B(n_242),
.C(n_276),
.Y(n_347)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_65),
.B(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_66),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_69),
.B(n_510),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.C(n_92),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_72),
.A2(n_73),
.B1(n_77),
.B2(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_77),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.C(n_90),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_79),
.B1(n_90),
.B2(n_96),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_83),
.B(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_84),
.A2(n_88),
.B1(n_245),
.B2(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_84),
.Y(n_478)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_88),
.A2(n_239),
.B1(n_240),
.B2(n_245),
.Y(n_238)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_88),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_88),
.B(n_136),
.C(n_242),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_90),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_90),
.A2(n_96),
.B1(n_311),
.B2(n_315),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_90),
.B(n_315),
.C(n_345),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_90),
.A2(n_96),
.B1(n_349),
.B2(n_350),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_92),
.B(n_505),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.C(n_107),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_93),
.A2(n_94),
.B1(n_487),
.B2(n_488),
.Y(n_486)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_96),
.B(n_347),
.C(n_350),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_97),
.B(n_107),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_98),
.B(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_103),
.A2(n_104),
.B1(n_136),
.B2(n_241),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_103),
.A2(n_104),
.B1(n_276),
.B2(n_302),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_133),
.C(n_136),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_104),
.B(n_276),
.C(n_327),
.Y(n_485)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_106),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_503),
.B(n_508),
.Y(n_110)
);

AOI21x1_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_469),
.B(n_500),
.Y(n_111)
);

AO21x1_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_321),
.B(n_353),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_284),
.B(n_320),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_260),
.B(n_283),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_115),
.B(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_223),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_116),
.B(n_223),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_175),
.C(n_205),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_117),
.B(n_282),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_146),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_118),
.B(n_147),
.C(n_158),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_132),
.C(n_137),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_119),
.B(n_279),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g513 ( 
.A(n_119),
.Y(n_513)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_124),
.CI(n_128),
.CON(n_119),
.SN(n_119)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_120),
.B(n_124),
.C(n_128),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx8_ASAP7_75t_L g365 ( 
.A(n_123),
.Y(n_365)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_127),
.Y(n_410)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_132),
.A2(n_137),
.B1(n_138),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_132),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_133),
.B(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_136),
.A2(n_241),
.B1(n_242),
.B2(n_244),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_136),
.Y(n_241)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_139),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_277)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_158),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_154),
.B1(n_155),
.B2(n_157),
.Y(n_149)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_150),
.A2(n_157),
.B1(n_191),
.B2(n_192),
.Y(n_388)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_165),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_160),
.B(n_161),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_159),
.B(n_166),
.C(n_173),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_164),
.B(n_406),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_173),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_170),
.Y(n_429)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_171),
.Y(n_406)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_171),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_174),
.B(n_372),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_174),
.B(n_384),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_174),
.B(n_420),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_175),
.B(n_205),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_186),
.C(n_188),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_176),
.A2(n_186),
.B1(n_187),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_176),
.Y(n_265)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_180),
.B1(n_181),
.B2(n_184),
.Y(n_177)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_178),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_180),
.A2(n_181),
.B1(n_292),
.B2(n_297),
.Y(n_291)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_181),
.B(n_293),
.C(n_294),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_188),
.B(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_195),
.C(n_201),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_189),
.A2(n_190),
.B1(n_456),
.B2(n_457),
.Y(n_455)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_195),
.A2(n_196),
.B1(n_201),
.B2(n_202),
.Y(n_457)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_200),
.Y(n_337)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx4_ASAP7_75t_SL g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_222),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_208),
.C(n_222),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_218),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_214),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_214),
.C(n_218),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_210),
.A2(n_335),
.B1(n_338),
.B2(n_339),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_210),
.Y(n_339)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_213),
.Y(n_296)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g328 ( 
.A(n_221),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_224),
.B(n_226),
.C(n_259),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_246),
.B1(n_258),
.B2(n_259),
.Y(n_225)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_238),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_228),
.B(n_229),
.C(n_238),
.Y(n_305)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_235),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_231),
.Y(n_317)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_235),
.Y(n_318)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_242),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_242),
.A2(n_244),
.B1(n_276),
.B2(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_242),
.A2(n_244),
.B1(n_379),
.B2(n_380),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_244),
.B(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_247),
.B(n_249),
.C(n_250),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_251),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_253),
.B(n_255),
.C(n_308),
.Y(n_307)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_281),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_261),
.B(n_281),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.C(n_278),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_262),
.A2(n_263),
.B1(n_462),
.B2(n_463),
.Y(n_461)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_266),
.B(n_278),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.C(n_277),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_267),
.B(n_449),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_269),
.B(n_277),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_274),
.C(n_276),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_270),
.A2(n_271),
.B1(n_274),
.B2(n_275),
.Y(n_376)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_273),
.Y(n_373)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_276),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_276),
.A2(n_302),
.B1(n_375),
.B2(n_376),
.Y(n_374)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_285),
.B(n_321),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_286),
.B(n_287),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_287),
.B(n_322),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_287),
.B(n_322),
.Y(n_468)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_304),
.CI(n_319),
.CON(n_287),
.SN(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_300),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_298),
.B2(n_299),
.Y(n_289)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_290),
.B(n_299),
.C(n_300),
.Y(n_342)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_291),
.Y(n_299)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_292),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

INVx4_ASAP7_75t_SL g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_307),
.C(n_309),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_316),
.Y(n_309)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_311),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_316),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_323),
.B(n_325),
.C(n_340),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_340),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_326),
.B(n_331),
.C(n_332),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_335),
.Y(n_338)
);

INVx6_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx8_ASAP7_75t_L g381 ( 
.A(n_337),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_343),
.B2(n_352),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_341),
.B(n_344),
.C(n_346),
.Y(n_496)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_343),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_346),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_350),
.Y(n_349)
);

OAI31xp33_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_465),
.A3(n_466),
.B(n_468),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_459),
.B(n_464),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_444),
.B(n_458),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_401),
.B(n_443),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_389),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_358),
.B(n_389),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_377),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_374),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_360),
.B(n_374),
.C(n_377),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_366),
.C(n_371),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_361),
.A2(n_362),
.B1(n_366),
.B2(n_367),
.Y(n_391)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx8_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_371),
.B(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_382),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_378),
.B(n_453),
.C(n_454),
.Y(n_452)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_388),
.Y(n_382)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_383),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_385),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_388),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_392),
.C(n_400),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_390),
.B(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_392),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_392),
.A2(n_400),
.B1(n_435),
.B2(n_441),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_397),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_393),
.Y(n_433)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_396),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_397),
.Y(n_434)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_400),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_437),
.B(n_442),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_422),
.B(n_436),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_411),
.B(n_421),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_407),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_419),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_412),
.B(n_419),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_414),
.B(n_418),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_413),
.B(n_414),
.Y(n_418)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_418),
.A2(n_424),
.B1(n_430),
.B2(n_431),
.Y(n_423)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_418),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_432),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_432),
.Y(n_436)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_424),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_425),
.A2(n_426),
.B(n_430),
.Y(n_438)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_433),
.A2(n_434),
.B(n_435),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_439),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_445),
.B(n_446),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_447),
.A2(n_448),
.B1(n_450),
.B2(n_451),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_452),
.C(n_455),
.Y(n_460)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_455),
.Y(n_451)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_461),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_460),
.B(n_461),
.Y(n_464)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_462),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_497),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_470),
.A2(n_501),
.B(n_502),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_489),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_471),
.B(n_489),
.Y(n_502)
);

BUFx24_ASAP7_75t_SL g512 ( 
.A(n_471),
.Y(n_512)
);

FAx1_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_480),
.CI(n_486),
.CON(n_471),
.SN(n_471)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_472),
.B(n_480),
.C(n_486),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_475),
.C(n_479),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_473),
.A2(n_474),
.B1(n_491),
.B2(n_492),
.Y(n_490)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_479),
.Y(n_491)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_484),
.C(n_485),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_481),
.A2(n_482),
.B1(n_494),
.B2(n_495),
.Y(n_493)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_485),
.Y(n_495)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_487),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_493),
.C(n_496),
.Y(n_489)
);

FAx1_ASAP7_75t_SL g499 ( 
.A(n_490),
.B(n_493),
.CI(n_496),
.CON(n_499),
.SN(n_499)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_491),
.Y(n_492)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_499),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_498),
.B(n_499),
.Y(n_501)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_499),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_507),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_504),
.B(n_507),
.Y(n_508)
);


endmodule