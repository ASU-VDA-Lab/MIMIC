module fake_netlist_6_993_n_817 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_817);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_817;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_179;
wire n_248;
wire n_222;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_787;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_45),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_88),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_126),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_6),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_81),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_6),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_51),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_161),
.Y(n_182)
);

NOR2xp67_ASAP7_75t_L g183 ( 
.A(n_18),
.B(n_63),
.Y(n_183)
);

NOR2xp67_ASAP7_75t_L g184 ( 
.A(n_13),
.B(n_21),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_64),
.B(n_17),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_120),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_83),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_170),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_99),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_47),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_14),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_103),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_30),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_46),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_62),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_33),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_95),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_40),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_29),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_102),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_35),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_91),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_70),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_138),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_68),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_109),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_4),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_139),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_100),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_84),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_80),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_141),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_135),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_66),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_151),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_14),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_133),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_76),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_113),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_112),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_89),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_31),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_86),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_124),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_90),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_52),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_104),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_147),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_8),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_166),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_156),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_116),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_71),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_106),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_2),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_41),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_125),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_4),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_38),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_0),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_177),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_192),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_208),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_207),
.B(n_0),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_1),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_1),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_219),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

AND2x6_ASAP7_75t_L g256 ( 
.A(n_191),
.B(n_19),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_225),
.B(n_183),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g258 ( 
.A1(n_209),
.A2(n_2),
.B(n_3),
.Y(n_258)
);

OA21x2_ASAP7_75t_L g259 ( 
.A1(n_229),
.A2(n_3),
.B(n_5),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_172),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_185),
.B(n_227),
.Y(n_261)
);

AND2x4_ASAP7_75t_L g262 ( 
.A(n_175),
.B(n_5),
.Y(n_262)
);

AND2x2_ASAP7_75t_SL g263 ( 
.A(n_229),
.B(n_7),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_175),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_213),
.B(n_226),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_221),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_213),
.Y(n_267)
);

BUFx8_ASAP7_75t_SL g268 ( 
.A(n_210),
.Y(n_268)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_221),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_221),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_179),
.B(n_7),
.Y(n_271)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_221),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_226),
.B(n_8),
.Y(n_273)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_173),
.Y(n_274)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_176),
.Y(n_275)
);

OAI22x1_ASAP7_75t_R g276 ( 
.A1(n_210),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_174),
.B(n_9),
.Y(n_277)
);

AND2x6_ASAP7_75t_L g278 ( 
.A(n_181),
.B(n_20),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_188),
.Y(n_279)
);

AND2x4_ASAP7_75t_L g280 ( 
.A(n_198),
.B(n_10),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_201),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_202),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_203),
.Y(n_283)
);

AND2x6_ASAP7_75t_L g284 ( 
.A(n_214),
.B(n_22),
.Y(n_284)
);

AND2x6_ASAP7_75t_L g285 ( 
.A(n_215),
.B(n_218),
.Y(n_285)
);

OA21x2_ASAP7_75t_L g286 ( 
.A1(n_230),
.A2(n_11),
.B(n_12),
.Y(n_286)
);

BUFx8_ASAP7_75t_SL g287 ( 
.A(n_182),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_238),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_236),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_237),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_178),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_180),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_249),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_267),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_257),
.B(n_184),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_264),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_249),
.Y(n_299)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_260),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_12),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_249),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_252),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_268),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_252),
.Y(n_307)
);

BUFx6f_ASAP7_75t_SL g308 ( 
.A(n_262),
.Y(n_308)
);

BUFx8_ASAP7_75t_SL g309 ( 
.A(n_268),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_248),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_252),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_254),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_287),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_261),
.B(n_242),
.Y(n_315)
);

NAND2xp33_ASAP7_75t_SL g316 ( 
.A(n_261),
.B(n_199),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_266),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_266),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_255),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_266),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_263),
.B(n_206),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_247),
.Y(n_323)
);

INVx5_ASAP7_75t_L g324 ( 
.A(n_256),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_270),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_263),
.B(n_262),
.Y(n_326)
);

NAND3xp33_ASAP7_75t_L g327 ( 
.A(n_265),
.B(n_212),
.C(n_187),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_247),
.Y(n_328)
);

NOR2x1p5_ASAP7_75t_L g329 ( 
.A(n_250),
.B(n_251),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_289),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_270),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_289),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_289),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_270),
.Y(n_334)
);

NOR2x1p5_ASAP7_75t_L g335 ( 
.A(n_250),
.B(n_186),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_290),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_290),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_290),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_246),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_245),
.Y(n_340)
);

AOI21x1_ASAP7_75t_L g341 ( 
.A1(n_251),
.A2(n_239),
.B(n_224),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_265),
.B(n_13),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_335),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_292),
.B(n_243),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_323),
.B(n_273),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_298),
.Y(n_346)
);

NOR3xp33_ASAP7_75t_L g347 ( 
.A(n_316),
.B(n_277),
.C(n_253),
.Y(n_347)
);

NAND2xp33_ASAP7_75t_L g348 ( 
.A(n_315),
.B(n_284),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_315),
.B(n_275),
.Y(n_349)
);

NOR3xp33_ASAP7_75t_L g350 ( 
.A(n_316),
.B(n_322),
.C(n_296),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_274),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_298),
.B(n_275),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_295),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_294),
.B(n_274),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_294),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_296),
.B(n_274),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_310),
.Y(n_357)
);

NOR3xp33_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_277),
.C(n_253),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_299),
.B(n_274),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_313),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_295),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_319),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_299),
.B(n_285),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_300),
.B(n_244),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_297),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_305),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_306),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_300),
.B(n_280),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_312),
.B(n_280),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_302),
.Y(n_371)
);

NOR2x1p5_ASAP7_75t_L g372 ( 
.A(n_301),
.B(n_312),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_302),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_303),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_303),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_307),
.B(n_311),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_327),
.B(n_244),
.Y(n_377)
);

INVx8_ASAP7_75t_L g378 ( 
.A(n_308),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_307),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_311),
.B(n_285),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_317),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_317),
.B(n_285),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_318),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_326),
.B(n_287),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_318),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_300),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_320),
.B(n_285),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_320),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_325),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_325),
.B(n_246),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_337),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_331),
.Y(n_392)
);

AOI221xp5_ASAP7_75t_L g393 ( 
.A1(n_326),
.A2(n_271),
.B1(n_228),
.B2(n_240),
.C(n_189),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_308),
.B(n_190),
.Y(n_394)
);

NAND3xp33_ASAP7_75t_L g395 ( 
.A(n_342),
.B(n_258),
.C(n_259),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_331),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_308),
.B(n_193),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_334),
.B(n_246),
.Y(n_398)
);

OR2x6_ASAP7_75t_L g399 ( 
.A(n_340),
.B(n_276),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_321),
.B(n_246),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_334),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_330),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_321),
.B(n_194),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_321),
.B(n_195),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_293),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_332),
.B(n_284),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_333),
.B(n_336),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_338),
.B(n_269),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_304),
.B(n_256),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_358),
.B(n_284),
.Y(n_410)
);

A2O1A1Ixp33_ASAP7_75t_L g411 ( 
.A1(n_377),
.A2(n_234),
.B(n_197),
.C(n_200),
.Y(n_411)
);

O2A1O1Ixp33_ASAP7_75t_L g412 ( 
.A1(n_344),
.A2(n_259),
.B(n_258),
.C(n_286),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_348),
.A2(n_339),
.B(n_324),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

AOI21x1_ASAP7_75t_L g415 ( 
.A1(n_363),
.A2(n_341),
.B(n_286),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_343),
.B(n_364),
.Y(n_416)
);

OAI321xp33_ASAP7_75t_L g417 ( 
.A1(n_395),
.A2(n_284),
.A3(n_278),
.B1(n_17),
.B2(n_18),
.C(n_15),
.Y(n_417)
);

INVx5_ASAP7_75t_L g418 ( 
.A(n_406),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_347),
.B(n_278),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_349),
.B(n_314),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_395),
.A2(n_231),
.B1(n_204),
.B2(n_205),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_370),
.B(n_278),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_357),
.B(n_278),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_374),
.A2(n_339),
.B(n_324),
.Y(n_424)
);

BUFx12f_ASAP7_75t_L g425 ( 
.A(n_386),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_406),
.A2(n_278),
.B(n_324),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_360),
.B(n_324),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_393),
.B(n_304),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_380),
.A2(n_339),
.B(n_324),
.Y(n_429)
);

AO21x1_ASAP7_75t_L g430 ( 
.A1(n_350),
.A2(n_256),
.B(n_15),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_362),
.B(n_256),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_365),
.B(n_366),
.Y(n_432)
);

AND2x2_ASAP7_75t_SL g433 ( 
.A(n_384),
.B(n_309),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_368),
.B(n_256),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_353),
.B(n_196),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_382),
.A2(n_269),
.B(n_272),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_369),
.B(n_211),
.Y(n_437)
);

NOR2x1_ASAP7_75t_L g438 ( 
.A(n_403),
.B(n_216),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_361),
.B(n_352),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_387),
.A2(n_222),
.B(n_235),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_355),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_353),
.B(n_217),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_376),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_353),
.B(n_405),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_354),
.A2(n_359),
.B(n_407),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_345),
.A2(n_351),
.B(n_398),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_390),
.A2(n_269),
.B(n_272),
.Y(n_447)
);

AOI21xp33_ASAP7_75t_L g448 ( 
.A1(n_356),
.A2(n_233),
.B(n_223),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_408),
.A2(n_269),
.B(n_272),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_367),
.B(n_220),
.Y(n_450)
);

O2A1O1Ixp33_ASAP7_75t_L g451 ( 
.A1(n_409),
.A2(n_404),
.B(n_402),
.C(n_401),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_394),
.B(n_309),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_372),
.A2(n_272),
.B1(n_23),
.B2(n_24),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_367),
.B(n_25),
.Y(n_454)
);

A2O1A1Ixp33_ASAP7_75t_L g455 ( 
.A1(n_397),
.A2(n_16),
.B(n_26),
.C(n_27),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_375),
.A2(n_105),
.B(n_28),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_391),
.A2(n_16),
.B1(n_32),
.B2(n_34),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_371),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_400),
.B(n_36),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_391),
.B(n_37),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_378),
.B(n_39),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_378),
.B(n_42),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_389),
.B(n_381),
.Y(n_463)
);

A2O1A1Ixp33_ASAP7_75t_L g464 ( 
.A1(n_373),
.A2(n_43),
.B(n_44),
.C(n_48),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_378),
.B(n_49),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_381),
.B(n_50),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_381),
.B(n_53),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_379),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_385),
.A2(n_396),
.B1(n_388),
.B2(n_392),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_383),
.A2(n_57),
.B(n_58),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_399),
.B(n_383),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_383),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_399),
.A2(n_65),
.B(n_67),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_392),
.A2(n_69),
.B(n_72),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_392),
.B(n_73),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_399),
.A2(n_74),
.B(n_75),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_364),
.B(n_77),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_343),
.B(n_78),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_343),
.A2(n_79),
.B1(n_82),
.B2(n_85),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_416),
.B(n_87),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_452),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_471),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_473),
.B(n_92),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_413),
.A2(n_429),
.B(n_445),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_444),
.B(n_93),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_441),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_420),
.B(n_428),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_412),
.A2(n_94),
.B(n_96),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g489 ( 
.A(n_414),
.Y(n_489)
);

NOR2x1_ASAP7_75t_SL g490 ( 
.A(n_418),
.B(n_98),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_439),
.B(n_101),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_410),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_444),
.B(n_111),
.Y(n_493)
);

OAI22xp33_ASAP7_75t_L g494 ( 
.A1(n_417),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_443),
.B(n_118),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_477),
.B(n_119),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_458),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_415),
.A2(n_121),
.B(n_122),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_423),
.A2(n_123),
.B(n_127),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_432),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_463),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_426),
.A2(n_446),
.B(n_434),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g503 ( 
.A(n_418),
.B(n_128),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_431),
.A2(n_171),
.B(n_130),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_478),
.B(n_129),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_437),
.B(n_131),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_425),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_427),
.A2(n_169),
.B(n_134),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_438),
.B(n_132),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_419),
.A2(n_136),
.B(n_137),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_422),
.A2(n_418),
.B(n_450),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_440),
.B(n_140),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_418),
.A2(n_142),
.B(n_143),
.Y(n_513)
);

BUFx4f_ASAP7_75t_L g514 ( 
.A(n_433),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_440),
.B(n_144),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_421),
.B(n_145),
.Y(n_516)
);

NAND2x1p5_ASAP7_75t_L g517 ( 
.A(n_461),
.B(n_465),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_469),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_424),
.A2(n_168),
.B(n_150),
.Y(n_519)
);

OAI21xp33_ASAP7_75t_L g520 ( 
.A1(n_473),
.A2(n_149),
.B(n_152),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_435),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_451),
.A2(n_153),
.B(n_154),
.Y(n_522)
);

AOI21x1_ASAP7_75t_L g523 ( 
.A1(n_436),
.A2(n_155),
.B(n_158),
.Y(n_523)
);

AO31x2_ASAP7_75t_L g524 ( 
.A1(n_430),
.A2(n_455),
.A3(n_411),
.B(n_464),
.Y(n_524)
);

NAND2x1p5_ASAP7_75t_L g525 ( 
.A(n_462),
.B(n_159),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_417),
.A2(n_163),
.B(n_164),
.Y(n_526)
);

AO31x2_ASAP7_75t_L g527 ( 
.A1(n_479),
.A2(n_165),
.A3(n_167),
.B(n_467),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_453),
.Y(n_528)
);

OAI21xp33_ASAP7_75t_L g529 ( 
.A1(n_457),
.A2(n_459),
.B(n_448),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_442),
.B(n_476),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_466),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_475),
.B(n_460),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_472),
.Y(n_533)
);

AO31x2_ASAP7_75t_L g534 ( 
.A1(n_454),
.A2(n_456),
.A3(n_470),
.B(n_474),
.Y(n_534)
);

AO31x2_ASAP7_75t_L g535 ( 
.A1(n_447),
.A2(n_430),
.A3(n_419),
.B(n_410),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_449),
.A2(n_445),
.B(n_423),
.Y(n_536)
);

AOI21xp33_ASAP7_75t_L g537 ( 
.A1(n_468),
.A2(n_416),
.B(n_393),
.Y(n_537)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_481),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_482),
.B(n_493),
.Y(n_539)
);

OR2x6_ASAP7_75t_L g540 ( 
.A(n_507),
.B(n_493),
.Y(n_540)
);

CKINVDCx14_ASAP7_75t_R g541 ( 
.A(n_514),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_514),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_485),
.B(n_489),
.Y(n_543)
);

NAND3xp33_ASAP7_75t_L g544 ( 
.A(n_487),
.B(n_537),
.C(n_483),
.Y(n_544)
);

AO31x2_ASAP7_75t_L g545 ( 
.A1(n_512),
.A2(n_515),
.A3(n_522),
.B(n_518),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_485),
.Y(n_546)
);

AO21x2_ASAP7_75t_L g547 ( 
.A1(n_488),
.A2(n_532),
.B(n_505),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_497),
.B(n_521),
.Y(n_548)
);

AO222x2_ASAP7_75t_SL g549 ( 
.A1(n_528),
.A2(n_500),
.B1(n_483),
.B2(n_486),
.C1(n_520),
.C2(n_494),
.Y(n_549)
);

AOI21xp33_ASAP7_75t_L g550 ( 
.A1(n_529),
.A2(n_506),
.B(n_480),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_533),
.B(n_501),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_501),
.B(n_491),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_530),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_517),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g555 ( 
.A(n_526),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_495),
.Y(n_556)
);

AOI21xp33_ASAP7_75t_L g557 ( 
.A1(n_529),
.A2(n_520),
.B(n_516),
.Y(n_557)
);

OA21x2_ASAP7_75t_L g558 ( 
.A1(n_502),
.A2(n_484),
.B(n_498),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_531),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_527),
.Y(n_560)
);

OA21x2_ASAP7_75t_L g561 ( 
.A1(n_536),
.A2(n_511),
.B(n_519),
.Y(n_561)
);

OAI21x1_ASAP7_75t_L g562 ( 
.A1(n_504),
.A2(n_508),
.B(n_523),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_496),
.A2(n_525),
.B1(n_509),
.B2(n_492),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_535),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_535),
.Y(n_565)
);

OAI21x1_ASAP7_75t_L g566 ( 
.A1(n_499),
.A2(n_510),
.B(n_513),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_527),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_503),
.A2(n_524),
.B1(n_535),
.B2(n_490),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_503),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_524),
.B(n_527),
.Y(n_570)
);

A2O1A1Ixp33_ASAP7_75t_L g571 ( 
.A1(n_524),
.A2(n_487),
.B(n_537),
.C(n_483),
.Y(n_571)
);

OAI21x1_ASAP7_75t_L g572 ( 
.A1(n_534),
.A2(n_484),
.B(n_536),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_534),
.B(n_487),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_532),
.A2(n_496),
.B(n_511),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_482),
.B(n_485),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_484),
.A2(n_536),
.B(n_502),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_481),
.Y(n_577)
);

AO21x1_ASAP7_75t_L g578 ( 
.A1(n_483),
.A2(n_515),
.B(n_512),
.Y(n_578)
);

AO21x2_ASAP7_75t_L g579 ( 
.A1(n_488),
.A2(n_515),
.B(n_512),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_482),
.Y(n_580)
);

CKINVDCx11_ASAP7_75t_R g581 ( 
.A(n_481),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_487),
.B(n_364),
.Y(n_582)
);

NOR2x1_ASAP7_75t_L g583 ( 
.A(n_509),
.B(n_512),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_487),
.B(n_364),
.Y(n_584)
);

AOI22x1_ASAP7_75t_L g585 ( 
.A1(n_488),
.A2(n_446),
.B1(n_531),
.B2(n_522),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_582),
.B(n_584),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_559),
.B(n_551),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_564),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_565),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_548),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_553),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_552),
.Y(n_592)
);

AO21x2_ASAP7_75t_L g593 ( 
.A1(n_578),
.A2(n_571),
.B(n_572),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_573),
.Y(n_594)
);

OAI211xp5_ASAP7_75t_L g595 ( 
.A1(n_544),
.A2(n_557),
.B(n_550),
.C(n_549),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_569),
.Y(n_596)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_562),
.A2(n_576),
.B(n_566),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_567),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_555),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_544),
.B(n_556),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_569),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_549),
.B(n_540),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_581),
.Y(n_603)
);

OA21x2_ASAP7_75t_L g604 ( 
.A1(n_560),
.A2(n_568),
.B(n_574),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_548),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_543),
.Y(n_606)
);

CKINVDCx11_ASAP7_75t_R g607 ( 
.A(n_538),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_570),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_543),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_570),
.Y(n_610)
);

OAI21x1_ASAP7_75t_L g611 ( 
.A1(n_585),
.A2(n_558),
.B(n_568),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_546),
.B(n_575),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_570),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_569),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_580),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_539),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_539),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_575),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_554),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_540),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_540),
.Y(n_621)
);

OAI21x1_ASAP7_75t_L g622 ( 
.A1(n_561),
.A2(n_583),
.B(n_563),
.Y(n_622)
);

OR2x6_ASAP7_75t_L g623 ( 
.A(n_542),
.B(n_583),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_545),
.B(n_541),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_545),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_608),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_600),
.A2(n_579),
.B1(n_547),
.B2(n_538),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_594),
.B(n_579),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_615),
.Y(n_629)
);

AO21x2_ASAP7_75t_L g630 ( 
.A1(n_611),
.A2(n_547),
.B(n_577),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_592),
.B(n_600),
.Y(n_631)
);

NAND2x1_ASAP7_75t_L g632 ( 
.A(n_598),
.B(n_604),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_594),
.B(n_588),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_586),
.A2(n_595),
.B1(n_602),
.B2(n_587),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_621),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_587),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_592),
.B(n_602),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_602),
.B(n_586),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_602),
.A2(n_624),
.B1(n_607),
.B2(n_617),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_588),
.B(n_589),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_589),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_608),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_599),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_599),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_624),
.B(n_591),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_616),
.A2(n_618),
.B1(n_623),
.B2(n_605),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_621),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_590),
.B(n_612),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_612),
.B(n_591),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_613),
.Y(n_650)
);

AOI222xp33_ASAP7_75t_L g651 ( 
.A1(n_606),
.A2(n_609),
.B1(n_620),
.B2(n_619),
.C1(n_603),
.C2(n_613),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_596),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_610),
.B(n_625),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_623),
.B(n_604),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_623),
.B(n_610),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_623),
.B(n_596),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_625),
.Y(n_657)
);

INVx6_ASAP7_75t_L g658 ( 
.A(n_596),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_596),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_596),
.B(n_601),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_601),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_601),
.B(n_614),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_601),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_601),
.B(n_614),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_604),
.B(n_593),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_614),
.B(n_604),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_614),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_657),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_633),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_657),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_631),
.B(n_593),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_641),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_641),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_640),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_631),
.B(n_614),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_628),
.B(n_593),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_638),
.A2(n_603),
.B1(n_622),
.B2(n_611),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_640),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_629),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_645),
.B(n_622),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_667),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_655),
.B(n_597),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_636),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_633),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_628),
.B(n_597),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_655),
.B(n_637),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_643),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_656),
.B(n_626),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_637),
.B(n_666),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_666),
.B(n_653),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_656),
.B(n_626),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_634),
.B(n_649),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_653),
.B(n_638),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_648),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_634),
.B(n_647),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_632),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_694),
.B(n_644),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_690),
.B(n_654),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_686),
.B(n_650),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_690),
.B(n_654),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_672),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_672),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_676),
.B(n_665),
.Y(n_703)
);

NOR3xp33_ASAP7_75t_L g704 ( 
.A(n_692),
.B(n_660),
.C(n_663),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_673),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_689),
.B(n_650),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_673),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_689),
.B(n_630),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_676),
.B(n_665),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_668),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_683),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_SL g712 ( 
.A1(n_695),
.A2(n_639),
.B(n_651),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_679),
.B(n_644),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_693),
.B(n_627),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_670),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_687),
.Y(n_716)
);

NOR2x1_ASAP7_75t_L g717 ( 
.A(n_681),
.B(n_643),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_686),
.B(n_626),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_674),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_671),
.B(n_630),
.Y(n_720)
);

NOR2xp67_ASAP7_75t_L g721 ( 
.A(n_696),
.B(n_642),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_674),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_678),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_678),
.Y(n_724)
);

AOI221xp5_ASAP7_75t_L g725 ( 
.A1(n_712),
.A2(n_684),
.B1(n_669),
.B2(n_671),
.C(n_677),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_701),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_708),
.B(n_680),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_698),
.B(n_685),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_718),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_703),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_701),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_702),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_702),
.Y(n_733)
);

NAND2x1_ASAP7_75t_L g734 ( 
.A(n_717),
.B(n_696),
.Y(n_734)
);

OR2x6_ASAP7_75t_L g735 ( 
.A(n_721),
.B(n_632),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_698),
.B(n_685),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_705),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_711),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_706),
.B(n_693),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_700),
.B(n_680),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_705),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_706),
.B(n_682),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_707),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_708),
.B(n_700),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_707),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_715),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_726),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_728),
.B(n_709),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_L g749 ( 
.A1(n_725),
.A2(n_704),
.B(n_651),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_744),
.B(n_699),
.Y(n_750)
);

NAND3xp33_ASAP7_75t_L g751 ( 
.A(n_725),
.B(n_738),
.C(n_697),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_731),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_730),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_L g754 ( 
.A1(n_734),
.A2(n_714),
.B1(n_709),
.B2(n_703),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_729),
.B(n_699),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_729),
.B(n_713),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_733),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_732),
.Y(n_758)
);

NOR3xp33_ASAP7_75t_L g759 ( 
.A(n_730),
.B(n_675),
.C(n_642),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_744),
.B(n_727),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_737),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_733),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_747),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_751),
.B(n_736),
.Y(n_764)
);

INVxp67_ASAP7_75t_SL g765 ( 
.A(n_754),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_748),
.B(n_740),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_749),
.A2(n_691),
.B1(n_688),
.B2(n_720),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_749),
.A2(n_716),
.B(n_719),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_757),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_768),
.A2(n_756),
.B(n_759),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_768),
.A2(n_753),
.B(n_735),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_764),
.B(n_760),
.Y(n_772)
);

AOI322xp5_ASAP7_75t_L g773 ( 
.A1(n_765),
.A2(n_753),
.A3(n_760),
.B1(n_727),
.B2(n_720),
.C1(n_742),
.C2(n_739),
.Y(n_773)
);

AOI31xp33_ASAP7_75t_L g774 ( 
.A1(n_767),
.A2(n_755),
.A3(n_750),
.B(n_761),
.Y(n_774)
);

OAI221xp5_ASAP7_75t_L g775 ( 
.A1(n_763),
.A2(n_758),
.B1(n_752),
.B2(n_762),
.C(n_741),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_769),
.Y(n_776)
);

OAI211xp5_ASAP7_75t_L g777 ( 
.A1(n_773),
.A2(n_646),
.B(n_722),
.C(n_723),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_L g778 ( 
.A(n_771),
.B(n_766),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_772),
.B(n_770),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_774),
.A2(n_775),
.B(n_776),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_770),
.B(n_755),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_777),
.Y(n_782)
);

NOR3xp33_ASAP7_75t_L g783 ( 
.A(n_779),
.B(n_781),
.C(n_778),
.Y(n_783)
);

NAND4xp75_ASAP7_75t_L g784 ( 
.A(n_782),
.B(n_780),
.C(n_662),
.D(n_724),
.Y(n_784)
);

NOR3xp33_ASAP7_75t_L g785 ( 
.A(n_783),
.B(n_663),
.C(n_661),
.Y(n_785)
);

OAI22xp33_ASAP7_75t_SL g786 ( 
.A1(n_782),
.A2(n_735),
.B1(n_743),
.B2(n_746),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_784),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_785),
.B(n_699),
.Y(n_788)
);

XNOR2xp5_ASAP7_75t_L g789 ( 
.A(n_786),
.B(n_647),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_784),
.Y(n_790)
);

INVxp33_ASAP7_75t_L g791 ( 
.A(n_785),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_787),
.A2(n_735),
.B1(n_718),
.B2(n_647),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_790),
.B(n_788),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_789),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_791),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_787),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_L g797 ( 
.A(n_789),
.B(n_745),
.Y(n_797)
);

NOR3xp33_ASAP7_75t_L g798 ( 
.A(n_787),
.B(n_663),
.C(n_661),
.Y(n_798)
);

INVx3_ASAP7_75t_SL g799 ( 
.A(n_795),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_796),
.A2(n_792),
.B1(n_794),
.B2(n_793),
.Y(n_800)
);

OAI22x1_ASAP7_75t_L g801 ( 
.A1(n_798),
.A2(n_664),
.B1(n_659),
.B2(n_662),
.Y(n_801)
);

AO22x2_ASAP7_75t_L g802 ( 
.A1(n_797),
.A2(n_664),
.B1(n_745),
.B2(n_635),
.Y(n_802)
);

XNOR2x1_ASAP7_75t_L g803 ( 
.A(n_793),
.B(n_664),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_799),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_803),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_800),
.A2(n_802),
.B1(n_801),
.B2(n_635),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_799),
.Y(n_807)
);

OAI21x1_ASAP7_75t_SL g808 ( 
.A1(n_804),
.A2(n_715),
.B(n_710),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_807),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_805),
.B(n_806),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_804),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_809),
.A2(n_658),
.B1(n_664),
.B2(n_635),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_811),
.A2(n_810),
.B1(n_808),
.B2(n_681),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_813),
.A2(n_630),
.B(n_661),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_814),
.B(n_812),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_815),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_816),
.A2(n_658),
.B1(n_667),
.B2(n_652),
.Y(n_817)
);


endmodule