module real_jpeg_26708_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_286, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_286;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_249;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_262;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_278;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_256;
wire n_274;
wire n_101;
wire n_182;
wire n_253;
wire n_273;
wire n_96;
wire n_269;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_SL g65 ( 
.A(n_0),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_1),
.Y(n_92)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_1),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_4),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_4),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_4),
.A2(n_20),
.B1(n_63),
.B2(n_64),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_4),
.A2(n_20),
.B1(n_42),
.B2(n_44),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_6),
.A2(n_18),
.B1(n_19),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_52),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_6),
.A2(n_52),
.B1(n_63),
.B2(n_64),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_6),
.A2(n_42),
.B1(n_44),
.B2(n_52),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_7),
.A2(n_18),
.B1(n_19),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_7),
.A2(n_29),
.B1(n_42),
.B2(n_44),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_7),
.A2(n_29),
.B1(n_63),
.B2(n_64),
.Y(n_201)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_8),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_11),
.A2(n_18),
.B1(n_19),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_36),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_SL g87 ( 
.A1(n_11),
.A2(n_24),
.B(n_26),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_11),
.A2(n_36),
.B1(n_63),
.B2(n_64),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_11),
.A2(n_36),
.B1(n_42),
.B2(n_44),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_11),
.B(n_25),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_11),
.A2(n_42),
.B(n_141),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g163 ( 
.A1(n_11),
.A2(n_60),
.B(n_64),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_11),
.B(n_41),
.Y(n_166)
);

AO21x1_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_278),
.B(n_282),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_67),
.B(n_277),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_30),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_15),
.B(n_30),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_15),
.B(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_15),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_21),
.B1(n_25),
.B2(n_28),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_17),
.A2(n_33),
.B(n_34),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_19),
.A2(n_23),
.B(n_36),
.C(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_21),
.A2(n_25),
.B1(n_35),
.B2(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_21),
.B(n_25),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx5_ASAP7_75t_SL g27 ( 
.A(n_26),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_26),
.A2(n_36),
.B(n_43),
.C(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_28),
.B(n_281),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_31),
.B(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_31),
.B(n_275),
.Y(n_276)
);

FAx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_37),
.CI(n_48),
.CON(n_31),
.SN(n_31)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_33),
.A2(n_34),
.B(n_51),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_35),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_36),
.A2(n_42),
.B(n_61),
.C(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_36),
.B(n_94),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_36),
.B(n_62),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_41),
.B1(n_45),
.B2(n_54),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_40),
.B(n_79),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_41),
.A2(n_54),
.B(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_44),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_80),
.Y(n_99)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_47),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.C(n_55),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_76),
.B1(n_82),
.B2(n_83),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_49),
.B(n_83),
.C(n_84),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_49),
.A2(n_82),
.B1(n_98),
.B2(n_122),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_49),
.B(n_122),
.C(n_217),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_49),
.A2(n_82),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_53),
.A2(n_55),
.B1(n_256),
.B2(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_53),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_55),
.A2(n_253),
.B1(n_254),
.B2(n_256),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_55),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_66),
.Y(n_55)
);

INVxp33_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_62),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_103),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_58),
.A2(n_62),
.B1(n_103),
.B2(n_110),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_58),
.A2(n_62),
.B1(n_66),
.B2(n_222),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_62),
.A2(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_63),
.B(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_91),
.Y(n_90)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_274),
.B(n_276),
.Y(n_67)
);

OAI321xp33_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_248),
.A3(n_267),
.B1(n_272),
.B2(n_273),
.C(n_286),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_230),
.B(n_247),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_211),
.B(n_229),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_133),
.B(n_194),
.C(n_210),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_119),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_73),
.B(n_119),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_95),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_74),
.B(n_96),
.C(n_106),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_84),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_76),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_128),
.C(n_131),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_76),
.A2(n_83),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_76),
.A2(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_76),
.B(n_236),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_81),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_86),
.B1(n_88),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_88),
.A2(n_126),
.B1(n_165),
.B2(n_168),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_88),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_88),
.B(n_178),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_88),
.B(n_155),
.C(n_167),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_116),
.B(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_90),
.B(n_91),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_90),
.A2(n_94),
.B1(n_115),
.B2(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_94),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_105),
.B2(n_106),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.C(n_104),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_100),
.B1(n_101),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_98),
.A2(n_107),
.B1(n_108),
.B2(n_122),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_99),
.Y(n_255)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_104),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_104),
.A2(n_123),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_104),
.A2(n_123),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_104),
.A2(n_123),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_104),
.B(n_254),
.C(n_256),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_104),
.B(n_261),
.C(n_266),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_113),
.B2(n_114),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_107),
.A2(n_108),
.B1(n_162),
.B2(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_107),
.B(n_114),
.Y(n_204)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_122),
.C(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_108),
.B(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_111),
.B(n_112),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_112),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_125),
.C(n_127),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_120),
.B(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_121),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_123),
.B(n_204),
.C(n_206),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_125),
.B(n_127),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_131),
.B1(n_132),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_128),
.B(n_175),
.Y(n_174)
);

INVx5_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_193),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_188),
.B(n_192),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_158),
.B(n_187),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_146),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_146),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_139),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_145),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_152),
.B2(n_153),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_155),
.C(n_156),
.Y(n_189)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_149),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_150),
.B(n_171),
.Y(n_180)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_154),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_155),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_157),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_155),
.A2(n_157),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_155),
.B(n_200),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_182),
.B(n_186),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_169),
.B(n_181),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_164),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_162),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_165),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_166),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_173),
.B(n_180),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_177),
.B(n_179),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_184),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_190),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_195),
.B(n_196),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_208),
.B2(n_209),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_203),
.C(n_209),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_200),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_208),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_212),
.B(n_213),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_228),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_219),
.B2(n_220),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_220),
.C(n_228),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_221),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_225),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_224),
.A2(n_225),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g258 ( 
.A1(n_225),
.A2(n_239),
.B(n_241),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_232),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_245),
.B2(n_246),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_238),
.C(n_246),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_250),
.C(n_257),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_250),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_244),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_245),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_259),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_259),
.Y(n_273)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_257),
.A2(n_258),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_266),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_270),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_284),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);


endmodule