module real_aes_9212_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_712;
wire n_183;
wire n_312;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g173 ( .A1(n_0), .A2(n_174), .B(n_177), .C(n_181), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_1), .B(n_165), .Y(n_184) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
NAND3xp33_ASAP7_75t_SL g723 ( .A(n_2), .B(n_439), .C(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_3), .B(n_175), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_4), .A2(n_134), .B(n_477), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_5), .A2(n_139), .B(n_142), .C(n_504), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_6), .A2(n_134), .B(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_7), .B(n_165), .Y(n_483) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_8), .A2(n_167), .B(n_242), .Y(n_241) );
AOI22xp33_ASAP7_75t_SL g101 ( .A1(n_9), .A2(n_102), .B1(n_719), .B2(n_720), .Y(n_101) );
AND2x6_ASAP7_75t_L g139 ( .A(n_10), .B(n_140), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_11), .A2(n_139), .B(n_142), .C(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g517 ( .A(n_12), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_13), .B(n_43), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_13), .B(n_43), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_14), .B(n_180), .Y(n_506) );
INVx1_ASAP7_75t_L g160 ( .A(n_15), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_16), .B(n_175), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_17), .A2(n_176), .B(n_537), .C(n_539), .Y(n_536) );
AOI222xp33_ASAP7_75t_SL g115 ( .A1(n_18), .A2(n_116), .B1(n_117), .B2(n_120), .C1(n_701), .C2(n_704), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_19), .B(n_165), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_20), .B(n_154), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g141 ( .A1(n_21), .A2(n_142), .B(n_145), .C(n_153), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_22), .A2(n_179), .B(n_235), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_23), .B(n_180), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g117 ( .A1(n_24), .A2(n_42), .B1(n_118), .B2(n_119), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_24), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_25), .B(n_180), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g451 ( .A(n_26), .Y(n_451) );
INVx1_ASAP7_75t_L g490 ( .A(n_27), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_28), .A2(n_142), .B(n_153), .C(n_245), .Y(n_244) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_29), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_30), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_31), .A2(n_78), .B1(n_714), .B2(n_715), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_31), .Y(n_715) );
INVx1_ASAP7_75t_L g468 ( .A(n_32), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_33), .A2(n_134), .B(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g137 ( .A(n_34), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_35), .A2(n_193), .B(n_194), .C(n_198), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_36), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_37), .A2(n_179), .B(n_480), .C(n_482), .Y(n_479) );
INVxp67_ASAP7_75t_L g469 ( .A(n_38), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_39), .B(n_247), .Y(n_246) );
CKINVDCx14_ASAP7_75t_R g478 ( .A(n_40), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_41), .A2(n_142), .B(n_153), .C(n_489), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_42), .Y(n_118) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_44), .A2(n_181), .B(n_515), .C(n_516), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_45), .B(n_133), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_46), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_47), .B(n_175), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_48), .B(n_134), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_49), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_50), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_51), .A2(n_193), .B(n_198), .C(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g178 ( .A(n_52), .Y(n_178) );
INVx1_ASAP7_75t_L g221 ( .A(n_53), .Y(n_221) );
INVx1_ASAP7_75t_L g523 ( .A(n_54), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_55), .B(n_134), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_56), .Y(n_162) );
CKINVDCx14_ASAP7_75t_R g513 ( .A(n_57), .Y(n_513) );
INVx1_ASAP7_75t_L g140 ( .A(n_58), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_59), .B(n_134), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_60), .B(n_165), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_61), .A2(n_152), .B(n_208), .C(n_210), .Y(n_207) );
INVx1_ASAP7_75t_L g159 ( .A(n_62), .Y(n_159) );
INVx1_ASAP7_75t_SL g481 ( .A(n_63), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_64), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_65), .B(n_175), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_66), .B(n_165), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_67), .B(n_176), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_68), .Y(n_108) );
INVx1_ASAP7_75t_L g454 ( .A(n_69), .Y(n_454) );
CKINVDCx16_ASAP7_75t_R g171 ( .A(n_70), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_71), .B(n_147), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_72), .A2(n_142), .B(n_198), .C(n_261), .Y(n_260) );
CKINVDCx16_ASAP7_75t_R g206 ( .A(n_73), .Y(n_206) );
INVx1_ASAP7_75t_L g726 ( .A(n_74), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_75), .A2(n_134), .B(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_76), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_77), .A2(n_134), .B(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_78), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_79), .A2(n_133), .B(n_464), .Y(n_463) );
CKINVDCx16_ASAP7_75t_R g487 ( .A(n_80), .Y(n_487) );
INVx1_ASAP7_75t_L g535 ( .A(n_81), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_82), .B(n_150), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_83), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_84), .A2(n_134), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g538 ( .A(n_85), .Y(n_538) );
INVx2_ASAP7_75t_L g157 ( .A(n_86), .Y(n_157) );
INVx1_ASAP7_75t_L g505 ( .A(n_87), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_88), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_89), .B(n_180), .Y(n_233) );
OR2x2_ASAP7_75t_L g110 ( .A(n_90), .B(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g123 ( .A(n_90), .B(n_112), .Y(n_123) );
INVx2_ASAP7_75t_L g439 ( .A(n_90), .Y(n_439) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_91), .A2(n_142), .B(n_198), .C(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_92), .B(n_134), .Y(n_191) );
INVx1_ASAP7_75t_L g195 ( .A(n_93), .Y(n_195) );
INVxp67_ASAP7_75t_L g211 ( .A(n_94), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_95), .B(n_167), .Y(n_518) );
INVx1_ASAP7_75t_L g228 ( .A(n_96), .Y(n_228) );
INVx1_ASAP7_75t_L g262 ( .A(n_97), .Y(n_262) );
INVx2_ASAP7_75t_L g526 ( .A(n_98), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_99), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g223 ( .A(n_100), .B(n_156), .Y(n_223) );
AOI22x1_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_115), .B1(n_709), .B2(n_711), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
BUFx2_ASAP7_75t_L g710 ( .A(n_105), .Y(n_710) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_107), .A2(n_712), .B(n_718), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_110), .Y(n_718) );
NOR2x2_ASAP7_75t_L g703 ( .A(n_111), .B(n_439), .Y(n_703) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g438 ( .A(n_112), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI22xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_124), .B1(n_438), .B2(n_440), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g705 ( .A(n_122), .Y(n_705) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g712 ( .A1(n_124), .A2(n_713), .B1(n_716), .B2(n_717), .Y(n_712) );
INVx1_ASAP7_75t_L g716 ( .A(n_124), .Y(n_716) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_SL g704 ( .A1(n_125), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_704) );
AND2x2_ASAP7_75t_SL g125 ( .A(n_126), .B(n_374), .Y(n_125) );
NOR5xp2_ASAP7_75t_L g126 ( .A(n_127), .B(n_305), .C(n_334), .D(n_354), .E(n_361), .Y(n_126) );
OAI211xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_185), .B(n_249), .C(n_292), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_129), .A2(n_377), .B1(n_379), .B2(n_380), .Y(n_376) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_164), .Y(n_129) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_130), .Y(n_252) );
AND2x4_ASAP7_75t_L g285 ( .A(n_130), .B(n_286), .Y(n_285) );
INVx5_ASAP7_75t_L g303 ( .A(n_130), .Y(n_303) );
AND2x2_ASAP7_75t_L g312 ( .A(n_130), .B(n_304), .Y(n_312) );
AND2x2_ASAP7_75t_L g324 ( .A(n_130), .B(n_189), .Y(n_324) );
AND2x2_ASAP7_75t_L g420 ( .A(n_130), .B(n_288), .Y(n_420) );
OR2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_161), .Y(n_130) );
AOI21xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_141), .B(n_154), .Y(n_131) );
BUFx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_139), .Y(n_134) );
NAND2x1p5_ASAP7_75t_L g229 ( .A(n_135), .B(n_139), .Y(n_229) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
INVx1_ASAP7_75t_L g152 ( .A(n_136), .Y(n_152) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g143 ( .A(n_137), .Y(n_143) );
INVx1_ASAP7_75t_L g236 ( .A(n_137), .Y(n_236) );
INVx1_ASAP7_75t_L g144 ( .A(n_138), .Y(n_144) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_138), .Y(n_148) );
INVx3_ASAP7_75t_L g176 ( .A(n_138), .Y(n_176) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_138), .Y(n_180) );
INVx1_ASAP7_75t_L g247 ( .A(n_138), .Y(n_247) );
BUFx3_ASAP7_75t_L g153 ( .A(n_139), .Y(n_153) );
INVx4_ASAP7_75t_SL g183 ( .A(n_139), .Y(n_183) );
INVx5_ASAP7_75t_L g172 ( .A(n_142), .Y(n_172) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
BUFx3_ASAP7_75t_L g182 ( .A(n_143), .Y(n_182) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_143), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_149), .B(n_151), .Y(n_145) );
INVx2_ASAP7_75t_L g150 ( .A(n_147), .Y(n_150) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx4_ASAP7_75t_L g209 ( .A(n_148), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_150), .A2(n_195), .B(n_196), .C(n_197), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_150), .A2(n_197), .B(n_221), .C(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g453 ( .A1(n_150), .A2(n_454), .B(n_455), .C(n_456), .Y(n_453) );
O2A1O1Ixp5_ASAP7_75t_L g504 ( .A1(n_150), .A2(n_456), .B(n_505), .C(n_506), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_151), .A2(n_175), .B(n_490), .C(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_152), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_155), .B(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g163 ( .A(n_156), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_156), .A2(n_191), .B(n_192), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_156), .A2(n_218), .B(n_219), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_156), .A2(n_229), .B(n_487), .C(n_488), .Y(n_486) );
OA21x2_ASAP7_75t_L g510 ( .A1(n_156), .A2(n_511), .B(n_518), .Y(n_510) );
AND2x2_ASAP7_75t_SL g156 ( .A(n_157), .B(n_158), .Y(n_156) );
AND2x2_ASAP7_75t_L g168 ( .A(n_157), .B(n_158), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_163), .A2(n_501), .B(n_507), .Y(n_500) );
INVx2_ASAP7_75t_L g286 ( .A(n_164), .Y(n_286) );
AND2x2_ASAP7_75t_L g304 ( .A(n_164), .B(n_258), .Y(n_304) );
AND2x2_ASAP7_75t_L g323 ( .A(n_164), .B(n_257), .Y(n_323) );
AND2x2_ASAP7_75t_L g363 ( .A(n_164), .B(n_303), .Y(n_363) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_169), .B(n_184), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_166), .B(n_200), .Y(n_199) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_166), .A2(n_227), .B(n_237), .Y(n_226) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_166), .A2(n_259), .B(n_267), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_166), .B(n_268), .Y(n_267) );
AO21x2_ASAP7_75t_L g449 ( .A1(n_166), .A2(n_450), .B(n_457), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_166), .B(n_493), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_166), .B(n_508), .Y(n_507) );
INVx4_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_167), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_167), .A2(n_243), .B(n_244), .Y(n_242) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g239 ( .A(n_168), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_SL g170 ( .A1(n_171), .A2(n_172), .B(n_173), .C(n_183), .Y(n_170) );
INVx2_ASAP7_75t_L g193 ( .A(n_172), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_172), .A2(n_183), .B(n_206), .C(n_207), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_SL g464 ( .A1(n_172), .A2(n_183), .B(n_465), .C(n_466), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_172), .A2(n_183), .B(n_478), .C(n_479), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_SL g512 ( .A1(n_172), .A2(n_183), .B(n_513), .C(n_514), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_SL g522 ( .A1(n_172), .A2(n_183), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_SL g534 ( .A1(n_172), .A2(n_183), .B(n_535), .C(n_536), .Y(n_534) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_175), .B(n_211), .Y(n_210) );
OAI22xp33_ASAP7_75t_L g467 ( .A1(n_175), .A2(n_209), .B1(n_468), .B2(n_469), .Y(n_467) );
INVx5_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_176), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_179), .B(n_481), .Y(n_480) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g515 ( .A(n_180), .Y(n_515) );
INVx2_ASAP7_75t_L g456 ( .A(n_181), .Y(n_456) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_182), .Y(n_197) );
INVx1_ASAP7_75t_L g539 ( .A(n_182), .Y(n_539) );
INVx1_ASAP7_75t_L g198 ( .A(n_183), .Y(n_198) );
INVxp67_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_187), .B(n_213), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AOI322xp5_ASAP7_75t_L g422 ( .A1(n_188), .A2(n_224), .A3(n_277), .B1(n_285), .B2(n_339), .C1(n_423), .C2(n_426), .Y(n_422) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_201), .Y(n_188) );
INVx5_ASAP7_75t_L g254 ( .A(n_189), .Y(n_254) );
AND2x2_ASAP7_75t_L g271 ( .A(n_189), .B(n_256), .Y(n_271) );
BUFx2_ASAP7_75t_L g349 ( .A(n_189), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_189), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g426 ( .A(n_189), .B(n_333), .Y(n_426) );
OR2x6_ASAP7_75t_L g189 ( .A(n_190), .B(n_199), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_201), .B(n_215), .Y(n_280) );
INVx1_ASAP7_75t_L g307 ( .A(n_201), .Y(n_307) );
AND2x2_ASAP7_75t_L g320 ( .A(n_201), .B(n_240), .Y(n_320) );
AND2x2_ASAP7_75t_L g421 ( .A(n_201), .B(n_339), .Y(n_421) );
INVx3_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
OR2x2_ASAP7_75t_L g275 ( .A(n_202), .B(n_215), .Y(n_275) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_202), .Y(n_283) );
OR2x2_ASAP7_75t_L g290 ( .A(n_202), .B(n_240), .Y(n_290) );
AND2x2_ASAP7_75t_L g300 ( .A(n_202), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_202), .B(n_226), .Y(n_329) );
INVxp67_ASAP7_75t_L g353 ( .A(n_202), .Y(n_353) );
AND2x2_ASAP7_75t_L g360 ( .A(n_202), .B(n_224), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_202), .B(n_240), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_202), .B(n_225), .Y(n_386) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_212), .Y(n_202) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_203), .A2(n_476), .B(n_483), .Y(n_475) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_203), .A2(n_521), .B(n_527), .Y(n_520) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_203), .A2(n_533), .B(n_540), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_208), .A2(n_262), .B(n_263), .C(n_264), .Y(n_261) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_209), .B(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_209), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_224), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_215), .B(n_241), .Y(n_330) );
OR2x2_ASAP7_75t_L g352 ( .A(n_215), .B(n_225), .Y(n_352) );
AND2x2_ASAP7_75t_L g365 ( .A(n_215), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_215), .B(n_320), .Y(n_371) );
OAI211xp5_ASAP7_75t_SL g375 ( .A1(n_215), .A2(n_376), .B(n_381), .C(n_390), .Y(n_375) );
AND2x2_ASAP7_75t_L g436 ( .A(n_215), .B(n_240), .Y(n_436) );
INVx5_ASAP7_75t_SL g215 ( .A(n_216), .Y(n_215) );
OR2x2_ASAP7_75t_L g289 ( .A(n_216), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_216), .B(n_295), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_216), .B(n_284), .Y(n_296) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_216), .Y(n_298) );
OR2x2_ASAP7_75t_L g309 ( .A(n_216), .B(n_225), .Y(n_309) );
AND2x2_ASAP7_75t_SL g314 ( .A(n_216), .B(n_300), .Y(n_314) );
AND2x2_ASAP7_75t_L g339 ( .A(n_216), .B(n_225), .Y(n_339) );
AND2x2_ASAP7_75t_L g359 ( .A(n_216), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g397 ( .A(n_216), .B(n_224), .Y(n_397) );
OR2x2_ASAP7_75t_L g400 ( .A(n_216), .B(n_386), .Y(n_400) );
OR2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_223), .Y(n_216) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_240), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g343 ( .A1(n_225), .A2(n_344), .B(n_347), .C(n_353), .Y(n_343) );
INVx5_ASAP7_75t_SL g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_226), .B(n_240), .Y(n_274) );
AND2x2_ASAP7_75t_L g278 ( .A(n_226), .B(n_241), .Y(n_278) );
OR2x2_ASAP7_75t_L g284 ( .A(n_226), .B(n_240), .Y(n_284) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_230), .Y(n_227) );
OAI21xp5_ASAP7_75t_L g450 ( .A1(n_229), .A2(n_451), .B(n_452), .Y(n_450) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_229), .A2(n_502), .B(n_503), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_234), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_234), .A2(n_246), .B(n_248), .Y(n_245) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx2_ASAP7_75t_L g461 ( .A(n_239), .Y(n_461) );
INVx1_ASAP7_75t_SL g301 ( .A(n_240), .Y(n_301) );
OR2x2_ASAP7_75t_L g429 ( .A(n_240), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_269), .B(n_272), .C(n_281), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AOI31xp33_ASAP7_75t_L g354 ( .A1(n_251), .A2(n_355), .A3(n_357), .B(n_358), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_252), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_253), .B(n_285), .Y(n_291) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_254), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g311 ( .A(n_254), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g316 ( .A(n_254), .B(n_286), .Y(n_316) );
AND2x2_ASAP7_75t_L g326 ( .A(n_254), .B(n_285), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_254), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g346 ( .A(n_254), .B(n_303), .Y(n_346) );
AND2x2_ASAP7_75t_L g351 ( .A(n_254), .B(n_323), .Y(n_351) );
OR2x2_ASAP7_75t_L g370 ( .A(n_254), .B(n_256), .Y(n_370) );
OR2x2_ASAP7_75t_L g372 ( .A(n_254), .B(n_373), .Y(n_372) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_254), .Y(n_419) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g319 ( .A(n_256), .B(n_286), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_256), .B(n_303), .Y(n_342) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
BUFx2_ASAP7_75t_L g288 ( .A(n_258), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_266), .Y(n_259) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx3_ASAP7_75t_L g482 ( .A(n_265), .Y(n_482) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g379 ( .A(n_271), .B(n_303), .Y(n_379) );
AOI322xp5_ASAP7_75t_L g381 ( .A1(n_271), .A2(n_285), .A3(n_323), .B1(n_382), .B2(n_383), .C1(n_384), .C2(n_387), .Y(n_381) );
INVx1_ASAP7_75t_L g389 ( .A(n_271), .Y(n_389) );
NAND2xp33_ASAP7_75t_L g272 ( .A(n_273), .B(n_276), .Y(n_272) );
INVx1_ASAP7_75t_SL g383 ( .A(n_273), .Y(n_383) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
OR2x2_ASAP7_75t_L g335 ( .A(n_274), .B(n_280), .Y(n_335) );
INVx1_ASAP7_75t_L g366 ( .A(n_274), .Y(n_366) );
INVx2_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OAI32xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_285), .A3(n_287), .B1(n_289), .B2(n_291), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
AOI21xp33_ASAP7_75t_SL g321 ( .A1(n_284), .A2(n_299), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g336 ( .A(n_285), .Y(n_336) );
AND2x4_ASAP7_75t_L g333 ( .A(n_286), .B(n_303), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_286), .B(n_369), .Y(n_368) );
AOI322xp5_ASAP7_75t_L g398 ( .A1(n_287), .A2(n_314), .A3(n_333), .B1(n_366), .B2(n_399), .C1(n_401), .C2(n_402), .Y(n_398) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_287), .A2(n_364), .B1(n_428), .B2(n_429), .C(n_431), .Y(n_427) );
AND2x2_ASAP7_75t_L g315 ( .A(n_288), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g295 ( .A(n_290), .Y(n_295) );
OR2x2_ASAP7_75t_L g367 ( .A(n_290), .B(n_352), .Y(n_367) );
OAI31xp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_296), .A3(n_297), .B(n_302), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_293), .A2(n_326), .B1(n_327), .B2(n_331), .Y(n_325) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g338 ( .A(n_295), .B(n_339), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_297), .A2(n_338), .B1(n_391), .B2(n_394), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g380 ( .A(n_300), .B(n_349), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_300), .B(n_339), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_301), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g414 ( .A(n_301), .B(n_352), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_302), .A2(n_397), .B1(n_410), .B2(n_413), .Y(n_409) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx2_ASAP7_75t_L g318 ( .A(n_303), .Y(n_318) );
AND2x2_ASAP7_75t_L g401 ( .A(n_303), .B(n_323), .Y(n_401) );
OR2x2_ASAP7_75t_L g403 ( .A(n_303), .B(n_370), .Y(n_403) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_303), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_304), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_304), .B(n_349), .Y(n_357) );
OAI211xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_310), .B(n_313), .C(n_325), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AOI221xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B1(n_317), .B2(n_320), .C(n_321), .Y(n_313) );
INVxp67_ASAP7_75t_L g425 ( .A(n_316), .Y(n_425) );
INVx1_ASAP7_75t_L g392 ( .A(n_317), .Y(n_392) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x2_ASAP7_75t_L g356 ( .A(n_318), .B(n_323), .Y(n_356) );
INVx1_ASAP7_75t_L g373 ( .A(n_319), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_319), .B(n_346), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g388 ( .A(n_323), .Y(n_388) );
AND2x2_ASAP7_75t_L g394 ( .A(n_323), .B(n_349), .Y(n_394) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_SL g382 ( .A(n_330), .Y(n_382) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_333), .B(n_369), .Y(n_393) );
OAI221xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B1(n_337), .B2(n_340), .C(n_343), .Y(n_334) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g430 ( .A(n_339), .Y(n_430) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g348 ( .A(n_342), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_346), .B(n_405), .Y(n_404) );
AOI21xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_350), .B(n_352), .Y(n_347) );
OAI211xp5_ASAP7_75t_SL g395 ( .A1(n_350), .A2(n_396), .B(n_398), .C(n_404), .Y(n_395) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g407 ( .A(n_352), .Y(n_407) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI222xp33_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_364), .B1(n_367), .B2(n_368), .C1(n_371), .C2(n_372), .Y(n_361) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g437 ( .A(n_368), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_369), .B(n_412), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_369), .A2(n_416), .B1(n_418), .B2(n_421), .Y(n_415) );
INVx2_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
NOR4xp25_ASAP7_75t_L g374 ( .A(n_375), .B(n_395), .C(n_408), .D(n_427), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_377), .B(n_407), .Y(n_417) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g384 ( .A(n_382), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_385), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND3xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_415), .C(n_422), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx2_ASAP7_75t_L g424 ( .A(n_420), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
OAI21xp5_ASAP7_75t_SL g431 ( .A1(n_432), .A2(n_434), .B(n_437), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g708 ( .A(n_438), .Y(n_708) );
INVx2_ASAP7_75t_L g706 ( .A(n_440), .Y(n_706) );
OR2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_635), .Y(n_440) );
NAND5xp2_ASAP7_75t_L g441 ( .A(n_442), .B(n_564), .C(n_594), .D(n_615), .E(n_621), .Y(n_441) );
AOI221xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_497), .B1(n_528), .B2(n_530), .C(n_541), .Y(n_442) );
INVxp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_494), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_472), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_SL g615 ( .A1(n_447), .A2(n_484), .B(n_616), .C(n_619), .Y(n_615) );
AND2x2_ASAP7_75t_L g685 ( .A(n_447), .B(n_485), .Y(n_685) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_459), .Y(n_447) );
AND2x2_ASAP7_75t_L g543 ( .A(n_448), .B(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g547 ( .A(n_448), .B(n_544), .Y(n_547) );
OR2x2_ASAP7_75t_L g573 ( .A(n_448), .B(n_485), .Y(n_573) );
AND2x2_ASAP7_75t_L g575 ( .A(n_448), .B(n_475), .Y(n_575) );
AND2x2_ASAP7_75t_L g593 ( .A(n_448), .B(n_474), .Y(n_593) );
INVx1_ASAP7_75t_L g626 ( .A(n_448), .Y(n_626) );
INVx2_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
BUFx2_ASAP7_75t_L g496 ( .A(n_449), .Y(n_496) );
AND2x2_ASAP7_75t_L g529 ( .A(n_449), .B(n_475), .Y(n_529) );
AND2x2_ASAP7_75t_L g682 ( .A(n_449), .B(n_485), .Y(n_682) );
AND2x2_ASAP7_75t_L g563 ( .A(n_459), .B(n_473), .Y(n_563) );
OR2x2_ASAP7_75t_L g567 ( .A(n_459), .B(n_485), .Y(n_567) );
AND2x2_ASAP7_75t_L g592 ( .A(n_459), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_SL g639 ( .A(n_459), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_459), .B(n_601), .Y(n_687) );
AO21x2_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_462), .B(n_470), .Y(n_459) );
INVx1_ASAP7_75t_L g545 ( .A(n_460), .Y(n_545) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_463), .A2(n_471), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OAI322xp33_ASAP7_75t_L g688 ( .A1(n_472), .A2(n_624), .A3(n_647), .B1(n_668), .B2(n_689), .C1(n_691), .C2(n_692), .Y(n_688) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_473), .B(n_544), .Y(n_691) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_484), .Y(n_473) );
AND2x2_ASAP7_75t_L g495 ( .A(n_474), .B(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_L g560 ( .A(n_474), .B(n_485), .Y(n_560) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g601 ( .A(n_475), .B(n_485), .Y(n_601) );
AND2x2_ASAP7_75t_L g645 ( .A(n_475), .B(n_484), .Y(n_645) );
AND2x2_ASAP7_75t_L g528 ( .A(n_484), .B(n_529), .Y(n_528) );
OR2x2_ASAP7_75t_L g546 ( .A(n_484), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_484), .B(n_575), .Y(n_699) );
INVx3_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g494 ( .A(n_485), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_485), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g613 ( .A(n_485), .B(n_544), .Y(n_613) );
AND2x2_ASAP7_75t_L g640 ( .A(n_485), .B(n_575), .Y(n_640) );
OR2x2_ASAP7_75t_L g696 ( .A(n_485), .B(n_547), .Y(n_696) );
OR2x6_ASAP7_75t_L g485 ( .A(n_486), .B(n_492), .Y(n_485) );
INVx1_ASAP7_75t_SL g582 ( .A(n_494), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_495), .B(n_613), .Y(n_614) );
AND2x2_ASAP7_75t_L g648 ( .A(n_495), .B(n_638), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_495), .B(n_571), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_495), .B(n_693), .Y(n_692) );
OAI31xp33_ASAP7_75t_L g666 ( .A1(n_497), .A2(n_528), .A3(n_667), .B(n_669), .Y(n_666) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_509), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_498), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g649 ( .A(n_498), .B(n_584), .Y(n_649) );
OR2x2_ASAP7_75t_L g656 ( .A(n_498), .B(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g668 ( .A(n_498), .B(n_557), .Y(n_668) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
OR2x2_ASAP7_75t_L g602 ( .A(n_499), .B(n_603), .Y(n_602) );
BUFx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g530 ( .A(n_500), .B(n_531), .Y(n_530) );
INVx4_ASAP7_75t_L g551 ( .A(n_500), .Y(n_551) );
AND2x2_ASAP7_75t_L g588 ( .A(n_500), .B(n_532), .Y(n_588) );
AND2x2_ASAP7_75t_L g587 ( .A(n_509), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_SL g657 ( .A(n_509), .Y(n_657) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_519), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_510), .B(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g557 ( .A(n_510), .B(n_520), .Y(n_557) );
INVx2_ASAP7_75t_L g577 ( .A(n_510), .Y(n_577) );
AND2x2_ASAP7_75t_L g591 ( .A(n_510), .B(n_520), .Y(n_591) );
AND2x2_ASAP7_75t_L g598 ( .A(n_510), .B(n_554), .Y(n_598) );
BUFx3_ASAP7_75t_L g608 ( .A(n_510), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_510), .B(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g553 ( .A(n_519), .Y(n_553) );
AND2x2_ASAP7_75t_L g561 ( .A(n_519), .B(n_551), .Y(n_561) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g531 ( .A(n_520), .B(n_532), .Y(n_531) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_520), .Y(n_585) );
INVx2_ASAP7_75t_SL g568 ( .A(n_529), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_529), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_529), .B(n_638), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_530), .B(n_608), .Y(n_661) );
INVx1_ASAP7_75t_SL g695 ( .A(n_530), .Y(n_695) );
INVx1_ASAP7_75t_SL g603 ( .A(n_531), .Y(n_603) );
INVx1_ASAP7_75t_SL g554 ( .A(n_532), .Y(n_554) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_532), .Y(n_565) );
OR2x2_ASAP7_75t_L g576 ( .A(n_532), .B(n_551), .Y(n_576) );
AND2x2_ASAP7_75t_L g590 ( .A(n_532), .B(n_551), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_532), .B(n_580), .Y(n_642) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_546), .B(n_548), .C(n_559), .Y(n_541) );
AOI31xp33_ASAP7_75t_L g658 ( .A1(n_542), .A2(n_659), .A3(n_660), .B(n_661), .Y(n_658) );
AND2x2_ASAP7_75t_L g631 ( .A(n_543), .B(n_560), .Y(n_631) );
BUFx3_ASAP7_75t_L g571 ( .A(n_544), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_544), .B(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g607 ( .A(n_544), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_544), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_SL g562 ( .A(n_547), .Y(n_562) );
OAI222xp33_ASAP7_75t_L g671 ( .A1(n_547), .A2(n_672), .B1(n_675), .B2(n_676), .C1(n_677), .C2(n_678), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_555), .Y(n_548) );
INVx1_ASAP7_75t_L g677 ( .A(n_549), .Y(n_677) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_551), .B(n_554), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_551), .B(n_577), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_551), .B(n_552), .Y(n_647) );
INVx1_ASAP7_75t_L g698 ( .A(n_551), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_552), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g700 ( .A(n_552), .Y(n_700) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx2_ASAP7_75t_L g580 ( .A(n_553), .Y(n_580) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_554), .Y(n_623) );
AOI32xp33_ASAP7_75t_L g559 ( .A1(n_555), .A2(n_560), .A3(n_561), .B1(n_562), .B2(n_563), .Y(n_559) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_557), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g634 ( .A(n_557), .Y(n_634) );
OR2x2_ASAP7_75t_L g675 ( .A(n_557), .B(n_576), .Y(n_675) );
INVx1_ASAP7_75t_L g611 ( .A(n_558), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_560), .B(n_571), .Y(n_596) );
INVx3_ASAP7_75t_L g605 ( .A(n_560), .Y(n_605) );
AOI322xp5_ASAP7_75t_L g621 ( .A1(n_560), .A2(n_605), .A3(n_622), .B1(n_624), .B2(n_627), .C1(n_631), .C2(n_632), .Y(n_621) );
AND2x2_ASAP7_75t_L g597 ( .A(n_561), .B(n_598), .Y(n_597) );
INVxp67_ASAP7_75t_L g674 ( .A(n_561), .Y(n_674) );
A2O1A1O1Ixp25_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_566), .B(n_569), .C(n_577), .D(n_578), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_565), .B(n_608), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
OAI221xp5_ASAP7_75t_L g578 ( .A1(n_567), .A2(n_579), .B1(n_582), .B2(n_583), .C(n_586), .Y(n_578) );
INVx1_ASAP7_75t_SL g693 ( .A(n_567), .Y(n_693) );
AOI21xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_574), .B(n_576), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_571), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OAI221xp5_ASAP7_75t_SL g663 ( .A1(n_573), .A2(n_657), .B1(n_664), .B2(n_665), .C(n_666), .Y(n_663) );
OAI222xp33_ASAP7_75t_L g694 ( .A1(n_574), .A2(n_695), .B1(n_696), .B2(n_697), .C1(n_699), .C2(n_700), .Y(n_694) );
AND2x2_ASAP7_75t_L g652 ( .A(n_575), .B(n_638), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_575), .A2(n_590), .B(n_637), .Y(n_664) );
INVx1_ASAP7_75t_L g678 ( .A(n_575), .Y(n_678) );
INVx2_ASAP7_75t_SL g581 ( .A(n_576), .Y(n_581) );
AND2x2_ASAP7_75t_L g584 ( .A(n_577), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx1_ASAP7_75t_SL g618 ( .A(n_580), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_580), .B(n_590), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_581), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_581), .B(n_591), .Y(n_620) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OAI21xp5_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_589), .B(n_592), .Y(n_586) );
INVx1_ASAP7_75t_SL g604 ( .A(n_588), .Y(n_604) );
AND2x2_ASAP7_75t_L g651 ( .A(n_588), .B(n_634), .Y(n_651) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AND2x2_ASAP7_75t_L g690 ( .A(n_590), .B(n_608), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_591), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g676 ( .A(n_592), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_597), .B1(n_599), .B2(n_606), .C(n_609), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_602), .B1(n_604), .B2(n_605), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_603), .A2(n_610), .B1(n_612), .B2(n_614), .Y(n_609) );
OR2x2_ASAP7_75t_L g680 ( .A(n_604), .B(n_608), .Y(n_680) );
OR2x2_ASAP7_75t_L g683 ( .A(n_604), .B(n_618), .Y(n_683) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g679 ( .A1(n_625), .A2(n_680), .B1(n_681), .B2(n_683), .C(n_684), .Y(n_679) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVxp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND3xp33_ASAP7_75t_SL g635 ( .A(n_636), .B(n_650), .C(n_662), .Y(n_635) );
AOI222xp33_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_641), .B1(n_643), .B2(n_646), .C1(n_648), .C2(n_649), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_638), .B(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g660 ( .A(n_640), .Y(n_660) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B1(n_653), .B2(n_655), .C(n_658), .Y(n_650) );
INVx1_ASAP7_75t_L g665 ( .A(n_651), .Y(n_665) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI21xp33_ASAP7_75t_L g684 ( .A1(n_655), .A2(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
NOR5xp2_ASAP7_75t_L g662 ( .A(n_663), .B(n_671), .C(n_679), .D(n_688), .E(n_694), .Y(n_662) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
INVxp67_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g717 ( .A(n_713), .Y(n_717) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
endmodule