module fake_jpeg_7873_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_43),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_0),
.C(n_1),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_0),
.Y(n_61)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_62),
.Y(n_72)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_33),
.B1(n_22),
.B2(n_27),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_65),
.B1(n_17),
.B2(n_34),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_17),
.B(n_34),
.Y(n_84)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_33),
.B1(n_22),
.B2(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_31),
.Y(n_79)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_36),
.C(n_40),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_40),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_44),
.B1(n_25),
.B2(n_24),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_71),
.A2(n_76),
.B1(n_93),
.B2(n_96),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_44),
.B1(n_47),
.B2(n_46),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_73),
.A2(n_85),
.B1(n_88),
.B2(n_90),
.Y(n_110)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_77),
.Y(n_113)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_46),
.B(n_30),
.C(n_27),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_78),
.A2(n_66),
.B(n_23),
.C(n_32),
.Y(n_117)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_80),
.Y(n_116)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_23),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_47),
.B1(n_28),
.B2(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_87),
.Y(n_122)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_17),
.B1(n_24),
.B2(n_25),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_49),
.B1(n_69),
.B2(n_62),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_25),
.B1(n_24),
.B2(n_34),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_23),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_55),
.A2(n_28),
.B1(n_20),
.B2(n_29),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_18),
.B1(n_26),
.B2(n_20),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_68),
.B1(n_66),
.B2(n_26),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_55),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_98)
);

OAI22x1_ASAP7_75t_SL g105 ( 
.A1(n_98),
.A2(n_23),
.B1(n_26),
.B2(n_18),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_48),
.B(n_29),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_112),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_111),
.B1(n_118),
.B2(n_120),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_125),
.C(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_83),
.B(n_56),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_114),
.B(n_11),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_56),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_94),
.B(n_36),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_85),
.Y(n_134)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_123),
.B1(n_91),
.B2(n_35),
.Y(n_154)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_72),
.B(n_36),
.C(n_53),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_126),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_123),
.A2(n_72),
.B1(n_76),
.B2(n_78),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_128),
.A2(n_135),
.B1(n_148),
.B2(n_125),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_106),
.B(n_78),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_131),
.A2(n_134),
.B(n_140),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_41),
.C(n_37),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_110),
.B1(n_117),
.B2(n_121),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_141),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_75),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_115),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_105),
.A2(n_81),
.B1(n_75),
.B2(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_143),
.B(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_147),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_104),
.A2(n_77),
.B1(n_86),
.B2(n_82),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_115),
.A2(n_81),
.B1(n_92),
.B2(n_74),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_102),
.A2(n_92),
.B1(n_94),
.B2(n_26),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_150),
.B(n_35),
.Y(n_175)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_153),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_152),
.B(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_112),
.B(n_10),
.Y(n_156)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_159),
.B1(n_174),
.B2(n_179),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_145),
.A2(n_109),
.B1(n_101),
.B2(n_116),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_169),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_127),
.A2(n_119),
.B1(n_126),
.B2(n_124),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_162),
.A2(n_130),
.B1(n_139),
.B2(n_142),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_100),
.B(n_32),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_163),
.A2(n_4),
.B(n_5),
.Y(n_214)
);

OAI32xp33_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_32),
.A3(n_35),
.B1(n_31),
.B2(n_21),
.Y(n_165)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_21),
.Y(n_166)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_41),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_168),
.C(n_170),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_132),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_41),
.C(n_37),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_131),
.A2(n_147),
.B(n_143),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_171),
.A2(n_184),
.B(n_185),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_132),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_175),
.A2(n_187),
.B(n_189),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_31),
.Y(n_178)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_R g179 ( 
.A1(n_136),
.A2(n_37),
.B1(n_31),
.B2(n_35),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_181),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_0),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_182),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_119),
.C(n_107),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_1),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_140),
.A2(n_16),
.B1(n_15),
.B2(n_13),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

AO21x2_ASAP7_75t_SL g189 ( 
.A1(n_149),
.A2(n_1),
.B(n_2),
.Y(n_189)
);

OAI22x1_ASAP7_75t_SL g190 ( 
.A1(n_189),
.A2(n_141),
.B1(n_129),
.B2(n_139),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_190),
.A2(n_206),
.B1(n_189),
.B2(n_161),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_191),
.A2(n_210),
.B1(n_185),
.B2(n_189),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_186),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_192),
.B(n_197),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_158),
.B(n_129),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_201),
.Y(n_226)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

OAI211xp5_ASAP7_75t_SL g197 ( 
.A1(n_183),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_198),
.A2(n_204),
.B1(n_211),
.B2(n_165),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_182),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_199),
.B(n_202),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_183),
.B(n_157),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_177),
.A2(n_130),
.B1(n_142),
.B2(n_155),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_161),
.A2(n_155),
.B1(n_16),
.B2(n_15),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_159),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_164),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g213 ( 
.A(n_167),
.B(n_13),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_166),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_214),
.A2(n_217),
.B(n_163),
.Y(n_243)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_189),
.Y(n_215)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_164),
.B(n_5),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_160),
.Y(n_219)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_202),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_228),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_168),
.C(n_181),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_227),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_180),
.C(n_170),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_198),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_171),
.Y(n_229)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_232),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_234),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_217),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_233),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_178),
.C(n_175),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_187),
.C(n_184),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_236),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_203),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_196),
.A2(n_176),
.B1(n_173),
.B2(n_169),
.Y(n_238)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_172),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_242),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_240),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_163),
.B1(n_188),
.B2(n_8),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_211),
.B1(n_190),
.B2(n_209),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_208),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_218),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_163),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_219),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_248),
.B(n_256),
.Y(n_279)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_252),
.A2(n_197),
.B(n_214),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_217),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_255),
.Y(n_283)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_266),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_205),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_264),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_205),
.Y(n_264)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_243),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_247),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_224),
.C(n_227),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_275),
.C(n_284),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_260),
.B(n_226),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_282),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_220),
.B1(n_230),
.B2(n_193),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_272),
.A2(n_277),
.B1(n_252),
.B2(n_254),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_265),
.A2(n_235),
.B1(n_234),
.B2(n_193),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_273),
.A2(n_276),
.B1(n_254),
.B2(n_258),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_239),
.C(n_236),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_257),
.A2(n_216),
.B1(n_225),
.B2(n_245),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_216),
.B1(n_218),
.B2(n_242),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_259),
.B(n_188),
.Y(n_278)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g281 ( 
.A(n_255),
.Y(n_281)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_246),
.B(n_226),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_286),
.A2(n_288),
.B1(n_276),
.B2(n_249),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_246),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_289),
.C(n_284),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_274),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_267),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_283),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_247),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g292 ( 
.A(n_277),
.B(n_250),
.CI(n_264),
.CON(n_292),
.SN(n_292)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_297),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_282),
.B1(n_270),
.B2(n_251),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_280),
.C(n_267),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_295),
.C(n_287),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_272),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_298),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_302),
.C(n_293),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_SL g301 ( 
.A(n_296),
.B(n_273),
.Y(n_301)
);

AO21x1_ASAP7_75t_SL g318 ( 
.A1(n_301),
.A2(n_306),
.B(n_308),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_280),
.C(n_262),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_303),
.A2(n_6),
.B(n_7),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_305),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_309),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_290),
.B(n_207),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_294),
.B(n_210),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_310),
.B(n_312),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_260),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_321),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_306),
.A2(n_292),
.B(n_285),
.Y(n_315)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_315),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_289),
.B(n_231),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_317),
.B(n_320),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_7),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_300),
.A2(n_10),
.B(n_12),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_12),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_6),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_324),
.B(n_325),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_6),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_316),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_328),
.A2(n_319),
.B(n_7),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_318),
.B1(n_8),
.B2(n_9),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_330),
.B(n_332),
.C(n_329),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_327),
.B(n_323),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

OAI211xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_326),
.B(n_319),
.C(n_331),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_9),
.C(n_313),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_9),
.Y(n_338)
);


endmodule