module fake_jpeg_2889_n_471 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_471);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_471;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_10),
.B(n_17),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_3),
.B(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_55),
.Y(n_135)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_57),
.B(n_60),
.Y(n_127)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_34),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_58),
.Y(n_173)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_19),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_61),
.B(n_62),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_14),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_63),
.B(n_64),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_29),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_29),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_65),
.B(n_71),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_31),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_66),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_67),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_68),
.Y(n_186)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_74),
.Y(n_194)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_76),
.Y(n_180)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_77),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_79),
.B(n_89),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_42),
.B(n_16),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_80),
.B(n_81),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_37),
.B(n_16),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_82),
.Y(n_184)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_20),
.B(n_16),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_90),
.Y(n_182)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_91),
.Y(n_190)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_92),
.Y(n_178)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_37),
.B(n_13),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_102),
.B(n_106),
.Y(n_169)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_103),
.B(n_116),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_39),
.B(n_13),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_39),
.B(n_1),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_108),
.B(n_109),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_21),
.B(n_1),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_110),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_27),
.Y(n_112)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_27),
.Y(n_114)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_31),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_24),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_77),
.B(n_35),
.C(n_25),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_132),
.B(n_168),
.C(n_150),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_55),
.A2(n_35),
.B1(n_25),
.B2(n_45),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_138),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_112),
.A2(n_40),
.B1(n_27),
.B2(n_45),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_89),
.A2(n_21),
.B1(n_46),
.B2(n_41),
.Y(n_136)
);

NAND2x1_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_30),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_137),
.A2(n_157),
.B(n_134),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_73),
.A2(n_49),
.B1(n_46),
.B2(n_41),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_49),
.B1(n_36),
.B2(n_44),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_142),
.A2(n_152),
.B1(n_157),
.B2(n_167),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_115),
.A2(n_95),
.B1(n_92),
.B2(n_76),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_151),
.A2(n_192),
.B1(n_121),
.B2(n_123),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_97),
.A2(n_36),
.B1(n_44),
.B2(n_28),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_99),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_66),
.B(n_30),
.Y(n_159)
);

NAND2x1_ASAP7_75t_SL g206 ( 
.A(n_159),
.B(n_101),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_58),
.B(n_2),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_164),
.B(n_185),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_67),
.A2(n_30),
.B1(n_38),
.B2(n_4),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_69),
.B(n_30),
.C(n_38),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_SL g174 ( 
.A1(n_68),
.A2(n_58),
.B(n_114),
.Y(n_174)
);

OR2x2_ASAP7_75t_SL g210 ( 
.A(n_174),
.B(n_156),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_113),
.B(n_2),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_176),
.B(n_195),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_70),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_179),
.A2(n_191),
.B1(n_175),
.B2(n_130),
.Y(n_230)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_83),
.Y(n_181)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_74),
.B(n_11),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_104),
.B(n_2),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_187),
.B(n_188),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_74),
.B(n_5),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_105),
.B(n_6),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_189),
.B(n_122),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_111),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_98),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_111),
.B(n_9),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_127),
.B(n_110),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_197),
.B(n_199),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_82),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_140),
.Y(n_200)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_200),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_159),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_201),
.B(n_208),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_146),
.B(n_84),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_202),
.B(n_209),
.Y(n_277)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_203),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_204),
.A2(n_207),
.B1(n_257),
.B2(n_259),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_170),
.A2(n_86),
.B1(n_94),
.B2(n_100),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_205),
.A2(n_244),
.B1(n_216),
.B2(n_227),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_206),
.B(n_210),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_139),
.A2(n_11),
.B1(n_193),
.B2(n_133),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_139),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_148),
.B(n_153),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_211),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_169),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_212),
.B(n_225),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_155),
.B(n_119),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_213),
.B(n_240),
.Y(n_297)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_214),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_215),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_216),
.B(n_219),
.Y(n_289)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_129),
.Y(n_217)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_217),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_147),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_218),
.B(n_222),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_144),
.B(n_137),
.C(n_190),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_220),
.B(n_240),
.C(n_251),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_150),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_223),
.Y(n_304)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_154),
.Y(n_224)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_224),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_131),
.B(n_141),
.Y(n_225)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_181),
.Y(n_229)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_229),
.Y(n_301)
);

OA22x2_ASAP7_75t_L g300 ( 
.A1(n_230),
.A2(n_260),
.B1(n_233),
.B2(n_248),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_182),
.B(n_173),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_232),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_135),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g295 ( 
.A(n_234),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_158),
.B(n_160),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_235),
.Y(n_294)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_236),
.B(n_237),
.Y(n_299)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_149),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_166),
.Y(n_238)
);

INVx11_ASAP7_75t_L g308 ( 
.A(n_238),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_135),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_239),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_186),
.B(n_122),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_118),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_241),
.A2(n_242),
.B1(n_246),
.B2(n_247),
.Y(n_268)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_126),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_245),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g244 ( 
.A1(n_142),
.A2(n_152),
.B1(n_138),
.B2(n_125),
.Y(n_244)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_178),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_248),
.A2(n_249),
.B1(n_253),
.B2(n_254),
.Y(n_306)
);

INVx4_ASAP7_75t_SL g249 ( 
.A(n_196),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_196),
.B(n_165),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_252),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_165),
.B(n_171),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_194),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_179),
.A2(n_196),
.B1(n_191),
.B2(n_184),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_120),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_120),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_256),
.Y(n_286)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_124),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_171),
.B(n_124),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_257),
.B(n_261),
.C(n_258),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_194),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_258),
.B(n_259),
.Y(n_303)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_125),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_128),
.Y(n_260)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_184),
.B(n_194),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g262 ( 
.A(n_219),
.B(n_128),
.CI(n_145),
.CON(n_262),
.SN(n_262)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_262),
.A2(n_278),
.B(n_270),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_204),
.A2(n_145),
.B1(n_210),
.B2(n_213),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_263),
.A2(n_269),
.B1(n_271),
.B2(n_274),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_228),
.A2(n_226),
.B1(n_244),
.B2(n_205),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_220),
.A2(n_198),
.B1(n_231),
.B2(n_251),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_276),
.A2(n_281),
.B1(n_296),
.B2(n_302),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_206),
.A2(n_242),
.B(n_229),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_251),
.A2(n_257),
.B1(n_254),
.B2(n_255),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_261),
.A2(n_256),
.B1(n_236),
.B2(n_234),
.Y(n_290)
);

AO21x2_ASAP7_75t_L g312 ( 
.A1(n_290),
.A2(n_293),
.B(n_286),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_214),
.A2(n_221),
.B1(n_237),
.B2(n_261),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_291),
.B(n_305),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_203),
.A2(n_211),
.B1(n_245),
.B2(n_260),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_221),
.A2(n_241),
.B1(n_215),
.B2(n_239),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_297),
.B(n_290),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_240),
.B(n_249),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_270),
.C(n_289),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_300),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_238),
.A2(n_226),
.B1(n_204),
.B2(n_205),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_262),
.B(n_266),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_309),
.B(n_314),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_310),
.A2(n_306),
.B(n_268),
.Y(n_357)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_312),
.Y(n_346)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_275),
.Y(n_313)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_313),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_266),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_269),
.A2(n_302),
.B1(n_289),
.B2(n_271),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_315),
.A2(n_279),
.B1(n_295),
.B2(n_308),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_293),
.Y(n_347)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_275),
.Y(n_318)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_318),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_264),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_322),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_284),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_320),
.Y(n_362)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_280),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_321),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_263),
.B(n_276),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_289),
.B(n_267),
.C(n_270),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_300),
.C(n_288),
.Y(n_351)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_286),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_324),
.B(n_325),
.Y(n_366)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_299),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_292),
.B(n_284),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_326),
.B(n_332),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_273),
.A2(n_285),
.B(n_267),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_327),
.A2(n_344),
.B(n_287),
.Y(n_359)
);

AND2x6_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_282),
.Y(n_328)
);

AOI31xp33_ASAP7_75t_SL g372 ( 
.A1(n_328),
.A2(n_327),
.A3(n_342),
.B(n_343),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_277),
.B(n_305),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_329),
.B(n_337),
.Y(n_355)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_299),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_330),
.B(n_334),
.Y(n_361)
);

INVx8_ASAP7_75t_L g331 ( 
.A(n_279),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_331),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_265),
.B(n_272),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_272),
.B(n_304),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_304),
.B(n_307),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_336),
.Y(n_350)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_299),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_303),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_339),
.Y(n_356)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_303),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_307),
.B(n_283),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_341),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_283),
.B(n_301),
.Y(n_341)
);

AO21x1_ASAP7_75t_L g342 ( 
.A1(n_278),
.A2(n_281),
.B(n_298),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_342),
.A2(n_317),
.B(n_335),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_343),
.B(n_323),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_301),
.B(n_280),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_345),
.B(n_347),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_352),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_300),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_357),
.A2(n_364),
.B(n_369),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_359),
.B(n_312),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_333),
.A2(n_322),
.B1(n_314),
.B2(n_309),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_363),
.A2(n_367),
.B1(n_312),
.B2(n_325),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_310),
.A2(n_300),
.B(n_287),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_365),
.A2(n_368),
.B1(n_312),
.B2(n_337),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_333),
.A2(n_295),
.B1(n_308),
.B2(n_312),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_315),
.A2(n_311),
.B1(n_335),
.B2(n_316),
.Y(n_368)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_372),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_342),
.A2(n_316),
.B(n_311),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_373),
.A2(n_312),
.B(n_329),
.Y(n_385)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_354),
.Y(n_374)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_374),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_371),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_376),
.B(n_377),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_324),
.Y(n_377)
);

OA21x2_ASAP7_75t_L g378 ( 
.A1(n_346),
.A2(n_339),
.B(n_338),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_378),
.A2(n_385),
.B(n_386),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_379),
.A2(n_396),
.B1(n_367),
.B2(n_378),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_358),
.B(n_362),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g401 ( 
.A(n_380),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_358),
.B(n_313),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_384),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_383),
.A2(n_365),
.B1(n_355),
.B2(n_357),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_330),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_361),
.B(n_328),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_SL g405 ( 
.A(n_387),
.B(n_382),
.C(n_353),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_360),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_389),
.A2(n_390),
.B(n_392),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_350),
.B(n_318),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_321),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_391),
.B(n_393),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_350),
.B(n_360),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_363),
.B(n_331),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_345),
.B(n_331),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_394),
.B(n_375),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_366),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_369),
.C(n_347),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_406),
.C(n_394),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_383),
.A2(n_368),
.B1(n_346),
.B2(n_373),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_400),
.A2(n_404),
.B1(n_407),
.B2(n_408),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_385),
.A2(n_352),
.B1(n_351),
.B2(n_364),
.Y(n_404)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_405),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_388),
.B(n_369),
.C(n_355),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_378),
.A2(n_349),
.B1(n_353),
.B2(n_372),
.Y(n_408)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_409),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_379),
.A2(n_349),
.B1(n_359),
.B2(n_361),
.Y(n_410)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_410),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_395),
.A2(n_348),
.B(n_370),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_411),
.A2(n_395),
.B(n_376),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_378),
.A2(n_370),
.B1(n_348),
.B2(n_354),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_390),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_415),
.B(n_384),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_417),
.B(n_428),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_401),
.B(n_389),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_418),
.B(n_420),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_401),
.B(n_387),
.Y(n_420)
);

XNOR2x1_ASAP7_75t_SL g423 ( 
.A(n_406),
.B(n_375),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_423),
.B(n_424),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_425),
.B(n_426),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_377),
.Y(n_426)
);

FAx1_ASAP7_75t_L g427 ( 
.A(n_397),
.B(n_393),
.CI(n_396),
.CON(n_427),
.SN(n_427)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_427),
.B(n_397),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_412),
.B(n_392),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_429),
.A2(n_403),
.B1(n_407),
.B2(n_402),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_424),
.B(n_398),
.C(n_404),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_430),
.B(n_438),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_408),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_433),
.B(n_440),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_434),
.B(n_417),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_422),
.B(n_380),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_436),
.B(n_381),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_416),
.A2(n_410),
.B1(n_409),
.B2(n_414),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_411),
.C(n_405),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_439),
.B(n_425),
.C(n_421),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_442),
.A2(n_446),
.B1(n_448),
.B2(n_433),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_443),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_444),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_421),
.C(n_416),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_435),
.A2(n_427),
.B(n_419),
.Y(n_447)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_447),
.Y(n_456)
);

NOR2xp67_ASAP7_75t_L g448 ( 
.A(n_432),
.B(n_402),
.Y(n_448)
);

AOI21xp33_ASAP7_75t_L g449 ( 
.A1(n_440),
.A2(n_412),
.B(n_427),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_449),
.A2(n_414),
.B1(n_419),
.B2(n_429),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_450),
.A2(n_447),
.B(n_441),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_442),
.A2(n_400),
.B1(n_439),
.B2(n_414),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_451),
.B(n_454),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_452),
.B(n_446),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_445),
.A2(n_413),
.B1(n_403),
.B2(n_437),
.Y(n_454)
);

NOR2xp67_ASAP7_75t_L g464 ( 
.A(n_457),
.B(n_454),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_455),
.B(n_444),
.C(n_441),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_458),
.A2(n_459),
.B(n_460),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_453),
.B(n_437),
.C(n_431),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_461),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_462),
.B(n_461),
.Y(n_465)
);

OAI21x1_ASAP7_75t_L g466 ( 
.A1(n_464),
.A2(n_451),
.B(n_456),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_465),
.B(n_466),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_467),
.B(n_463),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_468),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_469),
.B(n_431),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_470),
.A2(n_391),
.B(n_399),
.Y(n_471)
);


endmodule