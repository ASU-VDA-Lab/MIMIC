module fake_jpeg_26554_n_42 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_42);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_42;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_3),
.Y(n_24)
);

OAI32xp33_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_9),
.A3(n_17),
.B1(n_15),
.B2(n_4),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_19),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_30),
.B(n_0),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_36),
.B(n_37),
.Y(n_38)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_33),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_32),
.C(n_23),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_40),
.A2(n_21),
.B(n_1),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_5),
.C(n_18),
.Y(n_42)
);


endmodule