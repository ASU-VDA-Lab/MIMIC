module fake_jpeg_1587_n_151 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_151);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx6f_ASAP7_75t_SL g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_57),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_51),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_60),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_46),
.B(n_45),
.C(n_49),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_3),
.B(n_6),
.C(n_7),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_55),
.A2(n_53),
.B1(n_52),
.B2(n_40),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_67),
.B(n_2),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_2),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_53),
.B1(n_52),
.B2(n_40),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_42),
.B1(n_43),
.B2(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_77),
.Y(n_94)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_60),
.B1(n_42),
.B2(n_61),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_82),
.B1(n_62),
.B2(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_1),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_84),
.Y(n_93)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_60),
.B1(n_48),
.B2(n_4),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_85),
.Y(n_102)
);

AOI32xp33_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_48),
.A3(n_18),
.B1(n_20),
.B2(n_39),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_97),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_9),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_64),
.C(n_62),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_24),
.C(n_36),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_69),
.B(n_6),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_10),
.B(n_11),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_82),
.B1(n_85),
.B2(n_87),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_108),
.B1(n_114),
.B2(n_12),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_99),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_110),
.C(n_37),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_111),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_69),
.B1(n_84),
.B2(n_22),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_130)
);

AO22x1_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_90),
.B1(n_92),
.B2(n_101),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_25),
.B1(n_35),
.B2(n_34),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_16),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_10),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_117),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_11),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_123),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_118),
.A2(n_17),
.B(n_32),
.Y(n_122)
);

NOR3xp33_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_127),
.C(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_12),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_107),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_126),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_14),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_131),
.C(n_114),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_130),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_138),
.C(n_136),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_110),
.C(n_108),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g139 ( 
.A(n_136),
.B(n_121),
.CI(n_128),
.CON(n_139),
.SN(n_139)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_139),
.B(n_142),
.Y(n_143)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_141),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_141),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_147),
.A2(n_135),
.B(n_134),
.Y(n_148)
);

AOI322xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_122),
.A3(n_139),
.B1(n_143),
.B2(n_111),
.C1(n_126),
.C2(n_130),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_149),
.B(n_118),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_111),
.Y(n_151)
);


endmodule