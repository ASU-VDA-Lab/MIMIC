module fake_jpeg_5446_n_11 (n_3, n_2, n_1, n_0, n_4, n_5, n_11);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_11;

wire n_10;
wire n_8;
wire n_9;
wire n_6;
wire n_7;

NAND2xp5_ASAP7_75t_SL g6 ( 
.A(n_3),
.B(n_2),
.Y(n_6)
);

OA22x2_ASAP7_75t_L g7 ( 
.A1(n_0),
.A2(n_5),
.B1(n_4),
.B2(n_1),
.Y(n_7)
);

XNOR2xp5_ASAP7_75t_L g8 ( 
.A(n_7),
.B(n_0),
.Y(n_8)
);

OAI22xp5_ASAP7_75t_SL g9 ( 
.A1(n_8),
.A2(n_7),
.B1(n_6),
.B2(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_9),
.Y(n_10)
);

MAJx2_ASAP7_75t_L g11 ( 
.A(n_10),
.B(n_1),
.C(n_2),
.Y(n_11)
);


endmodule