module real_aes_1150_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g223 ( .A(n_0), .B(n_130), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_1), .B(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_2), .B(n_119), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_3), .B(n_128), .Y(n_459) );
INVx1_ASAP7_75t_L g118 ( .A(n_4), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_5), .B(n_119), .Y(n_176) );
NAND2xp33_ASAP7_75t_SL g169 ( .A(n_6), .B(n_125), .Y(n_169) );
INVx1_ASAP7_75t_L g149 ( .A(n_7), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g731 ( .A(n_8), .Y(n_731) );
AND2x2_ASAP7_75t_L g174 ( .A(n_9), .B(n_109), .Y(n_174) );
AND2x2_ASAP7_75t_L g452 ( .A(n_10), .B(n_166), .Y(n_452) );
AND2x2_ASAP7_75t_L g461 ( .A(n_11), .B(n_141), .Y(n_461) );
INVx2_ASAP7_75t_L g110 ( .A(n_12), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_13), .B(n_128), .Y(n_514) );
CKINVDCx16_ASAP7_75t_R g423 ( .A(n_14), .Y(n_423) );
AOI221x1_ASAP7_75t_L g163 ( .A1(n_15), .A2(n_113), .B1(n_164), .B2(n_166), .C(n_168), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_16), .B(n_119), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_17), .B(n_119), .Y(n_499) );
INVx1_ASAP7_75t_L g426 ( .A(n_18), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_19), .A2(n_87), .B1(n_119), .B2(n_151), .Y(n_440) );
AOI221xp5_ASAP7_75t_SL g112 ( .A1(n_20), .A2(n_34), .B1(n_113), .B2(n_119), .C(n_126), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_21), .A2(n_113), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_22), .B(n_130), .Y(n_179) );
OR2x2_ASAP7_75t_L g111 ( .A(n_23), .B(n_86), .Y(n_111) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_23), .A2(n_86), .B(n_110), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_24), .B(n_128), .Y(n_140) );
INVxp67_ASAP7_75t_L g162 ( .A(n_25), .Y(n_162) );
AND2x2_ASAP7_75t_L g212 ( .A(n_26), .B(n_108), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_27), .A2(n_113), .B(n_222), .Y(n_221) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_28), .A2(n_166), .B(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_29), .B(n_128), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_30), .A2(n_113), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_31), .B(n_128), .Y(n_494) );
AND2x2_ASAP7_75t_L g114 ( .A(n_32), .B(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g125 ( .A(n_32), .B(n_118), .Y(n_125) );
INVx1_ASAP7_75t_L g158 ( .A(n_32), .Y(n_158) );
OR2x6_ASAP7_75t_L g424 ( .A(n_33), .B(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_35), .B(n_119), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_36), .A2(n_79), .B1(n_113), .B2(n_156), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_37), .B(n_128), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_38), .B(n_119), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_39), .B(n_130), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_40), .A2(n_113), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g226 ( .A(n_41), .B(n_108), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_42), .B(n_130), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_43), .B(n_108), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_44), .B(n_119), .Y(n_511) );
INVx1_ASAP7_75t_L g117 ( .A(n_45), .Y(n_117) );
INVx1_ASAP7_75t_L g122 ( .A(n_45), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_46), .B(n_128), .Y(n_450) );
AND2x2_ASAP7_75t_L g480 ( .A(n_47), .B(n_108), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_48), .B(n_119), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_49), .B(n_130), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_50), .B(n_130), .Y(n_493) );
AND2x2_ASAP7_75t_L g190 ( .A(n_51), .B(n_108), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_52), .B(n_119), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_53), .B(n_128), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_54), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_55), .B(n_119), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_56), .A2(n_113), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_SL g143 ( .A(n_57), .B(n_109), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_58), .B(n_130), .Y(n_187) );
AND2x2_ASAP7_75t_L g505 ( .A(n_59), .B(n_109), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_60), .A2(n_113), .B(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_61), .B(n_128), .Y(n_180) );
AND2x2_ASAP7_75t_SL g197 ( .A(n_62), .B(n_141), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_63), .B(n_130), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_64), .B(n_130), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_65), .A2(n_89), .B1(n_113), .B2(n_156), .Y(n_441) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_66), .A2(n_99), .B1(n_724), .B2(n_735), .C1(n_751), .C2(n_753), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_66), .A2(n_738), .B1(n_739), .B2(n_741), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_66), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_67), .B(n_128), .Y(n_502) );
OAI222xp33_ASAP7_75t_L g99 ( .A1(n_68), .A2(n_100), .B1(n_715), .B2(n_716), .C1(n_720), .C2(n_723), .Y(n_99) );
INVx1_ASAP7_75t_L g715 ( .A(n_68), .Y(n_715) );
INVx1_ASAP7_75t_L g115 ( .A(n_69), .Y(n_115) );
INVx1_ASAP7_75t_L g124 ( .A(n_69), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_70), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_71), .B(n_130), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_72), .A2(n_113), .B(n_484), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_73), .A2(n_113), .B(n_470), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_74), .A2(n_113), .B(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g496 ( .A(n_75), .B(n_109), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_76), .B(n_108), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_77), .B(n_119), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_78), .A2(n_81), .B1(n_119), .B2(n_151), .Y(n_195) );
INVx1_ASAP7_75t_L g427 ( .A(n_80), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_82), .B(n_130), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_83), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g473 ( .A(n_84), .B(n_141), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_85), .A2(n_113), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_88), .B(n_128), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_90), .A2(n_113), .B(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_91), .B(n_128), .Y(n_471) );
INVxp67_ASAP7_75t_L g165 ( .A(n_92), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_93), .B(n_119), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_94), .B(n_128), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_95), .A2(n_113), .B(n_138), .Y(n_137) );
BUFx2_ASAP7_75t_L g504 ( .A(n_96), .Y(n_504) );
BUFx2_ASAP7_75t_L g732 ( .A(n_97), .Y(n_732) );
BUFx2_ASAP7_75t_SL g757 ( .A(n_97), .Y(n_757) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OAI22xp5_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_419), .B1(n_428), .B2(n_711), .Y(n_101) );
INVx2_ASAP7_75t_L g717 ( .A(n_102), .Y(n_717) );
INVx4_ASAP7_75t_L g740 ( .A(n_102), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_102), .Y(n_741) );
OR2x6_ASAP7_75t_L g102 ( .A(n_103), .B(n_332), .Y(n_102) );
NAND3xp33_ASAP7_75t_SL g103 ( .A(n_104), .B(n_242), .C(n_282), .Y(n_103) );
O2A1O1Ixp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_144), .B(n_171), .C(n_198), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_105), .B(n_247), .Y(n_281) );
NOR2x1p5_ASAP7_75t_L g105 ( .A(n_106), .B(n_133), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g217 ( .A(n_107), .Y(n_217) );
INVx2_ASAP7_75t_L g233 ( .A(n_107), .Y(n_233) );
OR2x2_ASAP7_75t_L g245 ( .A(n_107), .B(n_134), .Y(n_245) );
AND2x2_ASAP7_75t_L g259 ( .A(n_107), .B(n_218), .Y(n_259) );
INVx1_ASAP7_75t_L g287 ( .A(n_107), .Y(n_287) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_107), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_107), .B(n_134), .Y(n_393) );
OA21x2_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_112), .B(n_132), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_108), .Y(n_189) );
AO21x2_ASAP7_75t_L g439 ( .A1(n_108), .A2(n_440), .B(n_441), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_108), .A2(n_468), .B(n_469), .Y(n_467) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AND2x4_ASAP7_75t_L g150 ( .A(n_110), .B(n_111), .Y(n_150) );
AND2x6_ASAP7_75t_L g113 ( .A(n_114), .B(n_116), .Y(n_113) );
BUFx3_ASAP7_75t_L g155 ( .A(n_114), .Y(n_155) );
AND2x6_ASAP7_75t_L g130 ( .A(n_115), .B(n_121), .Y(n_130) );
INVx2_ASAP7_75t_L g160 ( .A(n_115), .Y(n_160) );
AND2x4_ASAP7_75t_L g156 ( .A(n_116), .B(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
AND2x4_ASAP7_75t_L g128 ( .A(n_117), .B(n_123), .Y(n_128) );
INVx2_ASAP7_75t_L g153 ( .A(n_117), .Y(n_153) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_118), .Y(n_154) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_125), .Y(n_119) );
INVx1_ASAP7_75t_L g170 ( .A(n_120), .Y(n_170) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_123), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx5_ASAP7_75t_L g131 ( .A(n_125), .Y(n_131) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_129), .B(n_131), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_130), .B(n_504), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_131), .A2(n_139), .B(n_140), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_131), .A2(n_179), .B(n_180), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_131), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_131), .A2(n_209), .B(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_131), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_131), .A2(n_449), .B(n_450), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_131), .A2(n_458), .B(n_459), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_131), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_131), .A2(n_485), .B(n_486), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_131), .A2(n_493), .B(n_494), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_131), .A2(n_502), .B(n_503), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_131), .A2(n_514), .B(n_515), .Y(n_513) );
OR2x2_ASAP7_75t_L g214 ( .A(n_133), .B(n_215), .Y(n_214) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_133), .Y(n_349) );
AND2x2_ASAP7_75t_L g354 ( .A(n_133), .B(n_216), .Y(n_354) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g144 ( .A(n_134), .B(n_145), .Y(n_144) );
OR2x2_ASAP7_75t_L g213 ( .A(n_134), .B(n_146), .Y(n_213) );
OR2x2_ASAP7_75t_L g232 ( .A(n_134), .B(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g261 ( .A(n_134), .Y(n_261) );
AND2x4_ASAP7_75t_SL g300 ( .A(n_134), .B(n_146), .Y(n_300) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_134), .Y(n_304) );
OR2x2_ASAP7_75t_L g321 ( .A(n_134), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g331 ( .A(n_134), .B(n_238), .Y(n_331) );
INVx1_ASAP7_75t_L g360 ( .A(n_134), .Y(n_360) );
OR2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_143), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_137), .B(n_141), .Y(n_135) );
INVx2_ASAP7_75t_SL g193 ( .A(n_141), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_141), .A2(n_499), .B(n_500), .Y(n_498) );
BUFx4f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx3_ASAP7_75t_L g167 ( .A(n_142), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_144), .B(n_289), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_145), .B(n_218), .Y(n_235) );
AND2x2_ASAP7_75t_L g247 ( .A(n_145), .B(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g265 ( .A(n_145), .B(n_232), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_145), .B(n_286), .Y(n_285) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g238 ( .A(n_146), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g260 ( .A(n_146), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g295 ( .A(n_146), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_146), .B(n_218), .Y(n_319) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_163), .Y(n_146) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_151), .B1(n_156), .B2(n_161), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_150), .B(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_150), .B(n_165), .Y(n_164) );
NOR3xp33_ASAP7_75t_L g168 ( .A(n_150), .B(n_169), .C(n_170), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_150), .A2(n_176), .B(n_177), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_150), .A2(n_482), .B(n_483), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_150), .A2(n_511), .B(n_512), .Y(n_510) );
AND2x4_ASAP7_75t_L g151 ( .A(n_152), .B(n_155), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
NOR2x1p5_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g489 ( .A(n_166), .Y(n_489) );
INVx4_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI21x1_ASAP7_75t_L g219 ( .A1(n_167), .A2(n_220), .B(n_226), .Y(n_219) );
AO21x2_ASAP7_75t_L g445 ( .A1(n_167), .A2(n_446), .B(n_452), .Y(n_445) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_181), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_172), .B(n_251), .Y(n_250) );
AND2x4_ASAP7_75t_L g268 ( .A(n_172), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_172), .B(n_182), .Y(n_273) );
NAND3xp33_ASAP7_75t_L g288 ( .A(n_172), .B(n_289), .C(n_290), .Y(n_288) );
AND2x2_ASAP7_75t_L g336 ( .A(n_172), .B(n_241), .Y(n_336) );
INVx5_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g203 ( .A(n_173), .B(n_204), .Y(n_203) );
AND2x4_ASAP7_75t_SL g240 ( .A(n_173), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g256 ( .A(n_173), .Y(n_256) );
OR2x2_ASAP7_75t_L g279 ( .A(n_173), .B(n_269), .Y(n_279) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_173), .Y(n_296) );
AND2x2_ASAP7_75t_SL g314 ( .A(n_173), .B(n_202), .Y(n_314) );
AND2x4_ASAP7_75t_L g329 ( .A(n_173), .B(n_205), .Y(n_329) );
AND2x2_ASAP7_75t_L g343 ( .A(n_173), .B(n_182), .Y(n_343) );
OR2x2_ASAP7_75t_L g364 ( .A(n_173), .B(n_191), .Y(n_364) );
OR2x6_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
AND2x2_ASAP7_75t_L g418 ( .A(n_181), .B(n_296), .Y(n_418) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_191), .Y(n_181) );
AND2x4_ASAP7_75t_L g241 ( .A(n_182), .B(n_204), .Y(n_241) );
INVx2_ASAP7_75t_L g252 ( .A(n_182), .Y(n_252) );
AND2x2_ASAP7_75t_L g257 ( .A(n_182), .B(n_202), .Y(n_257) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_182), .Y(n_290) );
OR2x2_ASAP7_75t_L g313 ( .A(n_182), .B(n_205), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_182), .B(n_205), .Y(n_316) );
INVx1_ASAP7_75t_L g325 ( .A(n_182), .Y(n_325) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_189), .B(n_190), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_188), .Y(n_183) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_189), .A2(n_206), .B(n_212), .Y(n_205) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_189), .A2(n_206), .B(n_212), .Y(n_269) );
AOI21x1_ASAP7_75t_L g454 ( .A1(n_189), .A2(n_455), .B(n_461), .Y(n_454) );
AND2x2_ASAP7_75t_L g228 ( .A(n_191), .B(n_205), .Y(n_228) );
BUFx2_ASAP7_75t_L g277 ( .A(n_191), .Y(n_277) );
AND2x2_ASAP7_75t_L g372 ( .A(n_191), .B(n_252), .Y(n_372) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_192), .Y(n_202) );
AOI21x1_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_197), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
OAI221xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_213), .B1(n_214), .B2(n_227), .C(n_229), .Y(n_198) );
INVx1_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_203), .Y(n_200) );
NOR2x1_ASAP7_75t_L g274 ( .A(n_201), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_201), .B(n_268), .Y(n_308) );
OR2x2_ASAP7_75t_L g320 ( .A(n_201), .B(n_316), .Y(n_320) );
OR2x2_ASAP7_75t_L g323 ( .A(n_201), .B(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g412 ( .A(n_201), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x4_ASAP7_75t_L g251 ( .A(n_202), .B(n_252), .Y(n_251) );
OA33x2_ASAP7_75t_L g284 ( .A1(n_202), .A2(n_245), .A3(n_285), .B1(n_288), .B2(n_291), .B3(n_294), .Y(n_284) );
OR2x2_ASAP7_75t_L g315 ( .A(n_202), .B(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g339 ( .A(n_202), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g347 ( .A(n_202), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g367 ( .A(n_202), .B(n_241), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_202), .B(n_256), .Y(n_405) );
INVx2_ASAP7_75t_L g275 ( .A(n_203), .Y(n_275) );
AOI322xp5_ASAP7_75t_L g345 ( .A1(n_203), .A2(n_258), .A3(n_346), .B1(n_349), .B2(n_350), .C1(n_352), .C2(n_354), .Y(n_345) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_205), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_211), .Y(n_206) );
OR2x2_ASAP7_75t_L g327 ( .A(n_213), .B(n_306), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_213), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_SL g400 ( .A(n_213), .Y(n_400) );
INVx1_ASAP7_75t_SL g266 ( .A(n_214), .Y(n_266) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g299 ( .A(n_216), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g239 ( .A(n_218), .Y(n_239) );
INVx1_ASAP7_75t_L g248 ( .A(n_218), .Y(n_248) );
INVx1_ASAP7_75t_L g289 ( .A(n_218), .Y(n_289) );
OR2x2_ASAP7_75t_L g306 ( .A(n_218), .B(n_233), .Y(n_306) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_218), .Y(n_381) );
INVx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_225), .Y(n_220) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_SL g350 ( .A(n_228), .B(n_351), .Y(n_350) );
OAI21xp5_ASAP7_75t_SL g229 ( .A1(n_230), .A2(n_236), .B(n_240), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g303 ( .A1(n_230), .A2(n_304), .B(n_305), .C(n_307), .Y(n_303) );
AND2x4_ASAP7_75t_L g230 ( .A(n_231), .B(n_234), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g368 ( .A(n_232), .B(n_369), .Y(n_368) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_233), .Y(n_237) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
OR2x2_ASAP7_75t_L g392 ( .A(n_235), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
AND2x2_ASAP7_75t_SL g361 ( .A(n_238), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g369 ( .A(n_238), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_238), .B(n_360), .Y(n_377) );
INVx3_ASAP7_75t_SL g302 ( .A(n_241), .Y(n_302) );
AOI221xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_249), .B1(n_253), .B2(n_258), .C(n_262), .Y(n_242) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_248), .Y(n_293) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_251), .A2(n_278), .B(n_350), .Y(n_356) );
AND2x2_ASAP7_75t_L g382 ( .A(n_251), .B(n_329), .Y(n_382) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_252), .Y(n_270) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_256), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g391 ( .A(n_256), .B(n_313), .Y(n_391) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx2_ASAP7_75t_L g340 ( .A(n_259), .Y(n_340) );
OAI21xp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_267), .B(n_271), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
INVx2_ASAP7_75t_L g413 ( .A(n_268), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_269), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g342 ( .A(n_269), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_270), .B(n_292), .Y(n_291) );
OAI31xp33_ASAP7_75t_SL g271 ( .A1(n_272), .A2(n_274), .A3(n_276), .B(n_280), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_275), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
OR2x2_ASAP7_75t_L g353 ( .A(n_277), .B(n_279), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_277), .B(n_329), .Y(n_408) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NOR5xp2_ASAP7_75t_L g282 ( .A(n_283), .B(n_297), .C(n_309), .D(n_318), .E(n_326), .Y(n_282) );
INVxp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_287), .B(n_289), .Y(n_322) );
INVx1_ASAP7_75t_L g362 ( .A(n_287), .Y(n_362) );
INVxp67_ASAP7_75t_SL g399 ( .A(n_287), .Y(n_399) );
INVx1_ASAP7_75t_L g351 ( .A(n_290), .Y(n_351) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp33_ASAP7_75t_SL g294 ( .A(n_295), .B(n_296), .Y(n_294) );
OAI321xp33_ASAP7_75t_L g334 ( .A1(n_295), .A2(n_335), .A3(n_337), .B1(n_341), .B2(n_344), .C(n_345), .Y(n_334) );
INVx1_ASAP7_75t_L g388 ( .A(n_296), .Y(n_388) );
OAI21xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_301), .B(n_303), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_299), .A2(n_372), .B1(n_379), .B2(n_382), .Y(n_378) );
AND2x2_ASAP7_75t_L g407 ( .A(n_300), .B(n_381), .Y(n_407) );
INVx1_ASAP7_75t_L g317 ( .A(n_305), .Y(n_317) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_315), .B(n_317), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_316), .A2(n_327), .B1(n_328), .B2(n_330), .Y(n_326) );
INVx1_ASAP7_75t_L g389 ( .A(n_316), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_320), .B1(n_321), .B2(n_323), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_325), .B(n_329), .Y(n_328) );
OAI221xp5_ASAP7_75t_L g403 ( .A1(n_327), .A2(n_404), .B1(n_406), .B2(n_408), .C(n_409), .Y(n_403) );
INVx1_ASAP7_75t_L g410 ( .A(n_327), .Y(n_410) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_328), .A2(n_385), .B1(n_392), .B2(n_394), .C(n_395), .Y(n_384) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_330), .A2(n_356), .B(n_357), .Y(n_355) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_383), .Y(n_332) );
NOR3xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_355), .C(n_373), .Y(n_333) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_336), .Y(n_402) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g401 ( .A(n_344), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_346), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g394 ( .A(n_354), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_363), .B(n_365), .Y(n_357) );
INVxp67_ASAP7_75t_L g415 ( .A(n_358), .Y(n_415) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_SL g370 ( .A(n_361), .Y(n_370) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
OAI22xp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_368), .B1(n_370), .B2(n_371), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI21xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B(n_378), .Y(n_373) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g416 ( .A(n_379), .Y(n_416) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NOR3xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_403), .C(n_414), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_390), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI21xp5_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_401), .B(n_402), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_400), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g409 ( .A1(n_407), .A2(n_410), .B(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AOI21xp33_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B(n_417), .Y(n_414) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx4_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
CKINVDCx6p67_ASAP7_75t_R g718 ( .A(n_420), .Y(n_718) );
INVx3_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_422), .Y(n_421) );
AND2x6_ASAP7_75t_SL g422 ( .A(n_423), .B(n_424), .Y(n_422) );
OR2x6_ASAP7_75t_SL g713 ( .A(n_423), .B(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g722 ( .A(n_423), .B(n_424), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_423), .B(n_714), .Y(n_734) );
CKINVDCx5p33_ASAP7_75t_R g714 ( .A(n_424), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx4_ASAP7_75t_L g719 ( .A(n_428), .Y(n_719) );
OR2x6_ASAP7_75t_L g428 ( .A(n_429), .B(n_648), .Y(n_428) );
NAND3xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_564), .C(n_601), .Y(n_429) );
NOR3xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_532), .C(n_547), .Y(n_430) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_477), .B1(n_506), .B2(n_518), .C(n_519), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_434), .B(n_462), .Y(n_433) );
OAI22xp33_ASAP7_75t_SL g592 ( .A1(n_434), .A2(n_556), .B1(n_593), .B2(n_596), .Y(n_592) );
OR2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_442), .Y(n_434) );
OAI21xp33_ASAP7_75t_SL g602 ( .A1(n_435), .A2(n_603), .B(n_609), .Y(n_602) );
OR2x2_ASAP7_75t_L g631 ( .A(n_435), .B(n_464), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_435), .B(n_551), .Y(n_632) );
INVx2_ASAP7_75t_L g663 ( .A(n_435), .Y(n_663) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_436), .B(n_523), .Y(n_644) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g518 ( .A(n_437), .B(n_445), .Y(n_518) );
BUFx3_ASAP7_75t_L g544 ( .A(n_437), .Y(n_544) );
AND2x2_ASAP7_75t_L g680 ( .A(n_437), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g703 ( .A(n_437), .B(n_465), .Y(n_703) );
AND2x4_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
AND2x4_ASAP7_75t_L g476 ( .A(n_438), .B(n_439), .Y(n_476) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_443), .B(n_465), .Y(n_623) );
INVx1_ASAP7_75t_L g660 ( .A(n_443), .Y(n_660) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_453), .Y(n_443) );
AND2x2_ASAP7_75t_L g475 ( .A(n_444), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g681 ( .A(n_444), .Y(n_681) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g524 ( .A(n_445), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_445), .B(n_453), .Y(n_525) );
AND2x2_ASAP7_75t_L g546 ( .A(n_445), .B(n_466), .Y(n_546) );
AND2x2_ASAP7_75t_L g628 ( .A(n_445), .B(n_454), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_451), .Y(n_446) );
AND2x4_ASAP7_75t_SL g521 ( .A(n_453), .B(n_466), .Y(n_521) );
INVx1_ASAP7_75t_L g552 ( .A(n_453), .Y(n_552) );
INVx2_ASAP7_75t_L g560 ( .A(n_453), .Y(n_560) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_453), .Y(n_584) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_454), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_460), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_475), .Y(n_462) );
AND2x2_ASAP7_75t_L g699 ( .A(n_463), .B(n_562), .Y(n_699) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_474), .Y(n_464) );
NAND2x1p5_ASAP7_75t_L g558 ( .A(n_465), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g610 ( .A(n_465), .B(n_525), .Y(n_610) );
AND2x2_ASAP7_75t_L g627 ( .A(n_465), .B(n_628), .Y(n_627) );
INVx4_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_L g551 ( .A(n_466), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g567 ( .A(n_466), .Y(n_567) );
AND2x2_ASAP7_75t_L g611 ( .A(n_466), .B(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g618 ( .A(n_466), .B(n_619), .Y(n_618) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_466), .B(n_524), .Y(n_633) );
BUFx2_ASAP7_75t_L g643 ( .A(n_466), .Y(n_643) );
AND2x2_ASAP7_75t_L g668 ( .A(n_466), .B(n_628), .Y(n_668) );
AND2x2_ASAP7_75t_L g689 ( .A(n_466), .B(n_690), .Y(n_689) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_473), .Y(n_466) );
INVx1_ASAP7_75t_L g620 ( .A(n_474), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_475), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g650 ( .A(n_475), .B(n_521), .Y(n_650) );
INVx3_ASAP7_75t_L g557 ( .A(n_476), .Y(n_557) );
AND2x2_ASAP7_75t_L g690 ( .A(n_476), .B(n_612), .Y(n_690) );
INVx1_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_478), .A2(n_520), .B1(n_525), .B2(n_526), .Y(n_519) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_487), .Y(n_478) );
INVx4_ASAP7_75t_L g517 ( .A(n_479), .Y(n_517) );
INVx2_ASAP7_75t_L g554 ( .A(n_479), .Y(n_554) );
NAND2x1_ASAP7_75t_L g580 ( .A(n_479), .B(n_497), .Y(n_580) );
OR2x2_ASAP7_75t_L g595 ( .A(n_479), .B(n_530), .Y(n_595) );
OR2x2_ASAP7_75t_SL g622 ( .A(n_479), .B(n_594), .Y(n_622) );
AND2x2_ASAP7_75t_L g635 ( .A(n_479), .B(n_509), .Y(n_635) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_479), .Y(n_656) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx2_ASAP7_75t_L g535 ( .A(n_487), .Y(n_535) );
AND2x2_ASAP7_75t_L g667 ( .A(n_487), .B(n_641), .Y(n_667) );
NOR2x1_ASAP7_75t_SL g487 ( .A(n_488), .B(n_497), .Y(n_487) );
AND2x2_ASAP7_75t_L g508 ( .A(n_488), .B(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g684 ( .A(n_488), .B(n_607), .Y(n_684) );
AO21x1_ASAP7_75t_SL g488 ( .A1(n_489), .A2(n_490), .B(n_496), .Y(n_488) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_489), .A2(n_490), .B(n_496), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_495), .Y(n_490) );
OR2x2_ASAP7_75t_L g516 ( .A(n_497), .B(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g527 ( .A(n_497), .B(n_517), .Y(n_527) );
AND2x2_ASAP7_75t_L g573 ( .A(n_497), .B(n_530), .Y(n_573) );
OR2x2_ASAP7_75t_L g594 ( .A(n_497), .B(n_509), .Y(n_594) );
INVx2_ASAP7_75t_SL g600 ( .A(n_497), .Y(n_600) );
AND2x2_ASAP7_75t_L g606 ( .A(n_497), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g616 ( .A(n_497), .B(n_599), .Y(n_616) );
BUFx2_ASAP7_75t_L g638 ( .A(n_497), .Y(n_638) );
OR2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_505), .Y(n_497) );
INVx2_ASAP7_75t_L g685 ( .A(n_506), .Y(n_685) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_516), .Y(n_506) );
OR2x2_ASAP7_75t_L g710 ( .A(n_507), .B(n_554), .Y(n_710) );
INVx2_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_508), .B(n_517), .Y(n_576) );
AND2x2_ASAP7_75t_L g647 ( .A(n_508), .B(n_527), .Y(n_647) );
INVx1_ASAP7_75t_L g529 ( .A(n_509), .Y(n_529) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_509), .Y(n_538) );
INVx1_ASAP7_75t_L g571 ( .A(n_509), .Y(n_571) );
INVx2_ASAP7_75t_L g607 ( .A(n_509), .Y(n_607) );
NOR2xp67_ASAP7_75t_L g537 ( .A(n_517), .B(n_538), .Y(n_537) );
BUFx2_ASAP7_75t_L g597 ( .A(n_517), .Y(n_597) );
INVx2_ASAP7_75t_SL g673 ( .A(n_518), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_520), .A2(n_575), .B1(n_577), .B2(n_581), .Y(n_574) );
AND2x2_ASAP7_75t_SL g520 ( .A(n_521), .B(n_522), .Y(n_520) );
AND2x2_ASAP7_75t_L g701 ( .A(n_521), .B(n_557), .Y(n_701) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_523), .B(n_567), .Y(n_646) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g612 ( .A(n_524), .B(n_560), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_525), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g555 ( .A(n_526), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_526), .A2(n_670), .B1(n_674), .B2(n_676), .C(n_678), .Y(n_669) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
AND2x2_ASAP7_75t_L g539 ( .A(n_527), .B(n_540), .Y(n_539) );
INVxp67_ASAP7_75t_SL g563 ( .A(n_527), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_527), .B(n_570), .Y(n_625) );
INVx1_ASAP7_75t_SL g621 ( .A(n_528), .Y(n_621) );
AOI221xp5_ASAP7_75t_SL g649 ( .A1(n_528), .A2(n_539), .B1(n_650), .B2(n_651), .C(n_654), .Y(n_649) );
AOI322xp5_ASAP7_75t_L g682 ( .A1(n_528), .A2(n_600), .A3(n_627), .B1(n_683), .B2(n_685), .C1(n_686), .C2(n_689), .Y(n_682) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
BUFx2_ASAP7_75t_L g549 ( .A(n_529), .Y(n_549) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_530), .Y(n_541) );
INVx2_ASAP7_75t_L g599 ( .A(n_530), .Y(n_599) );
AND2x2_ASAP7_75t_L g640 ( .A(n_530), .B(n_641), .Y(n_640) );
INVx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OA21x2_ASAP7_75t_SL g532 ( .A1(n_533), .A2(n_539), .B(n_542), .Y(n_532) );
AOI211xp5_ASAP7_75t_L g702 ( .A1(n_533), .A2(n_703), .B(n_704), .C(n_708), .Y(n_702) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
OR2x2_ASAP7_75t_L g591 ( .A(n_535), .B(n_553), .Y(n_591) );
OR2x2_ASAP7_75t_L g675 ( .A(n_535), .B(n_570), .Y(n_675) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g615 ( .A(n_537), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g693 ( .A(n_540), .Y(n_693) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g579 ( .A(n_541), .Y(n_579) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
OR2x2_ASAP7_75t_L g548 ( .A(n_544), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g583 ( .A(n_546), .B(n_584), .Y(n_583) );
OAI322xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_550), .A3(n_553), .B1(n_555), .B2(n_556), .C1(n_561), .C2(n_563), .Y(n_547) );
INVx1_ASAP7_75t_L g589 ( .A(n_548), .Y(n_589) );
OR2x2_ASAP7_75t_L g561 ( .A(n_550), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_550), .B(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g572 ( .A(n_554), .B(n_573), .Y(n_572) );
OAI32xp33_ASAP7_75t_L g617 ( .A1(n_554), .A2(n_618), .A3(n_621), .B1(n_622), .B2(n_623), .Y(n_617) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx2_ASAP7_75t_L g562 ( .A(n_557), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_557), .B(n_620), .Y(n_619) );
NOR2x1_ASAP7_75t_L g659 ( .A(n_557), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g683 ( .A(n_557), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g604 ( .A(n_558), .Y(n_604) );
INVx1_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_562), .B(n_628), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_585), .Y(n_564) );
OAI21xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_568), .B(n_574), .Y(n_565) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x4_ASAP7_75t_SL g569 ( .A(n_570), .B(n_572), .Y(n_569) );
INVx3_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g634 ( .A(n_573), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_576), .A2(n_596), .B1(n_698), .B2(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g624 ( .A1(n_578), .A2(n_625), .B(n_626), .C(n_629), .Y(n_624) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx3_ASAP7_75t_L g706 ( .A(n_580), .Y(n_706) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g587 ( .A(n_584), .Y(n_587) );
AO21x1_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_588), .B(n_592), .Y(n_585) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g652 ( .A(n_587), .Y(n_652) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_593), .B(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx1_ASAP7_75t_L g608 ( .A(n_595), .Y(n_608) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g665 ( .A(n_598), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NOR3xp33_ASAP7_75t_L g601 ( .A(n_602), .B(n_624), .C(n_636), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
OAI21xp5_ASAP7_75t_SL g666 ( .A1(n_605), .A2(n_667), .B(n_668), .Y(n_666) );
AND2x4_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVx1_ASAP7_75t_L g641 ( .A(n_607), .Y(n_641) );
O2A1O1Ixp5_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_611), .B(n_613), .C(n_617), .Y(n_609) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_619), .Y(n_709) );
INVx2_ASAP7_75t_L g694 ( .A(n_622), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g708 ( .A1(n_623), .A2(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g688 ( .A(n_628), .Y(n_688) );
OAI31xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .A3(n_633), .B(n_634), .Y(n_629) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g707 ( .A(n_635), .Y(n_707) );
OAI21xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_642), .B(n_645), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
BUFx2_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g657 ( .A(n_640), .Y(n_657) );
AOI21xp33_ASAP7_75t_SL g704 ( .A1(n_642), .A2(n_705), .B(n_707), .Y(n_704) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx2_ASAP7_75t_L g672 ( .A(n_643), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_643), .B(n_663), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_643), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g653 ( .A(n_644), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
NAND5xp2_ASAP7_75t_L g648 ( .A(n_649), .B(n_669), .C(n_682), .D(n_691), .E(n_702), .Y(n_648) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_658), .B1(n_661), .B2(n_664), .C(n_666), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVxp67_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_695), .B(n_697), .Y(n_691) );
AND2x4_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OA22x2_ASAP7_75t_L g716 ( .A1(n_711), .A2(n_717), .B1(n_718), .B2(n_719), .Y(n_716) );
CKINVDCx5p33_ASAP7_75t_R g711 ( .A(n_712), .Y(n_711) );
CKINVDCx11_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx3_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_733), .Y(n_726) );
INVxp67_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g728 ( .A(n_729), .B(n_732), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_SL g752 ( .A(n_730), .B(n_732), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_730), .A2(n_755), .B(n_758), .Y(n_754) );
BUFx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx2_ASAP7_75t_R g744 ( .A(n_734), .Y(n_744) );
BUFx3_ASAP7_75t_L g749 ( .A(n_734), .Y(n_749) );
BUFx2_ASAP7_75t_L g759 ( .A(n_734), .Y(n_759) );
INVxp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_742), .B(n_745), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
NOR2xp33_ASAP7_75t_SL g745 ( .A(n_746), .B(n_750), .Y(n_745) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
BUFx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
CKINVDCx11_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
CKINVDCx8_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
endmodule