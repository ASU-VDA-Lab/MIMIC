module fake_jpeg_3655_n_322 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx8_ASAP7_75t_SL g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_47),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_46),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_23),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_54),
.Y(n_104)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_52),
.Y(n_93)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_1),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_26),
.B(n_3),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_59),
.B(n_4),
.Y(n_115)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_63),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_71),
.Y(n_107)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

BUFx6f_ASAP7_75t_SL g68 ( 
.A(n_43),
.Y(n_68)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_22),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_73),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_22),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_82),
.Y(n_121)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx5_ASAP7_75t_SL g116 ( 
.A(n_77),
.Y(n_116)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_27),
.B(n_3),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_84),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_24),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_37),
.B(n_3),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_5),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_18),
.B1(n_32),
.B2(n_34),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_87),
.A2(n_91),
.B1(n_97),
.B2(n_101),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_59),
.A2(n_39),
.B1(n_34),
.B2(n_24),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_21),
.B1(n_39),
.B2(n_34),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_130),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_49),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_27),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_98),
.B(n_133),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_45),
.A2(n_29),
.B1(n_41),
.B2(n_30),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_46),
.A2(n_42),
.B1(n_41),
.B2(n_30),
.Y(n_106)
);

BUFx24_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_55),
.A2(n_42),
.B1(n_36),
.B2(n_31),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_SL g170 ( 
.A(n_112),
.B(n_77),
.C(n_81),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_58),
.A2(n_36),
.B1(n_31),
.B2(n_29),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_69),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_115),
.B(n_12),
.Y(n_161)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_80),
.A2(n_38),
.B1(n_35),
.B2(n_9),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_126),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_56),
.A2(n_35),
.B1(n_8),
.B2(n_11),
.Y(n_126)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

OR2x2_ASAP7_75t_SL g138 ( 
.A(n_104),
.B(n_51),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_138),
.B(n_143),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_139),
.A2(n_173),
.B1(n_174),
.B2(n_176),
.Y(n_203)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_61),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_147),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_170),
.B1(n_116),
.B2(n_113),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_90),
.B(n_66),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_149),
.B(n_157),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_64),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_150),
.B(n_171),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_102),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_160),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_77),
.B(n_70),
.C(n_74),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_113),
.B(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_93),
.B(n_8),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_12),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_161),
.B(n_162),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_78),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_130),
.B(n_13),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_167),
.B(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_103),
.B(n_67),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_13),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_13),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_111),
.B(n_14),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_103),
.B(n_81),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_177),
.C(n_178),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_97),
.B(n_14),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_14),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_106),
.B(n_15),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_152),
.A2(n_92),
.B1(n_123),
.B2(n_100),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_180),
.A2(n_187),
.B1(n_190),
.B2(n_192),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_147),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_152),
.A2(n_99),
.B1(n_100),
.B2(n_123),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_163),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_164),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_193),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_148),
.A2(n_99),
.B1(n_131),
.B2(n_128),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_159),
.A2(n_131),
.B1(n_128),
.B2(n_111),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_94),
.B(n_116),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_86),
.B1(n_124),
.B2(n_77),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_196),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_95),
.B1(n_86),
.B2(n_124),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_166),
.A2(n_94),
.B1(n_134),
.B2(n_95),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_166),
.A2(n_94),
.B1(n_117),
.B2(n_150),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_166),
.A2(n_165),
.B1(n_160),
.B2(n_138),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_165),
.A2(n_142),
.B1(n_136),
.B2(n_145),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_180),
.B1(n_192),
.B2(n_187),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_158),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_233),
.Y(n_240)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_195),
.B(n_140),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_216),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_163),
.C(n_169),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_232),
.C(n_200),
.Y(n_248)
);

NOR3xp33_ASAP7_75t_SL g218 ( 
.A(n_191),
.B(n_153),
.C(n_156),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_226),
.C(n_231),
.Y(n_245)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_219),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_229),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_208),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_228),
.B(n_237),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_179),
.B(n_155),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_181),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_156),
.C(n_164),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_164),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_205),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_236),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_212),
.B(n_206),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_182),
.B(n_183),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_183),
.B(n_182),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_213),
.B(n_190),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_236),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_230),
.A2(n_184),
.B1(n_193),
.B2(n_196),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_247),
.B1(n_235),
.B2(n_223),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_204),
.B1(n_211),
.B2(n_201),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_259),
.C(n_232),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_225),
.A2(n_200),
.B(n_186),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_250),
.A2(n_252),
.B(n_223),
.Y(n_267)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_215),
.A2(n_185),
.B(n_202),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_251),
.B(n_224),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_215),
.A2(n_198),
.B(n_186),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_255),
.B(n_228),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_198),
.C(n_202),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_251),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_261),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_237),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_262),
.B(n_264),
.Y(n_282)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_239),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_259),
.C(n_250),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_266),
.A2(n_269),
.B1(n_276),
.B2(n_241),
.Y(n_278)
);

XNOR2x1_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_271),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_221),
.Y(n_268)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_253),
.A2(n_235),
.B1(n_234),
.B2(n_222),
.Y(n_269)
);

NOR3xp33_ASAP7_75t_SL g286 ( 
.A(n_270),
.B(n_272),
.C(n_273),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_251),
.A2(n_231),
.B(n_214),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_242),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_217),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_275),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_249),
.B(n_216),
.Y(n_275)
);

A2O1A1O1Ixp25_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_240),
.B(n_257),
.C(n_252),
.D(n_253),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_278),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_248),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_254),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_274),
.C(n_268),
.Y(n_291)
);

A2O1A1O1Ixp25_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_245),
.B(n_254),
.C(n_218),
.D(n_244),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_267),
.C(n_260),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_296),
.B1(n_280),
.B2(n_288),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_291),
.B(n_292),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_266),
.C(n_271),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_282),
.A2(n_269),
.B1(n_261),
.B2(n_270),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_294),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_286),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_287),
.A2(n_276),
.B(n_254),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_298),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_273),
.C(n_272),
.Y(n_298)
);

AOI211xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_278),
.B(n_283),
.C(n_286),
.Y(n_299)
);

AO21x1_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_256),
.B(n_243),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_303),
.A2(n_291),
.B(n_297),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_280),
.B1(n_277),
.B2(n_247),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_296),
.A2(n_279),
.B1(n_263),
.B2(n_258),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_309),
.B(n_311),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_301),
.A2(n_279),
.B(n_258),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_246),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_312),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_256),
.C(n_207),
.Y(n_312)
);

OAI321xp33_ASAP7_75t_L g313 ( 
.A1(n_308),
.A2(n_306),
.A3(n_299),
.B1(n_302),
.B2(n_305),
.C(n_304),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_313),
.A2(n_302),
.B(n_243),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_308),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_315),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_318),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_316),
.A3(n_314),
.B1(n_226),
.B2(n_220),
.C1(n_219),
.C2(n_222),
.Y(n_320)
);

NOR3xp33_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_207),
.C(n_185),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_319),
.Y(n_322)
);


endmodule