module fake_netlist_6_144_n_4749 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_305, n_72, n_532, n_173, n_250, n_372, n_468, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_521, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4749);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_532;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4749;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_4730;
wire n_801;
wire n_4452;
wire n_3766;
wire n_1613;
wire n_4598;
wire n_1458;
wire n_2576;
wire n_1234;
wire n_3254;
wire n_3684;
wire n_4649;
wire n_1674;
wire n_1199;
wire n_3392;
wire n_4670;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_4620;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_4738;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_700;
wire n_3783;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_4504;
wire n_3844;
wire n_4388;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_4395;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4517;
wire n_4168;
wire n_783;
wire n_4372;
wire n_2451;
wire n_1738;
wire n_4490;
wire n_2243;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_798;
wire n_3088;
wire n_3443;
wire n_3257;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_4686;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_4699;
wire n_2051;
wire n_4370;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_2847;
wire n_2557;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1009;
wire n_1930;
wire n_1743;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_2997;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1238;
wire n_4092;
wire n_4645;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_4578;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4591;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_4702;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_1371;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_873;
wire n_3946;
wire n_1985;
wire n_4213;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_4474;
wire n_852;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_4531;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_2247;
wire n_544;
wire n_1711;
wire n_1078;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_4666;
wire n_2470;
wire n_2321;
wire n_4446;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_836;
wire n_3345;
wire n_2074;
wire n_4417;
wire n_2447;
wire n_2919;
wire n_4501;
wire n_3678;
wire n_3440;
wire n_4617;
wire n_4733;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_4724;
wire n_945;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_4555;
wire n_4743;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_4696;
wire n_4692;
wire n_1572;
wire n_4308;
wire n_616;
wire n_658;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2510;
wire n_1954;
wire n_2044;
wire n_2739;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_3023;
wire n_1735;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_4325;
wire n_4602;
wire n_2212;
wire n_3929;
wire n_758;
wire n_3494;
wire n_3063;
wire n_3048;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_1455;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_4722;
wire n_4606;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_4187;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_538;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3737;
wire n_3624;
wire n_3077;
wire n_3979;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_4556;
wire n_539;
wire n_4563;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_4687;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_4619;
wire n_2378;
wire n_887;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_4414;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_4600;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_4646;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_4262;
wire n_4392;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_659;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_913;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4071;
wire n_4255;
wire n_4403;
wire n_3506;
wire n_4729;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_4605;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_4549;
wire n_4575;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_2300;
wire n_1986;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_564;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4349;
wire n_824;
wire n_686;
wire n_4102;
wire n_4297;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_577;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_4662;
wire n_1843;
wire n_619;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_4227;
wire n_2778;
wire n_2850;
wire n_572;
wire n_4314;
wire n_1909;
wire n_2080;
wire n_813;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_606;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_3910;
wire n_1699;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4415;
wire n_4296;
wire n_4009;
wire n_2633;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_630;
wire n_2059;
wire n_4507;
wire n_2198;
wire n_3319;
wire n_541;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_4499;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_4677;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_792;
wire n_3949;
wire n_4364;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_4732;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_4393;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_982;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_2832;
wire n_4581;
wire n_4226;
wire n_549;
wire n_1762;
wire n_4641;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_932;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_4377;
wire n_3446;
wire n_4158;
wire n_4366;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_905;
wire n_3630;
wire n_4698;
wire n_3518;
wire n_4445;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_993;
wire n_2692;
wire n_3842;
wire n_689;
wire n_3248;
wire n_2031;
wire n_4544;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_4477;
wire n_966;
wire n_3888;
wire n_4511;
wire n_2908;
wire n_3168;
wire n_764;
wire n_4468;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4337;
wire n_4161;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3055;
wire n_3092;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_4369;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_4454;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_4742;
wire n_1014;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_4520;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_4502;
wire n_882;
wire n_4503;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_586;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1875;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_4375;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4526;
wire n_4277;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1950;
wire n_1726;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_4441;
wire n_4613;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_4478;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_4717;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_4585;
wire n_4731;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_702;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_2254;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_4467;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_4427;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_4485;
wire n_4386;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_4681;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4523;
wire n_4220;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_690;
wire n_2347;
wire n_835;
wire n_2092;
wire n_1886;
wire n_1654;
wire n_816;
wire n_4371;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_4552;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_4043;
wire n_4673;
wire n_825;
wire n_4313;
wire n_728;
wire n_4353;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_4607;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_4381;
wire n_1624;
wire n_1124;
wire n_3873;
wire n_3983;
wire n_2980;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_4510;
wire n_696;
wire n_1515;
wire n_4473;
wire n_961;
wire n_4356;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_593;
wire n_4169;
wire n_4055;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_3271;
wire n_950;
wire n_4248;
wire n_2812;
wire n_4518;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_4361;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_4589;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_4367;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_4560;
wire n_590;
wire n_4737;
wire n_4685;
wire n_4394;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_4675;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_2431;
wire n_3073;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_1634;
wire n_2078;
wire n_3252;
wire n_2932;
wire n_595;
wire n_627;
wire n_3253;
wire n_1779;
wire n_1465;
wire n_3337;
wire n_3431;
wire n_3450;
wire n_1767;
wire n_3209;
wire n_4002;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_4603;
wire n_1391;
wire n_4663;
wire n_1523;
wire n_2558;
wire n_2893;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_4697;
wire n_2954;
wire n_3477;
wire n_4288;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4289;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_815;
wire n_3953;
wire n_1100;
wire n_4588;
wire n_585;
wire n_4653;
wire n_1487;
wire n_4435;
wire n_2691;
wire n_3421;
wire n_2913;
wire n_840;
wire n_3614;
wire n_874;
wire n_4471;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_4728;
wire n_898;
wire n_4385;
wire n_1952;
wire n_865;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_2535;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_4191;
wire n_4636;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_4701;
wire n_4651;
wire n_1451;
wire n_3941;
wire n_639;
wire n_963;
wire n_2767;
wire n_794;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_4576;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_4615;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_872;
wire n_1139;
wire n_1714;
wire n_3922;
wire n_3179;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_542;
wire n_2897;
wire n_644;
wire n_682;
wire n_2537;
wire n_847;
wire n_851;
wire n_3970;
wire n_4389;
wire n_4483;
wire n_4345;
wire n_2554;
wire n_996;
wire n_4661;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_3171;
wire n_1913;
wire n_791;
wire n_4621;
wire n_4216;
wire n_3608;
wire n_4540;
wire n_837;
wire n_4315;
wire n_4664;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_4713;
wire n_4098;
wire n_4021;
wire n_4476;
wire n_765;
wire n_987;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_4688;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_4674;
wire n_2191;
wire n_2717;
wire n_1723;
wire n_4481;
wire n_1246;
wire n_4528;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_4475;
wire n_899;
wire n_738;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_3580;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_705;
wire n_3775;
wire n_3537;
wire n_4669;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_4443;
wire n_3887;
wire n_4634;
wire n_1022;
wire n_614;
wire n_2307;
wire n_2069;
wire n_3704;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_4123;
wire n_1431;
wire n_4096;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_4587;
wire n_4286;
wire n_3119;
wire n_1809;
wire n_4280;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_4379;
wire n_3731;
wire n_1822;
wire n_947;
wire n_2936;
wire n_3224;
wire n_4718;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_4525;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_4218;
wire n_4440;
wire n_4402;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_2848;
wire n_1849;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_4541;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4551;
wire n_4264;
wire n_4484;
wire n_2857;
wire n_3693;
wire n_4497;
wire n_3788;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_4459;
wire n_1299;
wire n_4545;
wire n_4708;
wire n_2896;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_4627;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3325;
wire n_3203;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_4464;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_4624;
wire n_2837;
wire n_4175;
wire n_4700;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_4659;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_2127;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_4455;
wire n_4453;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_4514;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_1507;
wire n_2482;
wire n_552;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4564;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2424;
wire n_2296;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_4487;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_623;
wire n_1048;
wire n_1398;
wire n_1201;
wire n_884;
wire n_716;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_4592;
wire n_4573;
wire n_2589;
wire n_4535;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_3393;
wire n_683;
wire n_811;
wire n_2442;
wire n_1207;
wire n_3627;
wire n_3451;
wire n_1791;
wire n_1368;
wire n_3480;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_4695;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_4401;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_4368;
wire n_1478;
wire n_589;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2581;
wire n_1363;
wire n_2294;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3591;
wire n_767;
wire n_3641;
wire n_1314;
wire n_600;
wire n_964;
wire n_1837;
wire n_2218;
wire n_831;
wire n_2788;
wire n_4533;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_1410;
wire n_4746;
wire n_2389;
wire n_1440;
wire n_2892;
wire n_2132;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1564;
wire n_1736;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_4658;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_3909;
wire n_3944;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2323;
wire n_1220;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2301;
wire n_2209;
wire n_3582;
wire n_4665;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_4431;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_4387;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_4633;
wire n_4654;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_642;
wire n_995;
wire n_2329;
wire n_1092;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_4584;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_4362;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_1784;
wire n_2990;
wire n_3847;
wire n_1286;
wire n_1775;
wire n_2115;
wire n_1773;
wire n_4430;
wire n_2552;
wire n_2410;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_1093;
wire n_4428;
wire n_4597;
wire n_1783;
wire n_1533;
wire n_2929;
wire n_1597;
wire n_2780;
wire n_3323;
wire n_3226;
wire n_3364;
wire n_4020;
wire n_4176;
wire n_4489;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_4404;
wire n_651;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_1531;
wire n_4618;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_4261;
wire n_1745;
wire n_4679;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_4496;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_4513;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_3646;
wire n_2801;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_4706;
wire n_2648;
wire n_4747;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_4570;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_3188;
wire n_1459;
wire n_3742;
wire n_4410;
wire n_1892;
wire n_2462;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4056;
wire n_1617;
wire n_4034;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_4622;
wire n_4721;
wire n_3093;
wire n_3175;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_4693;
wire n_2928;
wire n_4206;
wire n_4448;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_3284;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_1881;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_906;
wire n_2289;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2863;
wire n_3299;
wire n_1419;
wire n_1390;
wire n_3663;
wire n_4132;
wire n_2995;
wire n_2955;
wire n_1731;
wire n_2158;
wire n_3360;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_4614;
wire n_4609;
wire n_1437;
wire n_4438;
wire n_2135;
wire n_3956;
wire n_4707;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4676;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_4355;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_4422;
wire n_3917;
wire n_663;
wire n_2803;
wire n_3314;
wire n_2100;
wire n_856;
wire n_3525;
wire n_3016;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2993;
wire n_3688;
wire n_3566;
wire n_3004;
wire n_4647;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_4126;
wire n_1129;
wire n_3870;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_2181;
wire n_1995;
wire n_1594;
wire n_3751;
wire n_664;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_4632;
wire n_1429;
wire n_4655;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_4470;
wire n_587;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_4546;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_4583;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_4704;
wire n_4714;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_828;
wire n_2142;
wire n_4067;
wire n_4357;
wire n_4252;
wire n_607;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_4509;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_2327;
wire n_820;
wire n_951;
wire n_4374;
wire n_2201;
wire n_725;
wire n_952;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_4668;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4635;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3250;
wire n_1934;
wire n_3276;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_4582;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_617;
wire n_3886;
wire n_2924;
wire n_807;
wire n_845;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_4420;
wire n_4710;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_4574;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3926;
wire n_3797;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_4690;
wire n_1187;
wire n_4405;
wire n_610;
wire n_4234;
wire n_4413;
wire n_4304;
wire n_1403;
wire n_1669;
wire n_4558;
wire n_1852;
wire n_4488;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_4211;
wire n_4667;
wire n_4182;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_621;
wire n_1037;
wire n_1397;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_923;
wire n_1409;
wire n_4230;
wire n_4656;
wire n_1841;
wire n_4660;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_4637;
wire n_4274;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4270;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_4397;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_4155;
wire n_2740;
wire n_746;
wire n_4238;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_4611;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_3042;
wire n_1356;
wire n_1589;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_4610;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_4472;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_3249;
wire n_1320;
wire n_2716;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_4725;
wire n_4590;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_4406;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_4380;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_4398;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_3238;
wire n_2472;
wire n_1262;
wire n_2171;
wire n_1213;
wire n_1891;
wire n_2235;
wire n_3529;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4192;
wire n_4109;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_4565;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4159;
wire n_4195;
wire n_4567;
wire n_3784;
wire n_2298;
wire n_2326;
wire n_782;
wire n_1539;
wire n_4554;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_4586;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_4595;
wire n_4626;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4174;
wire n_2964;
wire n_1870;
wire n_4144;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_4734;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_662;
wire n_3475;
wire n_4442;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_4434;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_4680;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_711;
wire n_579;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_4515;
wire n_4689;
wire n_3845;
wire n_4616;
wire n_1682;
wire n_2017;
wire n_4516;
wire n_1695;
wire n_2699;
wire n_2046;
wire n_2272;
wire n_3029;
wire n_2200;
wire n_1828;
wire n_4547;
wire n_4258;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_4548;
wire n_4643;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_3878;
wire n_4601;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_4623;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_4553;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_4739;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_2479;
wire n_3050;
wire n_1823;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_4135;
wire n_2871;
wire n_4279;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_3858;
wire n_1845;
wire n_4183;
wire n_1489;
wire n_4321;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_543;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_4644;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_4040;
wire n_4561;
wire n_804;
wire n_4461;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4209;
wire n_4111;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_879;
wire n_959;
wire n_2310;
wire n_4608;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_4716;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_799;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_2195;
wire n_1633;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_3528;
wire n_4682;
wire n_3489;
wire n_4571;
wire n_4343;
wire n_2835;
wire n_4715;
wire n_4530;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_4694;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_4672;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_652;
wire n_2154;
wire n_2727;
wire n_3377;
wire n_4604;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_4378;
wire n_4407;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_3762;
wire n_3469;
wire n_3932;
wire n_2266;
wire n_2960;
wire n_3958;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_4519;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_4358;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_4524;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_4469;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_2083;
wire n_1269;
wire n_1931;
wire n_2834;
wire n_4572;
wire n_3207;
wire n_2668;
wire n_672;
wire n_4424;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_655;
wire n_4726;
wire n_706;
wire n_1045;
wire n_1794;
wire n_786;
wire n_1650;
wire n_1962;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_4736;
wire n_4317;
wire n_834;
wire n_4493;
wire n_4723;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_743;
wire n_766;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2671;
wire n_2885;
wire n_2761;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_2888;
wire n_3711;
wire n_3776;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_4650;
wire n_660;
wire n_2062;
wire n_4539;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_4421;
wire n_4719;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_4498;
wire n_2070;
wire n_2588;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_4492;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_817;
wire n_4423;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_1476;
wire n_841;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_4376;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_4203;
wire n_3808;
wire n_1742;
wire n_3190;
wire n_4505;
wire n_4657;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_4365;
wire n_1826;
wire n_566;
wire n_1023;
wire n_2951;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_4512;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_853;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_4542;
wire n_3199;
wire n_2931;
wire n_875;
wire n_680;
wire n_4462;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_4450;
wire n_4536;
wire n_4741;
wire n_4543;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_4630;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_4550;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_4652;
wire n_3503;
wire n_3160;
wire n_2796;
wire n_1065;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_4534;
wire n_1536;
wire n_3846;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_4408;
wire n_4577;
wire n_1132;
wire n_4748;
wire n_643;
wire n_698;
wire n_1074;
wire n_4439;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_4639;
wire n_2787;
wire n_2969;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_4494;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_4295;
wire n_1120;
wire n_832;
wire n_1583;
wire n_4480;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_2946;
wire n_2746;
wire n_814;
wire n_4579;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_691;
wire n_535;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3860;
wire n_3583;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3701;
wire n_3154;
wire n_4027;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_3473;
wire n_4557;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_4432;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_4352;
wire n_744;
wire n_971;
wire n_4391;
wire n_4416;
wire n_2702;
wire n_3241;
wire n_946;
wire n_4593;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_4342;
wire n_4465;
wire n_3622;
wire n_4568;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_4495;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_3551;
wire n_4436;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_4569;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_4559;
wire n_1347;
wire n_4106;
wire n_795;
wire n_3604;
wire n_1501;
wire n_1221;
wire n_3334;
wire n_4373;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_647;
wire n_4160;
wire n_4231;
wire n_844;
wire n_4711;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_4740;
wire n_2117;
wire n_2234;
wire n_4631;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2465;
wire n_1112;
wire n_2275;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_4720;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_2255;
wire n_2112;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_3486;
wire n_4678;
wire n_4086;
wire n_908;
wire n_752;
wire n_2649;
wire n_2721;
wire n_944;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_576;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_2862;
wire n_2615;
wire n_2265;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_4625;
wire n_4409;
wire n_2744;
wire n_4309;
wire n_4363;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_4521;
wire n_2437;
wire n_2444;
wire n_839;
wire n_1215;
wire n_2743;
wire n_3962;
wire n_4629;
wire n_4638;
wire n_708;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_4166;
wire n_626;
wire n_990;
wire n_1500;
wire n_1537;
wire n_779;
wire n_1821;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_2242;
wire n_1266;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4744;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3256;
wire n_3868;
wire n_1276;
wire n_3802;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4142;
wire n_2466;
wire n_2111;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3697;
wire n_3643;
wire n_771;
wire n_1584;
wire n_2425;
wire n_924;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_4265;
wire n_3680;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_4532;
wire n_719;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_4383;
wire n_4491;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_2666;
wire n_4105;
wire n_1851;
wire n_1585;
wire n_1799;
wire n_1090;
wire n_2564;
wire n_2147;
wire n_592;
wire n_4486;
wire n_4244;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_829;
wire n_1156;
wire n_1362;
wire n_4259;
wire n_3123;
wire n_2600;
wire n_984;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_4612;
wire n_868;
wire n_3038;
wire n_570;
wire n_3086;
wire n_2033;
wire n_859;
wire n_735;
wire n_4104;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_3285;
wire n_4208;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_4529;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_4537;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_4346;
wire n_4351;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_4316;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_4640;
wire n_3521;
wire n_3233;
wire n_4599;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_4437;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4390;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_4628;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_4396;
wire n_4508;
wire n_1763;
wire n_4594;
wire n_1998;
wire n_3066;
wire n_4727;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_3989;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_4451;
wire n_1606;
wire n_4332;
wire n_810;
wire n_4108;
wire n_1133;
wire n_4460;
wire n_635;
wire n_1194;
wire n_3374;
wire n_4429;
wire n_4506;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_4538;
wire n_2640;
wire n_3695;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_4293;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_553;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_849;
wire n_3383;
wire n_3709;
wire n_4684;
wire n_753;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_3187;
wire n_2540;
wire n_4412;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_4580;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_4522;
wire n_4148;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_679;
wire n_4057;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_4263;
wire n_1819;
wire n_2055;
wire n_1260;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_4447;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_3017;
wire n_1890;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_3903;
wire n_730;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_2333;
wire n_1868;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_4463;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3896;
wire n_2774;
wire n_3815;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_4648;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3333;
wire n_3274;
wire n_3186;
wire n_640;
wire n_4129;
wire n_1322;
wire n_4457;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_722;
wire n_4500;
wire n_862;
wire n_2105;
wire n_3079;
wire n_4360;
wire n_3085;
wire n_2098;
wire n_4433;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3584;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_4745;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4566;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_4482;
wire n_4275;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_900;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_4426;
wire n_2912;
wire n_827;
wire n_4703;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_4425;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_4449;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_4030;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_439),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_265),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_339),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_136),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_523),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_258),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_451),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_351),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_504),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_206),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_58),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_514),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_457),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_284),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_36),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_482),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_378),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_7),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_417),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_527),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_500),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_506),
.Y(n_554)
);

BUFx10_ASAP7_75t_L g555 ( 
.A(n_425),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_365),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_178),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_336),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_519),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_388),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_230),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_200),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_5),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_418),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_144),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_278),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_384),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_453),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_287),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_467),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_294),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_13),
.Y(n_572)
);

BUFx2_ASAP7_75t_R g573 ( 
.A(n_230),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_250),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_526),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_39),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_359),
.Y(n_577)
);

BUFx10_ASAP7_75t_L g578 ( 
.A(n_472),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_204),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_325),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_375),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_12),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_139),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_77),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_125),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_495),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_405),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_398),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_316),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_505),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_221),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_445),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_461),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_25),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_242),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_386),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_229),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_36),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_216),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_247),
.Y(n_600)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_414),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_124),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_218),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_332),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_24),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_358),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_328),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_125),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_236),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_390),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_165),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_420),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_471),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_120),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_304),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_222),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_272),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_383),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_130),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_401),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_73),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_355),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_222),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_77),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_320),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_160),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_138),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_431),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_529),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_185),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_291),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_473),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_124),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_442),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_183),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_489),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_91),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_213),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_174),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_63),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_164),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_464),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_511),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_128),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_501),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_496),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_479),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_10),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_337),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_34),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_433),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_340),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_347),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_18),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_306),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_186),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_324),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_8),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_137),
.Y(n_659)
);

BUFx2_ASAP7_75t_SL g660 ( 
.A(n_338),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_382),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_158),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_271),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_117),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_466),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_465),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_204),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_276),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_183),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_173),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_211),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_228),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_42),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_400),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_288),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_395),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_245),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_81),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_91),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_281),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_12),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_481),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_136),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_406),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_193),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_93),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_456),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_427),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_32),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_223),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_39),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_233),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_364),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_33),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_190),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_202),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_282),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_517),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_497),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_97),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_155),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_402),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_530),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_237),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_396),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_58),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_205),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_102),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_54),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_34),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_235),
.Y(n_711)
);

CKINVDCx14_ASAP7_75t_R g712 ( 
.A(n_6),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_107),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_28),
.Y(n_714)
);

BUFx10_ASAP7_75t_L g715 ( 
.A(n_385),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_148),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_333),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_71),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_486),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_470),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_193),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_478),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_253),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_25),
.Y(n_724)
);

CKINVDCx14_ASAP7_75t_R g725 ( 
.A(n_221),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_86),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_408),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_38),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_455),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_99),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_32),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_51),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_363),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_196),
.Y(n_734)
);

BUFx10_ASAP7_75t_L g735 ( 
.A(n_444),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_354),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_352),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_528),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_14),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_518),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_89),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_493),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_397),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_318),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_210),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_205),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_220),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_515),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_286),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_341),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_255),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_73),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_119),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_525),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_61),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_68),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_132),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_452),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_298),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_319),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_208),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_147),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_17),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_192),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_380),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_379),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_361),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_95),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_476),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_113),
.Y(n_770)
);

BUFx10_ASAP7_75t_L g771 ( 
.A(n_262),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_454),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_423),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_175),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_321),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_84),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_176),
.Y(n_777)
);

CKINVDCx14_ASAP7_75t_R g778 ( 
.A(n_75),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_463),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_447),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_426),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_60),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_432),
.Y(n_783)
);

INVx1_ASAP7_75t_SL g784 ( 
.A(n_389),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_374),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_97),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_7),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_201),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_200),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_317),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_160),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_297),
.Y(n_792)
);

CKINVDCx16_ASAP7_75t_R g793 ( 
.A(n_104),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_203),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_508),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_53),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_263),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_20),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_260),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_213),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_177),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_83),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_13),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_299),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_268),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_399),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_111),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_441),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_47),
.Y(n_809)
);

BUFx5_ASAP7_75t_L g810 ( 
.A(n_458),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_43),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_367),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_121),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_71),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_201),
.Y(n_815)
);

CKINVDCx14_ASAP7_75t_R g816 ( 
.A(n_135),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_251),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_231),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_422),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_258),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_412),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_278),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_218),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_507),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_531),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_311),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_81),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_323),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_309),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_43),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_498),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_8),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_30),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_236),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_250),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_233),
.Y(n_836)
);

BUFx5_ASAP7_75t_L g837 ( 
.A(n_108),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_169),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_217),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_197),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_301),
.Y(n_841)
);

CKINVDCx16_ASAP7_75t_R g842 ( 
.A(n_182),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_326),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_56),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_74),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_238),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_107),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_421),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_219),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_371),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_313),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_212),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_357),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_38),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_305),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_303),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_211),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_460),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_366),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_123),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_438),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_103),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_262),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_231),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_161),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_260),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_334),
.Y(n_867)
);

BUFx10_ASAP7_75t_L g868 ( 
.A(n_40),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_20),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_387),
.Y(n_870)
);

BUFx10_ASAP7_75t_L g871 ( 
.A(n_122),
.Y(n_871)
);

BUFx10_ASAP7_75t_L g872 ( 
.A(n_145),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_302),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_404),
.Y(n_874)
);

CKINVDCx16_ASAP7_75t_R g875 ( 
.A(n_105),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_314),
.Y(n_876)
);

CKINVDCx14_ASAP7_75t_R g877 ( 
.A(n_134),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_295),
.Y(n_878)
);

CKINVDCx14_ASAP7_75t_R g879 ( 
.A(n_129),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_188),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_407),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_223),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_448),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_82),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_449),
.Y(n_885)
);

BUFx10_ASAP7_75t_L g886 ( 
.A(n_148),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_217),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_377),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_219),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_151),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_255),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_169),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_67),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_167),
.Y(n_894)
);

CKINVDCx16_ASAP7_75t_R g895 ( 
.A(n_149),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_369),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_83),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_79),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_203),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_440),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_289),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_310),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_424),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_480),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_435),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_66),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_238),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_163),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_232),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_403),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_416),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_155),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_41),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_273),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_104),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_487),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_512),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_63),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_162),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_185),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_349),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_207),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_192),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_28),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_120),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_206),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_413),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_837),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_746),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_837),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_712),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_837),
.Y(n_932)
);

NOR2xp67_ASAP7_75t_L g933 ( 
.A(n_747),
.B(n_0),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_567),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_725),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_837),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_837),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_837),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_837),
.Y(n_939)
);

INVxp33_ASAP7_75t_SL g940 ( 
.A(n_692),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_543),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_837),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_747),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_540),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_540),
.Y(n_945)
);

INVxp33_ASAP7_75t_L g946 ( 
.A(n_739),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_778),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_546),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_546),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_746),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_554),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_551),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_551),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_553),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_553),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_762),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_564),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_564),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_571),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_571),
.Y(n_960)
);

CKINVDCx14_ASAP7_75t_R g961 ( 
.A(n_816),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_877),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_542),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_577),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_577),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_580),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_557),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_580),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_572),
.Y(n_969)
);

INVxp67_ASAP7_75t_SL g970 ( 
.A(n_698),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_762),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_836),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_747),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_599),
.Y(n_974)
);

INVxp33_ASAP7_75t_SL g975 ( 
.A(n_836),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_606),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_606),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_607),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_607),
.Y(n_979)
);

CKINVDCx14_ASAP7_75t_R g980 ( 
.A(n_879),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_622),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_567),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_622),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_629),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_793),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_609),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_868),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_629),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_643),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_643),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_641),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_655),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_655),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_554),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_661),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_793),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_842),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_661),
.Y(n_998)
);

INVxp67_ASAP7_75t_SL g999 ( 
.A(n_760),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_842),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_542),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_875),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_542),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_875),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_895),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_542),
.Y(n_1006)
);

CKINVDCx16_ASAP7_75t_R g1007 ( 
.A(n_895),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_542),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_534),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_884),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_884),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_884),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_884),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_884),
.Y(n_1014)
);

INVxp33_ASAP7_75t_SL g1015 ( 
.A(n_561),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_897),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_641),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_897),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_897),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_897),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_897),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_562),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_908),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_908),
.Y(n_1024)
);

INVxp33_ASAP7_75t_L g1025 ( 
.A(n_536),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_908),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_908),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_563),
.Y(n_1028)
);

INVxp33_ASAP7_75t_SL g1029 ( 
.A(n_565),
.Y(n_1029)
);

CKINVDCx16_ASAP7_75t_R g1030 ( 
.A(n_868),
.Y(n_1030)
);

INVxp67_ASAP7_75t_L g1031 ( 
.A(n_868),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_908),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_583),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_666),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_717),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_576),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_666),
.Y(n_1037)
);

INVxp33_ASAP7_75t_SL g1038 ( 
.A(n_579),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_582),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_688),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_688),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_705),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_705),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_717),
.Y(n_1044)
);

CKINVDCx14_ASAP7_75t_R g1045 ( 
.A(n_628),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_727),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_727),
.Y(n_1047)
);

CKINVDCx14_ASAP7_75t_R g1048 ( 
.A(n_628),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_662),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_737),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_585),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_737),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_748),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_748),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_766),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_591),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_554),
.Y(n_1057)
);

INVxp67_ASAP7_75t_L g1058 ( 
.A(n_871),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_766),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_594),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_767),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_767),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_595),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_769),
.Y(n_1064)
);

INVxp33_ASAP7_75t_L g1065 ( 
.A(n_536),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_602),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_769),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_603),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_773),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_773),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_608),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_806),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_871),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_671),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_616),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_619),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_806),
.Y(n_1077)
);

INVxp33_ASAP7_75t_L g1078 ( 
.A(n_538),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_621),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_819),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_819),
.Y(n_1081)
);

INVxp67_ASAP7_75t_SL g1082 ( 
.A(n_647),
.Y(n_1082)
);

INVxp33_ASAP7_75t_L g1083 ( 
.A(n_538),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_824),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_824),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_850),
.Y(n_1086)
);

CKINVDCx16_ASAP7_75t_R g1087 ( 
.A(n_871),
.Y(n_1087)
);

INVxp33_ASAP7_75t_L g1088 ( 
.A(n_547),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_850),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_855),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_623),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_627),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_855),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_867),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_867),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_810),
.Y(n_1096)
);

CKINVDCx16_ASAP7_75t_R g1097 ( 
.A(n_872),
.Y(n_1097)
);

INVxp67_ASAP7_75t_SL g1098 ( 
.A(n_647),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_870),
.Y(n_1099)
);

INVxp67_ASAP7_75t_SL g1100 ( 
.A(n_888),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_630),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_810),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_870),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_883),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_635),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_685),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_637),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_883),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_905),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_905),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_910),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_910),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_858),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_917),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_917),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_638),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_872),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_927),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_686),
.Y(n_1119)
);

CKINVDCx16_ASAP7_75t_R g1120 ( 
.A(n_872),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_927),
.Y(n_1121)
);

CKINVDCx16_ASAP7_75t_R g1122 ( 
.A(n_886),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_691),
.Y(n_1123)
);

INVxp67_ASAP7_75t_L g1124 ( 
.A(n_886),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_691),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_810),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_640),
.Y(n_1127)
);

CKINVDCx16_ASAP7_75t_R g1128 ( 
.A(n_886),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_810),
.Y(n_1129)
);

CKINVDCx14_ASAP7_75t_R g1130 ( 
.A(n_888),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_815),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_644),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_815),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_648),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_839),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_839),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_547),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_656),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_554),
.Y(n_1139)
);

INVxp67_ASAP7_75t_SL g1140 ( 
.A(n_858),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_923),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_901),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_663),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_901),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_923),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_925),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_925),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_904),
.Y(n_1148)
);

INVxp67_ASAP7_75t_SL g1149 ( 
.A(n_904),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_566),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_554),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_566),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_598),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_598),
.Y(n_1154)
);

NOR2xp67_ASAP7_75t_L g1155 ( 
.A(n_568),
.B(n_0),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_600),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_550),
.B(n_1),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_600),
.Y(n_1158)
);

INVxp67_ASAP7_75t_SL g1159 ( 
.A(n_568),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_611),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_611),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_614),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_614),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_810),
.Y(n_1164)
);

INVxp33_ASAP7_75t_SL g1165 ( 
.A(n_664),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_617),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_617),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_667),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_624),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_668),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_555),
.Y(n_1171)
);

INVxp33_ASAP7_75t_L g1172 ( 
.A(n_624),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_626),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_626),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_633),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_689),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_633),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_650),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_650),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_810),
.Y(n_1180)
);

CKINVDCx16_ASAP7_75t_R g1181 ( 
.A(n_771),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_654),
.Y(n_1182)
);

CKINVDCx16_ASAP7_75t_R g1183 ( 
.A(n_771),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_654),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_658),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_583),
.Y(n_1186)
);

INVxp67_ASAP7_75t_SL g1187 ( 
.A(n_568),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_658),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_673),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_555),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_678),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_679),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_669),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_669),
.Y(n_1194)
);

INVxp67_ASAP7_75t_SL g1195 ( 
.A(n_665),
.Y(n_1195)
);

INVxp67_ASAP7_75t_SL g1196 ( 
.A(n_610),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_670),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_670),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_681),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_672),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_672),
.B(n_1),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_694),
.Y(n_1202)
);

INVxp67_ASAP7_75t_SL g1203 ( 
.A(n_610),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_683),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_696),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_683),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_695),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_700),
.Y(n_1208)
);

INVxp33_ASAP7_75t_SL g1209 ( 
.A(n_701),
.Y(n_1209)
);

CKINVDCx16_ASAP7_75t_R g1210 ( 
.A(n_771),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_695),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_710),
.Y(n_1212)
);

CKINVDCx16_ASAP7_75t_R g1213 ( 
.A(n_771),
.Y(n_1213)
);

INVxp33_ASAP7_75t_SL g1214 ( 
.A(n_704),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_710),
.Y(n_1215)
);

CKINVDCx20_ASAP7_75t_R g1216 ( 
.A(n_786),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_718),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_799),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_718),
.Y(n_1219)
);

INVxp33_ASAP7_75t_L g1220 ( 
.A(n_724),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_706),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_707),
.Y(n_1222)
);

INVxp67_ASAP7_75t_SL g1223 ( 
.A(n_646),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_724),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_741),
.Y(n_1225)
);

INVxp33_ASAP7_75t_SL g1226 ( 
.A(n_708),
.Y(n_1226)
);

INVxp67_ASAP7_75t_SL g1227 ( 
.A(n_646),
.Y(n_1227)
);

INVxp33_ASAP7_75t_L g1228 ( 
.A(n_741),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_709),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_713),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_751),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_751),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_756),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_756),
.Y(n_1234)
);

INVxp33_ASAP7_75t_L g1235 ( 
.A(n_761),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_761),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_605),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_763),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_763),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_721),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_605),
.Y(n_1241)
);

CKINVDCx14_ASAP7_75t_R g1242 ( 
.A(n_555),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_764),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_764),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_631),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_800),
.Y(n_1246)
);

INVxp33_ASAP7_75t_L g1247 ( 
.A(n_800),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_723),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_834),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_834),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_838),
.Y(n_1251)
);

INVxp67_ASAP7_75t_SL g1252 ( 
.A(n_651),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_838),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_846),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_846),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_852),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_852),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_854),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_854),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_864),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_728),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_864),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_578),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_811),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_730),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_866),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_866),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_880),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_880),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_892),
.Y(n_1270)
);

INVxp33_ASAP7_75t_SL g1271 ( 
.A(n_731),
.Y(n_1271)
);

BUFx2_ASAP7_75t_L g1272 ( 
.A(n_732),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_892),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_918),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_918),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_651),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_639),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_734),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_812),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_812),
.Y(n_1280)
);

NOR2xp67_ASAP7_75t_L g1281 ( 
.A(n_776),
.B(n_2),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_821),
.Y(n_1282)
);

INVxp33_ASAP7_75t_SL g1283 ( 
.A(n_745),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_821),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_639),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_714),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_818),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_714),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_726),
.Y(n_1289)
);

INVxp67_ASAP7_75t_SL g1290 ( 
.A(n_894),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_898),
.Y(n_1291)
);

INVxp67_ASAP7_75t_SL g1292 ( 
.A(n_676),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_578),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_726),
.Y(n_1294)
);

BUFx12f_ASAP7_75t_L g1295 ( 
.A(n_931),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_961),
.B(n_578),
.Y(n_1296)
);

CKINVDCx8_ASAP7_75t_R g1297 ( 
.A(n_1007),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1292),
.B(n_1140),
.Y(n_1298)
);

INVx5_ASAP7_75t_L g1299 ( 
.A(n_951),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_963),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_980),
.B(n_715),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_951),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_951),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_951),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1144),
.B(n_676),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1045),
.B(n_715),
.Y(n_1306)
);

BUFx8_ASAP7_75t_SL g1307 ( 
.A(n_941),
.Y(n_1307)
);

INVx5_ASAP7_75t_L g1308 ( 
.A(n_951),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_994),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_963),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1001),
.Y(n_1311)
);

BUFx12f_ASAP7_75t_L g1312 ( 
.A(n_931),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1001),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1159),
.B(n_631),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1149),
.B(n_533),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1187),
.B(n_631),
.Y(n_1316)
);

INVx4_ASAP7_75t_L g1317 ( 
.A(n_1009),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1003),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1048),
.B(n_715),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_991),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_985),
.Y(n_1321)
);

INVx5_ASAP7_75t_L g1322 ( 
.A(n_994),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_934),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1195),
.B(n_535),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1003),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_994),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_935),
.Y(n_1327)
);

BUFx12f_ASAP7_75t_L g1328 ( 
.A(n_935),
.Y(n_1328)
);

INVx4_ASAP7_75t_L g1329 ( 
.A(n_1009),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1130),
.B(n_601),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1006),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1157),
.B(n_631),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_994),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_934),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1006),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1142),
.B(n_537),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_994),
.Y(n_1337)
);

BUFx12f_ASAP7_75t_L g1338 ( 
.A(n_947),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1008),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1057),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1008),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1142),
.B(n_539),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_982),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1057),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1010),
.Y(n_1345)
);

INVx5_ASAP7_75t_L g1346 ( 
.A(n_1057),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_982),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1142),
.B(n_541),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1155),
.B(n_735),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1157),
.B(n_631),
.Y(n_1350)
);

BUFx12f_ASAP7_75t_L g1351 ( 
.A(n_947),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1010),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1082),
.B(n_625),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1057),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1057),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1098),
.B(n_645),
.Y(n_1356)
);

INVx4_ASAP7_75t_L g1357 ( 
.A(n_1022),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1035),
.B(n_544),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1242),
.B(n_735),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1011),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1011),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1139),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1035),
.B(n_545),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1028),
.B(n_735),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1044),
.B(n_548),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1044),
.B(n_549),
.Y(n_1366)
);

AND2x6_ASAP7_75t_L g1367 ( 
.A(n_928),
.B(n_780),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_SL g1368 ( 
.A(n_1181),
.B(n_573),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1100),
.B(n_653),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1063),
.B(n_735),
.Y(n_1370)
);

BUFx8_ASAP7_75t_SL g1371 ( 
.A(n_941),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1113),
.B(n_552),
.Y(n_1372)
);

BUFx12f_ASAP7_75t_L g1373 ( 
.A(n_962),
.Y(n_1373)
);

BUFx12f_ASAP7_75t_L g1374 ( 
.A(n_962),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1091),
.B(n_744),
.Y(n_1375)
);

INVx5_ASAP7_75t_L g1376 ( 
.A(n_1139),
.Y(n_1376)
);

BUFx12f_ASAP7_75t_L g1377 ( 
.A(n_985),
.Y(n_1377)
);

BUFx8_ASAP7_75t_L g1378 ( 
.A(n_1208),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1113),
.B(n_556),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1012),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1196),
.B(n_765),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1012),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1092),
.B(n_784),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_970),
.B(n_558),
.Y(n_1384)
);

AND2x6_ASAP7_75t_L g1385 ( 
.A(n_928),
.B(n_780),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1013),
.Y(n_1386)
);

BUFx12f_ASAP7_75t_L g1387 ( 
.A(n_996),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1013),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_991),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1139),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_999),
.B(n_1290),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1203),
.B(n_559),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1107),
.B(n_921),
.Y(n_1393)
);

INVx5_ASAP7_75t_L g1394 ( 
.A(n_1139),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1014),
.Y(n_1395)
);

INVx5_ASAP7_75t_L g1396 ( 
.A(n_1139),
.Y(n_1396)
);

BUFx8_ASAP7_75t_L g1397 ( 
.A(n_1017),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1223),
.B(n_550),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_933),
.B(n_1227),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1014),
.Y(n_1400)
);

BUFx12f_ASAP7_75t_L g1401 ( 
.A(n_996),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1252),
.B(n_1148),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1016),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_943),
.B(n_780),
.Y(n_1404)
);

INVx4_ASAP7_75t_L g1405 ( 
.A(n_1022),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1171),
.B(n_1190),
.Y(n_1406)
);

BUFx12f_ASAP7_75t_L g1407 ( 
.A(n_997),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1016),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1151),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_940),
.B(n_574),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1116),
.B(n_1143),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_1151),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1018),
.Y(n_1413)
);

AND2x6_ASAP7_75t_L g1414 ( 
.A(n_942),
.B(n_780),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_943),
.B(n_780),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1036),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1018),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1151),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1151),
.Y(n_1419)
);

BUFx8_ASAP7_75t_L g1420 ( 
.A(n_1017),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_997),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_973),
.B(n_1019),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_973),
.B(n_807),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1000),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1151),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1171),
.B(n_560),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1019),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1020),
.B(n_807),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1020),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1000),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1190),
.B(n_569),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1189),
.B(n_570),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1245),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_940),
.B(n_574),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1021),
.B(n_659),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1240),
.B(n_575),
.Y(n_1436)
);

INVx5_ASAP7_75t_L g1437 ( 
.A(n_1245),
.Y(n_1437)
);

INVx5_ASAP7_75t_L g1438 ( 
.A(n_1245),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1015),
.B(n_659),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1245),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1123),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1015),
.B(n_803),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1245),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1021),
.B(n_803),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1023),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1023),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1024),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1029),
.B(n_830),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1024),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1026),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1026),
.Y(n_1451)
);

INVx5_ASAP7_75t_L g1452 ( 
.A(n_1186),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1027),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1027),
.Y(n_1454)
);

INVx5_ASAP7_75t_L g1455 ( 
.A(n_1186),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1248),
.B(n_581),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1032),
.B(n_830),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_SL g1458 ( 
.A(n_1183),
.B(n_1210),
.Y(n_1458)
);

INVx5_ASAP7_75t_L g1459 ( 
.A(n_1237),
.Y(n_1459)
);

INVx4_ASAP7_75t_L g1460 ( 
.A(n_1036),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1032),
.B(n_586),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1263),
.B(n_587),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1029),
.B(n_752),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1281),
.B(n_753),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1038),
.B(n_755),
.Y(n_1465)
);

CKINVDCx6p67_ASAP7_75t_R g1466 ( 
.A(n_1213),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1237),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_SL g1468 ( 
.A(n_975),
.B(n_588),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_944),
.B(n_589),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1241),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_945),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1241),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1263),
.B(n_1293),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1208),
.B(n_590),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1277),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1293),
.B(n_592),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_930),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1125),
.B(n_593),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_932),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1277),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1038),
.B(n_757),
.Y(n_1481)
);

CKINVDCx16_ASAP7_75t_R g1482 ( 
.A(n_1030),
.Y(n_1482)
);

INVx5_ASAP7_75t_L g1483 ( 
.A(n_1096),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_936),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1131),
.B(n_596),
.Y(n_1485)
);

AND2x6_ASAP7_75t_L g1486 ( 
.A(n_937),
.B(n_584),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1150),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_938),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1133),
.B(n_604),
.Y(n_1489)
);

BUFx12f_ASAP7_75t_L g1490 ( 
.A(n_1002),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_939),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1165),
.B(n_768),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_948),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_949),
.B(n_612),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1152),
.Y(n_1495)
);

BUFx8_ASAP7_75t_L g1496 ( 
.A(n_1145),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1153),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1002),
.Y(n_1498)
);

INVx6_ASAP7_75t_L g1499 ( 
.A(n_1087),
.Y(n_1499)
);

CKINVDCx16_ASAP7_75t_R g1500 ( 
.A(n_1097),
.Y(n_1500)
);

INVx5_ASAP7_75t_L g1501 ( 
.A(n_1102),
.Y(n_1501)
);

INVx4_ASAP7_75t_L g1502 ( 
.A(n_1039),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_952),
.B(n_613),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1276),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_953),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1154),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1279),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_954),
.B(n_615),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1135),
.B(n_620),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_955),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1039),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_957),
.B(n_632),
.Y(n_1512)
);

INVx2_ASAP7_75t_SL g1513 ( 
.A(n_1051),
.Y(n_1513)
);

INVx4_ASAP7_75t_L g1514 ( 
.A(n_1051),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1136),
.B(n_634),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1056),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1145),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_1156),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1165),
.B(n_1283),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1209),
.B(n_1283),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1280),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1004),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1229),
.B(n_642),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_SL g1524 ( 
.A(n_975),
.B(n_618),
.Y(n_1524)
);

NOR2x1_ASAP7_75t_L g1525 ( 
.A(n_1282),
.B(n_660),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_958),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_959),
.B(n_649),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1229),
.B(n_652),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_960),
.B(n_674),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1158),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1272),
.B(n_675),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1160),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1284),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1272),
.B(n_680),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_1161),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1162),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_SL g1537 ( 
.A(n_1120),
.B(n_636),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1209),
.B(n_770),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1141),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_964),
.B(n_682),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_946),
.B(n_684),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_965),
.B(n_687),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1004),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1146),
.B(n_697),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1214),
.B(n_1226),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1126),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_929),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1129),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1214),
.B(n_774),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1147),
.B(n_699),
.Y(n_1550)
);

INVx3_ASAP7_75t_L g1551 ( 
.A(n_1163),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_966),
.B(n_702),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1166),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1167),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1056),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1169),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_968),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_976),
.B(n_977),
.Y(n_1558)
);

XNOR2x2_ASAP7_75t_L g1559 ( 
.A(n_1176),
.B(n_597),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_978),
.B(n_979),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1060),
.B(n_719),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1173),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1174),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1005),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1060),
.B(n_720),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_981),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_950),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1164),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_983),
.B(n_729),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_1066),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1175),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_984),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1066),
.Y(n_1573)
);

BUFx12f_ASAP7_75t_L g1574 ( 
.A(n_1005),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_988),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_989),
.B(n_733),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1226),
.B(n_777),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_1177),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_990),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1178),
.Y(n_1580)
);

BUFx8_ASAP7_75t_SL g1581 ( 
.A(n_967),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_992),
.B(n_736),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1179),
.Y(n_1583)
);

INVxp33_ASAP7_75t_SL g1584 ( 
.A(n_1068),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1182),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1068),
.B(n_738),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1184),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1180),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_993),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1071),
.Y(n_1590)
);

INVx5_ASAP7_75t_L g1591 ( 
.A(n_1122),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_995),
.B(n_740),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_998),
.B(n_742),
.Y(n_1593)
);

BUFx8_ASAP7_75t_SL g1594 ( 
.A(n_967),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_971),
.Y(n_1595)
);

AND2x6_ASAP7_75t_L g1596 ( 
.A(n_1034),
.B(n_677),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_L g1597 ( 
.A(n_1185),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1033),
.Y(n_1598)
);

BUFx12f_ASAP7_75t_L g1599 ( 
.A(n_1071),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1075),
.B(n_1076),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1320),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1320),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1546),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1546),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1310),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1310),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1435),
.B(n_1037),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1311),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1399),
.B(n_1040),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1298),
.B(n_1271),
.Y(n_1610)
);

INVx1_ASAP7_75t_SL g1611 ( 
.A(n_1307),
.Y(n_1611)
);

BUFx4f_ASAP7_75t_L g1612 ( 
.A(n_1484),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1471),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1323),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1493),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1548),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1548),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1398),
.B(n_1041),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1398),
.B(n_1042),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1568),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1302),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1311),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1335),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1335),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1323),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1399),
.B(n_1043),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1505),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1399),
.B(n_1046),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1339),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1389),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1435),
.B(n_1047),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1510),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1302),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1389),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1302),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1526),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1557),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1566),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1435),
.B(n_1050),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1314),
.B(n_1316),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1314),
.B(n_1052),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1314),
.B(n_1053),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1541),
.Y(n_1643)
);

NOR2x1_ASAP7_75t_L g1644 ( 
.A(n_1317),
.B(n_657),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1568),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1517),
.Y(n_1646)
);

CKINVDCx20_ASAP7_75t_R g1647 ( 
.A(n_1307),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1334),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1588),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1444),
.B(n_1054),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1339),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_SL g1652 ( 
.A1(n_1410),
.A2(n_912),
.B1(n_915),
.B2(n_909),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1315),
.B(n_1271),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1572),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_1334),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1575),
.Y(n_1656)
);

INVx2_ASAP7_75t_SL g1657 ( 
.A(n_1517),
.Y(n_1657)
);

INVx3_ASAP7_75t_L g1658 ( 
.A(n_1302),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1341),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1588),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1579),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1477),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1547),
.B(n_1218),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1444),
.B(n_1055),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1341),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1345),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1345),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1444),
.B(n_1059),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1316),
.B(n_1061),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1477),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1303),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1303),
.Y(n_1672)
);

BUFx6f_ASAP7_75t_L g1673 ( 
.A(n_1303),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1479),
.Y(n_1674)
);

NOR2x1_ASAP7_75t_L g1675 ( 
.A(n_1317),
.B(n_693),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1479),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1343),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_L g1678 ( 
.A(n_1329),
.B(n_1357),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1316),
.B(n_1062),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1491),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1491),
.Y(n_1681)
);

AND2x2_ASAP7_75t_SL g1682 ( 
.A(n_1468),
.B(n_1201),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1324),
.B(n_1075),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1330),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1303),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1358),
.B(n_1076),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1336),
.B(n_1064),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1484),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1300),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1361),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1313),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1318),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1371),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1342),
.B(n_1067),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1325),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_SL g1696 ( 
.A(n_1297),
.B(n_703),
.Y(n_1696)
);

INVxp67_ASAP7_75t_L g1697 ( 
.A(n_1330),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1457),
.B(n_1069),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1363),
.B(n_1079),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1361),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1386),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1371),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1331),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1457),
.B(n_1070),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1352),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1360),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1380),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1386),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1348),
.B(n_1072),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1382),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1395),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_SL g1712 ( 
.A(n_1591),
.B(n_1128),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1457),
.B(n_1077),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1388),
.Y(n_1714)
);

CKINVDCx8_ASAP7_75t_R g1715 ( 
.A(n_1482),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1395),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1400),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1558),
.B(n_1080),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1381),
.B(n_1081),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1417),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1400),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1591),
.B(n_1079),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1326),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1484),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_SL g1725 ( 
.A(n_1591),
.B(n_722),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1343),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1484),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1365),
.B(n_1101),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1326),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1558),
.B(n_1084),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1326),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1347),
.B(n_1085),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1558),
.B(n_1423),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1403),
.Y(n_1734)
);

INVx3_ASAP7_75t_L g1735 ( 
.A(n_1326),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1347),
.B(n_1086),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1488),
.Y(n_1737)
);

INVxp67_ASAP7_75t_L g1738 ( 
.A(n_1463),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1488),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1461),
.B(n_1089),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1488),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1488),
.Y(n_1742)
);

INVx4_ASAP7_75t_L g1743 ( 
.A(n_1483),
.Y(n_1743)
);

OA21x2_ASAP7_75t_L g1744 ( 
.A1(n_1429),
.A2(n_1093),
.B(n_1090),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1441),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1403),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1441),
.Y(n_1747)
);

INVx3_ASAP7_75t_L g1748 ( 
.A(n_1337),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1408),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1408),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1423),
.B(n_1094),
.Y(n_1751)
);

CKINVDCx11_ASAP7_75t_R g1752 ( 
.A(n_1466),
.Y(n_1752)
);

AND2x6_ASAP7_75t_L g1753 ( 
.A(n_1332),
.B(n_1095),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1539),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1539),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1381),
.B(n_1099),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1337),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1413),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1392),
.B(n_1103),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1589),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1589),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1495),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1413),
.Y(n_1763)
);

NAND2xp33_ASAP7_75t_L g1764 ( 
.A(n_1486),
.B(n_1201),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1495),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1375),
.A2(n_1105),
.B1(n_1127),
.B2(n_1101),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_1337),
.Y(n_1767)
);

OA21x2_ASAP7_75t_L g1768 ( 
.A1(n_1445),
.A2(n_1350),
.B(n_1332),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1427),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1495),
.Y(n_1770)
);

AND2x6_ASAP7_75t_L g1771 ( 
.A(n_1332),
.B(n_1104),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1427),
.Y(n_1772)
);

INVx3_ASAP7_75t_L g1773 ( 
.A(n_1337),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1446),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1446),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1495),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1350),
.B(n_1108),
.Y(n_1777)
);

BUFx6f_ASAP7_75t_L g1778 ( 
.A(n_1340),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1366),
.B(n_1105),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1506),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1350),
.B(n_1109),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1451),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1461),
.B(n_1110),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1340),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1461),
.B(n_1111),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1451),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1454),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1522),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1353),
.B(n_1112),
.Y(n_1789)
);

NAND2xp33_ASAP7_75t_SL g1790 ( 
.A(n_1383),
.B(n_919),
.Y(n_1790)
);

AND3x2_ASAP7_75t_L g1791 ( 
.A(n_1359),
.B(n_972),
.C(n_956),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1353),
.B(n_1114),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_L g1793 ( 
.A(n_1340),
.Y(n_1793)
);

INVxp67_ASAP7_75t_L g1794 ( 
.A(n_1463),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1454),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1356),
.B(n_1115),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1404),
.B(n_1118),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1506),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1467),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1467),
.Y(n_1800)
);

AO21x2_ASAP7_75t_L g1801 ( 
.A1(n_1349),
.A2(n_1121),
.B(n_1188),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1467),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1467),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1404),
.B(n_1415),
.Y(n_1804)
);

AND2x6_ASAP7_75t_L g1805 ( 
.A(n_1306),
.B(n_1193),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1340),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1470),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1423),
.B(n_1033),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1506),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1506),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1518),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1393),
.B(n_1504),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1518),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1518),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1470),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1470),
.Y(n_1816)
);

BUFx6f_ASAP7_75t_L g1817 ( 
.A(n_1344),
.Y(n_1817)
);

AND2x4_ASAP7_75t_L g1818 ( 
.A(n_1404),
.B(n_1194),
.Y(n_1818)
);

BUFx2_ASAP7_75t_L g1819 ( 
.A(n_1596),
.Y(n_1819)
);

BUFx3_ASAP7_75t_L g1820 ( 
.A(n_1415),
.Y(n_1820)
);

BUFx6f_ASAP7_75t_L g1821 ( 
.A(n_1344),
.Y(n_1821)
);

BUFx6f_ASAP7_75t_L g1822 ( 
.A(n_1344),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1518),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1344),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1470),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1532),
.Y(n_1826)
);

BUFx6f_ASAP7_75t_L g1827 ( 
.A(n_1354),
.Y(n_1827)
);

INVx3_ASAP7_75t_L g1828 ( 
.A(n_1354),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1522),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1354),
.Y(n_1830)
);

OAI21x1_ASAP7_75t_L g1831 ( 
.A1(n_1305),
.A2(n_1286),
.B(n_1285),
.Y(n_1831)
);

BUFx6f_ASAP7_75t_L g1832 ( 
.A(n_1354),
.Y(n_1832)
);

BUFx2_ASAP7_75t_L g1833 ( 
.A(n_1596),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1532),
.Y(n_1834)
);

INVx3_ASAP7_75t_L g1835 ( 
.A(n_1355),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1532),
.Y(n_1836)
);

NAND2xp33_ASAP7_75t_SL g1837 ( 
.A(n_1349),
.B(n_783),
.Y(n_1837)
);

BUFx6f_ASAP7_75t_L g1838 ( 
.A(n_1355),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1472),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1596),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_1581),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1504),
.B(n_1285),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1532),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1535),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1356),
.B(n_1369),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1535),
.Y(n_1846)
);

OAI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1369),
.A2(n_1127),
.B1(n_1134),
.B2(n_1132),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1535),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1535),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1472),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1553),
.Y(n_1851)
);

CKINVDCx6p67_ASAP7_75t_R g1852 ( 
.A(n_1591),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1567),
.B(n_1264),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1553),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1472),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1472),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1564),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1553),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1553),
.Y(n_1859)
);

BUFx6f_ASAP7_75t_L g1860 ( 
.A(n_1355),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1475),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1556),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1556),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1355),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1415),
.B(n_1197),
.Y(n_1865)
);

INVx3_ASAP7_75t_L g1866 ( 
.A(n_1409),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1475),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1475),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1475),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1556),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1480),
.Y(n_1871)
);

INVx3_ASAP7_75t_L g1872 ( 
.A(n_1409),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1480),
.Y(n_1873)
);

AND2x4_ASAP7_75t_SL g1874 ( 
.A(n_1564),
.B(n_969),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1480),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1372),
.B(n_1132),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1507),
.B(n_1286),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1480),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1556),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_1319),
.B(n_1134),
.Y(n_1880)
);

BUFx6f_ASAP7_75t_L g1881 ( 
.A(n_1409),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1562),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1409),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1447),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1562),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1447),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1447),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_R g1888 ( 
.A(n_1416),
.B(n_1138),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1562),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1447),
.Y(n_1890)
);

INVx3_ASAP7_75t_L g1891 ( 
.A(n_1412),
.Y(n_1891)
);

BUFx6f_ASAP7_75t_L g1892 ( 
.A(n_1412),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1379),
.B(n_1138),
.Y(n_1893)
);

BUFx3_ASAP7_75t_L g1894 ( 
.A(n_1449),
.Y(n_1894)
);

OAI21x1_ASAP7_75t_L g1895 ( 
.A1(n_1478),
.A2(n_1289),
.B(n_1288),
.Y(n_1895)
);

AND2x2_ASAP7_75t_SL g1896 ( 
.A(n_1524),
.B(n_1198),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1449),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1562),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1563),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1563),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1507),
.B(n_1288),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_1412),
.Y(n_1902)
);

BUFx8_ASAP7_75t_L g1903 ( 
.A(n_1295),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1521),
.B(n_1533),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1449),
.Y(n_1905)
);

OAI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1474),
.A2(n_1137),
.B(n_1168),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1563),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1563),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1552),
.B(n_1168),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1449),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1571),
.Y(n_1911)
);

INVx3_ASAP7_75t_L g1912 ( 
.A(n_1412),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1410),
.A2(n_974),
.B1(n_986),
.B2(n_969),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1521),
.B(n_1289),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1450),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1595),
.B(n_987),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1450),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1533),
.B(n_1294),
.Y(n_1918)
);

AND2x4_ASAP7_75t_L g1919 ( 
.A(n_1428),
.B(n_1200),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1450),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1450),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1571),
.Y(n_1922)
);

BUFx6f_ASAP7_75t_L g1923 ( 
.A(n_1418),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1571),
.Y(n_1924)
);

AND2x4_ASAP7_75t_L g1925 ( 
.A(n_1428),
.B(n_1204),
.Y(n_1925)
);

OA21x2_ASAP7_75t_L g1926 ( 
.A1(n_1569),
.A2(n_1582),
.B(n_1576),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1384),
.B(n_1465),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1465),
.B(n_1170),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1453),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1428),
.B(n_1422),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1571),
.Y(n_1931)
);

INVx3_ASAP7_75t_L g1932 ( 
.A(n_1418),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1453),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1453),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1453),
.Y(n_1935)
);

BUFx6f_ASAP7_75t_L g1936 ( 
.A(n_1418),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1592),
.B(n_1170),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1578),
.Y(n_1938)
);

INVx3_ASAP7_75t_L g1939 ( 
.A(n_1418),
.Y(n_1939)
);

NAND2xp33_ASAP7_75t_L g1940 ( 
.A(n_1486),
.B(n_1191),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1578),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1578),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1422),
.B(n_1206),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1485),
.B(n_1191),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1422),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1845),
.B(n_1927),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1640),
.B(n_1593),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1768),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1820),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1605),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1738),
.B(n_1584),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1820),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1808),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1605),
.Y(n_1954)
);

BUFx6f_ASAP7_75t_SL g1955 ( 
.A(n_1682),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1752),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1808),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1804),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1663),
.B(n_1321),
.Y(n_1959)
);

AND3x1_ASAP7_75t_L g1960 ( 
.A(n_1766),
.B(n_1368),
.C(n_1537),
.Y(n_1960)
);

INVx5_ASAP7_75t_L g1961 ( 
.A(n_1753),
.Y(n_1961)
);

INVx3_ASAP7_75t_L g1962 ( 
.A(n_1768),
.Y(n_1962)
);

AND2x2_ASAP7_75t_SL g1963 ( 
.A(n_1764),
.B(n_1519),
.Y(n_1963)
);

BUFx6f_ASAP7_75t_SL g1964 ( 
.A(n_1682),
.Y(n_1964)
);

INVx2_ASAP7_75t_SL g1965 ( 
.A(n_1812),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1759),
.B(n_1593),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1606),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1804),
.B(n_1593),
.Y(n_1968)
);

AOI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1764),
.A2(n_1520),
.B1(n_1545),
.B2(n_1519),
.Y(n_1969)
);

AND2x4_ASAP7_75t_L g1970 ( 
.A(n_1733),
.B(n_1469),
.Y(n_1970)
);

INVx2_ASAP7_75t_SL g1971 ( 
.A(n_1812),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1804),
.B(n_1469),
.Y(n_1972)
);

INVx3_ASAP7_75t_L g1973 ( 
.A(n_1768),
.Y(n_1973)
);

BUFx6f_ASAP7_75t_L g1974 ( 
.A(n_1753),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1606),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1603),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1608),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1610),
.B(n_1329),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1608),
.Y(n_1979)
);

NAND2xp33_ASAP7_75t_L g1980 ( 
.A(n_1753),
.B(n_1771),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_1753),
.Y(n_1981)
);

AOI22xp33_ASAP7_75t_L g1982 ( 
.A1(n_1753),
.A2(n_1486),
.B1(n_1434),
.B2(n_1442),
.Y(n_1982)
);

NAND2xp33_ASAP7_75t_L g1983 ( 
.A(n_1753),
.B(n_1486),
.Y(n_1983)
);

INVx2_ASAP7_75t_SL g1984 ( 
.A(n_1657),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_L g1985 ( 
.A(n_1794),
.B(n_1584),
.Y(n_1985)
);

AOI21x1_ASAP7_75t_L g1986 ( 
.A1(n_1674),
.A2(n_1509),
.B(n_1489),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1622),
.Y(n_1987)
);

BUFx6f_ASAP7_75t_L g1988 ( 
.A(n_1771),
.Y(n_1988)
);

OR2x2_ASAP7_75t_SL g1989 ( 
.A(n_1916),
.B(n_1500),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1622),
.Y(n_1990)
);

BUFx6f_ASAP7_75t_L g1991 ( 
.A(n_1771),
.Y(n_1991)
);

BUFx3_ASAP7_75t_L g1992 ( 
.A(n_1614),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1603),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1687),
.B(n_1469),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1623),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1604),
.Y(n_1996)
);

CKINVDCx20_ASAP7_75t_R g1997 ( 
.A(n_1913),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1694),
.B(n_1494),
.Y(n_1998)
);

INVx3_ASAP7_75t_L g1999 ( 
.A(n_1930),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1623),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1624),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_SL g2002 ( 
.A(n_1896),
.Y(n_2002)
);

BUFx6f_ASAP7_75t_L g2003 ( 
.A(n_1771),
.Y(n_2003)
);

CKINVDCx20_ASAP7_75t_R g2004 ( 
.A(n_1874),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1618),
.B(n_1411),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1604),
.Y(n_2006)
);

NAND3xp33_ASAP7_75t_L g2007 ( 
.A(n_1906),
.B(n_1442),
.C(n_1439),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1709),
.B(n_1494),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1684),
.B(n_1357),
.Y(n_2009)
);

INVx3_ASAP7_75t_L g2010 ( 
.A(n_1930),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1624),
.Y(n_2011)
);

INVx8_ASAP7_75t_L g2012 ( 
.A(n_1805),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1629),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1629),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_SL g2015 ( 
.A(n_1653),
.B(n_1405),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1683),
.B(n_1405),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1651),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1616),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_1697),
.B(n_1460),
.Y(n_2019)
);

BUFx6f_ASAP7_75t_L g2020 ( 
.A(n_1771),
.Y(n_2020)
);

CKINVDCx6p67_ASAP7_75t_R g2021 ( 
.A(n_1752),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1801),
.B(n_1494),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1651),
.Y(n_2023)
);

INVx4_ASAP7_75t_L g2024 ( 
.A(n_1771),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1659),
.Y(n_2025)
);

BUFx10_ASAP7_75t_L g2026 ( 
.A(n_1686),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1659),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1616),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1665),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1665),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1643),
.B(n_1460),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1801),
.B(n_1503),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1666),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1801),
.B(n_1503),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1666),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1667),
.Y(n_2036)
);

INVx1_ASAP7_75t_SL g2037 ( 
.A(n_1663),
.Y(n_2037)
);

INVx11_ASAP7_75t_L g2038 ( 
.A(n_1903),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1617),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1667),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_L g2041 ( 
.A(n_1847),
.B(n_1502),
.Y(n_2041)
);

CKINVDCx6p67_ASAP7_75t_R g2042 ( 
.A(n_1647),
.Y(n_2042)
);

BUFx10_ASAP7_75t_L g2043 ( 
.A(n_1699),
.Y(n_2043)
);

INVxp67_ASAP7_75t_SL g2044 ( 
.A(n_1894),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1690),
.Y(n_2045)
);

INVx2_ASAP7_75t_SL g2046 ( 
.A(n_1657),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1733),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1904),
.Y(n_2048)
);

INVx2_ASAP7_75t_SL g2049 ( 
.A(n_1732),
.Y(n_2049)
);

BUFx8_ASAP7_75t_SL g2050 ( 
.A(n_1647),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1904),
.Y(n_2051)
);

HB1xp67_ASAP7_75t_L g2052 ( 
.A(n_1602),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_1819),
.B(n_1502),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1626),
.B(n_1503),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1819),
.B(n_1511),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1690),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1700),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1626),
.B(n_1508),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1930),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1700),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1701),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1613),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1615),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1627),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1618),
.B(n_1523),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1632),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_1909),
.B(n_1511),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1701),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1708),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1708),
.Y(n_2070)
);

BUFx6f_ASAP7_75t_L g2071 ( 
.A(n_1635),
.Y(n_2071)
);

AND2x6_ASAP7_75t_L g2072 ( 
.A(n_1678),
.B(n_1364),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1636),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1711),
.Y(n_2074)
);

AND3x2_ASAP7_75t_L g2075 ( 
.A(n_1725),
.B(n_1458),
.C(n_1424),
.Y(n_2075)
);

BUFx6f_ASAP7_75t_L g2076 ( 
.A(n_1635),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1711),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1716),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1637),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1728),
.B(n_1508),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1638),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1716),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_1717),
.Y(n_2083)
);

NOR2xp33_ASAP7_75t_L g2084 ( 
.A(n_1937),
.B(n_1514),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_L g2085 ( 
.A(n_1944),
.B(n_1514),
.Y(n_2085)
);

OR2x2_ASAP7_75t_SL g2086 ( 
.A(n_1916),
.B(n_1499),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1717),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1654),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1721),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1721),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1734),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1656),
.Y(n_2092)
);

INVx3_ASAP7_75t_L g2093 ( 
.A(n_1734),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1746),
.Y(n_2094)
);

BUFx6f_ASAP7_75t_L g2095 ( 
.A(n_1635),
.Y(n_2095)
);

INVx3_ASAP7_75t_L g2096 ( 
.A(n_1746),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1617),
.Y(n_2097)
);

INVx3_ASAP7_75t_L g2098 ( 
.A(n_1749),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1749),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1779),
.B(n_1719),
.Y(n_2100)
);

BUFx2_ASAP7_75t_L g2101 ( 
.A(n_1602),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1756),
.B(n_1508),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1635),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1750),
.Y(n_2104)
);

BUFx3_ASAP7_75t_L g2105 ( 
.A(n_1614),
.Y(n_2105)
);

INVx2_ASAP7_75t_SL g2106 ( 
.A(n_1732),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1661),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1750),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_L g2109 ( 
.A(n_1635),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_1758),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1758),
.Y(n_2111)
);

INVxp67_ASAP7_75t_SL g2112 ( 
.A(n_1894),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1763),
.Y(n_2113)
);

NAND2xp33_ASAP7_75t_L g2114 ( 
.A(n_1805),
.B(n_1486),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1763),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1769),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1769),
.Y(n_2117)
);

OR2x6_ASAP7_75t_L g2118 ( 
.A(n_1833),
.B(n_1599),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1772),
.Y(n_2119)
);

NOR2xp33_ASAP7_75t_L g2120 ( 
.A(n_1876),
.B(n_1416),
.Y(n_2120)
);

INVx3_ASAP7_75t_L g2121 ( 
.A(n_1772),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_1619),
.B(n_1528),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_L g2123 ( 
.A(n_1893),
.B(n_1555),
.Y(n_2123)
);

INVx3_ASAP7_75t_L g2124 ( 
.A(n_1774),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1609),
.B(n_1512),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1774),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1775),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1775),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1751),
.Y(n_2129)
);

INVx2_ASAP7_75t_SL g2130 ( 
.A(n_1732),
.Y(n_2130)
);

BUFx2_ASAP7_75t_L g2131 ( 
.A(n_1630),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1782),
.Y(n_2132)
);

CKINVDCx5p33_ASAP7_75t_R g2133 ( 
.A(n_1693),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1751),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_L g2135 ( 
.A(n_1928),
.B(n_1555),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1782),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_SL g2137 ( 
.A(n_1833),
.B(n_1513),
.Y(n_2137)
);

BUFx6f_ASAP7_75t_SL g2138 ( 
.A(n_1896),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1786),
.Y(n_2139)
);

NAND3xp33_ASAP7_75t_L g2140 ( 
.A(n_1940),
.B(n_1448),
.C(n_1439),
.Y(n_2140)
);

CKINVDCx6p67_ASAP7_75t_R g2141 ( 
.A(n_1852),
.Y(n_2141)
);

BUFx3_ASAP7_75t_L g2142 ( 
.A(n_1625),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1628),
.B(n_1512),
.Y(n_2143)
);

INVxp67_ASAP7_75t_SL g2144 ( 
.A(n_1799),
.Y(n_2144)
);

INVxp33_ASAP7_75t_SL g2145 ( 
.A(n_1888),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1786),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_SL g2147 ( 
.A(n_1840),
.B(n_1516),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_1619),
.B(n_1531),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_SL g2149 ( 
.A(n_1840),
.B(n_1600),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1945),
.Y(n_2150)
);

INVxp33_ASAP7_75t_SL g2151 ( 
.A(n_1696),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_1639),
.B(n_1668),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1945),
.Y(n_2153)
);

CKINVDCx20_ASAP7_75t_R g2154 ( 
.A(n_1874),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1918),
.Y(n_2155)
);

NOR2x1p5_ASAP7_75t_L g2156 ( 
.A(n_1852),
.B(n_1295),
.Y(n_2156)
);

BUFx10_ASAP7_75t_L g2157 ( 
.A(n_1791),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1918),
.Y(n_2158)
);

INVxp67_ASAP7_75t_SL g2159 ( 
.A(n_1799),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1787),
.Y(n_2160)
);

AOI21x1_ASAP7_75t_L g2161 ( 
.A1(n_1674),
.A2(n_1544),
.B(n_1515),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1620),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1787),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1620),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1795),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1645),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_1639),
.B(n_1534),
.Y(n_2167)
);

INVx4_ASAP7_75t_L g2168 ( 
.A(n_1612),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1795),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1645),
.Y(n_2170)
);

INVx3_ASAP7_75t_L g2171 ( 
.A(n_1800),
.Y(n_2171)
);

CKINVDCx5p33_ASAP7_75t_R g2172 ( 
.A(n_1693),
.Y(n_2172)
);

INVx3_ASAP7_75t_L g2173 ( 
.A(n_1800),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1649),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1649),
.Y(n_2175)
);

INVx3_ASAP7_75t_L g2176 ( 
.A(n_1802),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1660),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1660),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1744),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1689),
.Y(n_2180)
);

OAI22xp33_ASAP7_75t_SL g2181 ( 
.A1(n_1789),
.A2(n_1464),
.B1(n_1448),
.B2(n_1434),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1689),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1691),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1744),
.Y(n_2184)
);

BUFx6f_ASAP7_75t_SL g2185 ( 
.A(n_1625),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1792),
.B(n_1520),
.Y(n_2186)
);

OAI22xp33_ASAP7_75t_L g2187 ( 
.A1(n_1796),
.A2(n_1785),
.B1(n_1783),
.B2(n_1781),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1744),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1842),
.Y(n_2189)
);

NAND2xp33_ASAP7_75t_L g2190 ( 
.A(n_1805),
.B(n_1596),
.Y(n_2190)
);

BUFx3_ASAP7_75t_L g2191 ( 
.A(n_1648),
.Y(n_2191)
);

BUFx6f_ASAP7_75t_L g2192 ( 
.A(n_1672),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_1740),
.B(n_1545),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1691),
.Y(n_2194)
);

BUFx6f_ASAP7_75t_L g2195 ( 
.A(n_1672),
.Y(n_2195)
);

BUFx6f_ASAP7_75t_L g2196 ( 
.A(n_1672),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1692),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1842),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1877),
.Y(n_2199)
);

BUFx2_ASAP7_75t_L g2200 ( 
.A(n_1630),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1692),
.Y(n_2201)
);

BUFx10_ASAP7_75t_L g2202 ( 
.A(n_1702),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1695),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1695),
.Y(n_2204)
);

BUFx6f_ASAP7_75t_L g2205 ( 
.A(n_1672),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1703),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1703),
.Y(n_2207)
);

INVx2_ASAP7_75t_SL g2208 ( 
.A(n_1736),
.Y(n_2208)
);

AO21x2_ASAP7_75t_L g2209 ( 
.A1(n_1895),
.A2(n_1550),
.B(n_1431),
.Y(n_2209)
);

NAND2xp33_ASAP7_75t_L g2210 ( 
.A(n_1805),
.B(n_1596),
.Y(n_2210)
);

NOR2xp33_ASAP7_75t_L g2211 ( 
.A(n_1853),
.B(n_1570),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_1877),
.Y(n_2212)
);

NOR2x1p5_ASAP7_75t_L g2213 ( 
.A(n_1853),
.B(n_1312),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1705),
.Y(n_2214)
);

INVxp33_ASAP7_75t_L g2215 ( 
.A(n_1601),
.Y(n_2215)
);

BUFx6f_ASAP7_75t_L g2216 ( 
.A(n_1672),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1705),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_1641),
.B(n_1642),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_SL g2219 ( 
.A(n_1740),
.B(n_1736),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1706),
.Y(n_2220)
);

NAND3xp33_ASAP7_75t_L g2221 ( 
.A(n_1940),
.B(n_1492),
.C(n_1481),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1901),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1901),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1914),
.Y(n_2224)
);

INVx2_ASAP7_75t_SL g2225 ( 
.A(n_1736),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_1669),
.B(n_1512),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1706),
.Y(n_2227)
);

INVx3_ASAP7_75t_L g2228 ( 
.A(n_1802),
.Y(n_2228)
);

NAND3xp33_ASAP7_75t_L g2229 ( 
.A(n_1837),
.B(n_1492),
.C(n_1481),
.Y(n_2229)
);

BUFx10_ASAP7_75t_L g2230 ( 
.A(n_1702),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1707),
.Y(n_2231)
);

INVx3_ASAP7_75t_L g2232 ( 
.A(n_1803),
.Y(n_2232)
);

INVx2_ASAP7_75t_SL g2233 ( 
.A(n_1740),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1914),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1760),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_1662),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_SL g2237 ( 
.A(n_1607),
.B(n_1573),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_1670),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_1679),
.B(n_1527),
.Y(n_2239)
);

INVx3_ASAP7_75t_L g2240 ( 
.A(n_1803),
.Y(n_2240)
);

OAI22xp5_ASAP7_75t_SL g2241 ( 
.A1(n_1652),
.A2(n_974),
.B1(n_1049),
.B2(n_986),
.Y(n_2241)
);

NOR2xp33_ASAP7_75t_L g2242 ( 
.A(n_1677),
.B(n_1570),
.Y(n_2242)
);

INVxp67_ASAP7_75t_SL g2243 ( 
.A(n_1807),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_1676),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1761),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1680),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1707),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1710),
.Y(n_2248)
);

AO22x2_ASAP7_75t_L g2249 ( 
.A1(n_1607),
.A2(n_1370),
.B1(n_660),
.B2(n_711),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1710),
.Y(n_2250)
);

BUFx3_ASAP7_75t_L g2251 ( 
.A(n_1648),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1714),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_1926),
.B(n_1527),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1681),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1714),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1720),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1720),
.Y(n_2257)
);

BUFx4f_ASAP7_75t_L g2258 ( 
.A(n_1805),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1777),
.Y(n_2259)
);

NOR2x1p5_ASAP7_75t_L g2260 ( 
.A(n_1841),
.B(n_1312),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1926),
.B(n_1527),
.Y(n_2261)
);

INVx4_ASAP7_75t_L g2262 ( 
.A(n_1612),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1807),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_1815),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1815),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_SL g2266 ( 
.A(n_1607),
.B(n_1573),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1816),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1919),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1919),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_SL g2270 ( 
.A(n_1631),
.B(n_1590),
.Y(n_2270)
);

OR2x2_ASAP7_75t_L g2271 ( 
.A(n_1634),
.B(n_1421),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1919),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1816),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_1631),
.B(n_1590),
.Y(n_2274)
);

INVx3_ASAP7_75t_L g2275 ( 
.A(n_1825),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1925),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1825),
.Y(n_2277)
);

INVx3_ASAP7_75t_L g2278 ( 
.A(n_1839),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_1631),
.B(n_1391),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1839),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_1850),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1797),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1925),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_1850),
.Y(n_2284)
);

CKINVDCx5p33_ASAP7_75t_R g2285 ( 
.A(n_1841),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1797),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_SL g2287 ( 
.A(n_1650),
.B(n_1664),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1797),
.Y(n_2288)
);

AOI22xp33_ASAP7_75t_L g2289 ( 
.A1(n_1818),
.A2(n_1529),
.B1(n_1542),
.B2(n_1540),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1818),
.Y(n_2290)
);

INVxp67_ASAP7_75t_L g2291 ( 
.A(n_1790),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_1855),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_SL g2293 ( 
.A(n_1650),
.B(n_1561),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_1855),
.Y(n_2294)
);

NAND3xp33_ASAP7_75t_L g2295 ( 
.A(n_1837),
.B(n_1549),
.C(n_1538),
.Y(n_2295)
);

BUFx6f_ASAP7_75t_SL g2296 ( 
.A(n_1655),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_1650),
.B(n_1565),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1925),
.Y(n_2298)
);

INVx8_ASAP7_75t_L g2299 ( 
.A(n_1805),
.Y(n_2299)
);

OR2x2_ASAP7_75t_L g2300 ( 
.A(n_1634),
.B(n_1430),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1818),
.Y(n_2301)
);

NOR2xp67_ASAP7_75t_L g2302 ( 
.A(n_2229),
.B(n_1599),
.Y(n_2302)
);

OR2x2_ASAP7_75t_L g2303 ( 
.A(n_2037),
.B(n_1646),
.Y(n_2303)
);

INVx2_ASAP7_75t_SL g2304 ( 
.A(n_2101),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2150),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_1946),
.B(n_2100),
.Y(n_2306)
);

NOR2xp33_ASAP7_75t_L g2307 ( 
.A(n_1951),
.B(n_1985),
.Y(n_2307)
);

AND2x6_ASAP7_75t_L g2308 ( 
.A(n_1948),
.B(n_1644),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2153),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_SL g2310 ( 
.A(n_1965),
.B(n_1675),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1958),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1976),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_1976),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1993),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1993),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1996),
.Y(n_2316)
);

INVx1_ASAP7_75t_SL g2317 ( 
.A(n_2101),
.Y(n_2317)
);

INVxp67_ASAP7_75t_L g2318 ( 
.A(n_2052),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1996),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2006),
.Y(n_2320)
);

NAND2x1p5_ASAP7_75t_L g2321 ( 
.A(n_2024),
.B(n_1655),
.Y(n_2321)
);

BUFx6f_ASAP7_75t_L g2322 ( 
.A(n_1992),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_L g2323 ( 
.A(n_2186),
.B(n_1790),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_L g2324 ( 
.A(n_2007),
.B(n_1788),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2006),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2018),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2018),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2005),
.B(n_1677),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2028),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2259),
.B(n_1926),
.Y(n_2330)
);

CKINVDCx5p33_ASAP7_75t_R g2331 ( 
.A(n_2145),
.Y(n_2331)
);

XNOR2x1_ASAP7_75t_L g2332 ( 
.A(n_1960),
.B(n_1559),
.Y(n_2332)
);

CKINVDCx20_ASAP7_75t_R g2333 ( 
.A(n_2050),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2028),
.Y(n_2334)
);

NAND2x1p5_ASAP7_75t_L g2335 ( 
.A(n_2024),
.B(n_1865),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2039),
.Y(n_2336)
);

INVx2_ASAP7_75t_SL g2337 ( 
.A(n_2131),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2259),
.B(n_1718),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2039),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_1950),
.Y(n_2340)
);

INVxp33_ASAP7_75t_L g2341 ( 
.A(n_1959),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2097),
.Y(n_2342)
);

OAI21xp5_ASAP7_75t_L g2343 ( 
.A1(n_1948),
.A2(n_1895),
.B(n_1831),
.Y(n_2343)
);

BUFx6f_ASAP7_75t_L g2344 ( 
.A(n_1992),
.Y(n_2344)
);

CKINVDCx16_ASAP7_75t_R g2345 ( 
.A(n_2202),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2097),
.Y(n_2346)
);

AND2x6_ASAP7_75t_L g2347 ( 
.A(n_1974),
.B(n_1668),
.Y(n_2347)
);

INVxp67_ASAP7_75t_L g2348 ( 
.A(n_2131),
.Y(n_2348)
);

AND2x2_ASAP7_75t_SL g2349 ( 
.A(n_1963),
.B(n_1498),
.Y(n_2349)
);

INVx1_ASAP7_75t_SL g2350 ( 
.A(n_2200),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2162),
.Y(n_2351)
);

XOR2xp5_ASAP7_75t_L g2352 ( 
.A(n_2241),
.B(n_1049),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2162),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_SL g2354 ( 
.A(n_1965),
.B(n_1664),
.Y(n_2354)
);

HB1xp67_ASAP7_75t_L g2355 ( 
.A(n_2200),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2005),
.B(n_1726),
.Y(n_2356)
);

XOR2xp5_ASAP7_75t_L g2357 ( 
.A(n_2145),
.B(n_1074),
.Y(n_2357)
);

INVxp33_ASAP7_75t_L g2358 ( 
.A(n_1959),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2164),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2164),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_1950),
.Y(n_2361)
);

CKINVDCx16_ASAP7_75t_R g2362 ( 
.A(n_2202),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2166),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2065),
.B(n_1726),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_L g2365 ( 
.A(n_2120),
.B(n_1074),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2166),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2175),
.Y(n_2367)
);

AND2x6_ASAP7_75t_L g2368 ( 
.A(n_1974),
.B(n_1704),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2175),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_2065),
.B(n_2122),
.Y(n_2370)
);

CKINVDCx5p33_ASAP7_75t_R g2371 ( 
.A(n_2050),
.Y(n_2371)
);

CKINVDCx20_ASAP7_75t_R g2372 ( 
.A(n_2042),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2122),
.B(n_1829),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2047),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2059),
.Y(n_2375)
);

INVxp33_ASAP7_75t_L g2376 ( 
.A(n_2211),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2170),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2170),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2174),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2174),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2177),
.Y(n_2381)
);

NAND2x1p5_ASAP7_75t_L g2382 ( 
.A(n_2024),
.B(n_1865),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2177),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2178),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2178),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_2148),
.B(n_1857),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_2148),
.B(n_1538),
.Y(n_2387)
);

AND2x4_ASAP7_75t_L g2388 ( 
.A(n_2105),
.B(n_1745),
.Y(n_2388)
);

OAI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_2179),
.A2(n_1831),
.B(n_1730),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_1971),
.B(n_1549),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2189),
.Y(n_2391)
);

CKINVDCx20_ASAP7_75t_R g2392 ( 
.A(n_2042),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2189),
.Y(n_2393)
);

CKINVDCx20_ASAP7_75t_R g2394 ( 
.A(n_2004),
.Y(n_2394)
);

NAND2xp33_ASAP7_75t_SL g2395 ( 
.A(n_2002),
.B(n_1712),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_1969),
.B(n_1577),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2198),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2198),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2199),
.Y(n_2399)
);

AND2x2_ASAP7_75t_L g2400 ( 
.A(n_1971),
.B(n_1577),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2199),
.Y(n_2401)
);

BUFx6f_ASAP7_75t_L g2402 ( 
.A(n_2105),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_1984),
.B(n_1543),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2212),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_1984),
.B(n_1586),
.Y(n_2405)
);

OR2x2_ASAP7_75t_L g2406 ( 
.A(n_2271),
.B(n_1880),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_2123),
.B(n_1747),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2218),
.B(n_1718),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2212),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2222),
.Y(n_2410)
);

NAND2x1p5_ASAP7_75t_L g2411 ( 
.A(n_1974),
.B(n_1981),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2222),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2223),
.Y(n_2413)
);

INVx1_ASAP7_75t_SL g2414 ( 
.A(n_2271),
.Y(n_2414)
);

NOR2xp67_ASAP7_75t_L g2415 ( 
.A(n_2295),
.B(n_1328),
.Y(n_2415)
);

XOR2xp5_ASAP7_75t_L g2416 ( 
.A(n_2133),
.B(n_1106),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2223),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2224),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2224),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_1999),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_1999),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_1954),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_1999),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2046),
.B(n_1704),
.Y(n_2424)
);

AND2x4_ASAP7_75t_L g2425 ( 
.A(n_2142),
.B(n_1754),
.Y(n_2425)
);

XNOR2x2_ASAP7_75t_L g2426 ( 
.A(n_2140),
.B(n_690),
.Y(n_2426)
);

OR2x2_ASAP7_75t_L g2427 ( 
.A(n_2300),
.B(n_1611),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2187),
.B(n_1730),
.Y(n_2428)
);

CKINVDCx16_ASAP7_75t_R g2429 ( 
.A(n_2202),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2010),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2010),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2010),
.Y(n_2432)
);

XNOR2xp5_ASAP7_75t_L g2433 ( 
.A(n_2151),
.B(n_1106),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2282),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2282),
.Y(n_2435)
);

OR2x6_ASAP7_75t_L g2436 ( 
.A(n_2118),
.B(n_1377),
.Y(n_2436)
);

NOR2xp33_ASAP7_75t_L g2437 ( 
.A(n_2067),
.B(n_1119),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2286),
.Y(n_2438)
);

XOR2xp5_ASAP7_75t_L g2439 ( 
.A(n_2133),
.B(n_1119),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2286),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2288),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2102),
.B(n_1664),
.Y(n_2442)
);

AOI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2253),
.A2(n_1612),
.B(n_1688),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2046),
.B(n_1432),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2288),
.Y(n_2445)
);

XNOR2x2_ASAP7_75t_L g2446 ( 
.A(n_2135),
.B(n_716),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2290),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_2172),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2152),
.B(n_1436),
.Y(n_2449)
);

XOR2xp5_ASAP7_75t_L g2450 ( 
.A(n_2172),
.B(n_1216),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2290),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2301),
.Y(n_2452)
);

CKINVDCx5p33_ASAP7_75t_R g2453 ( 
.A(n_2285),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2301),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2180),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2180),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2182),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2182),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_1954),
.Y(n_2459)
);

CKINVDCx20_ASAP7_75t_R g2460 ( 
.A(n_2004),
.Y(n_2460)
);

BUFx6f_ASAP7_75t_L g2461 ( 
.A(n_2142),
.Y(n_2461)
);

AND2x2_ASAP7_75t_L g2462 ( 
.A(n_2152),
.B(n_1456),
.Y(n_2462)
);

NOR2xp33_ASAP7_75t_L g2463 ( 
.A(n_1963),
.B(n_1755),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2183),
.Y(n_2464)
);

XOR2x2_ASAP7_75t_L g2465 ( 
.A(n_2151),
.B(n_1722),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2183),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2194),
.Y(n_2467)
);

CKINVDCx20_ASAP7_75t_R g2468 ( 
.A(n_2154),
.Y(n_2468)
);

AND2x4_ASAP7_75t_L g2469 ( 
.A(n_2191),
.B(n_1698),
.Y(n_2469)
);

CKINVDCx20_ASAP7_75t_R g2470 ( 
.A(n_2154),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2194),
.Y(n_2471)
);

AOI21xp5_ASAP7_75t_L g2472 ( 
.A1(n_2261),
.A2(n_1727),
.B(n_1724),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2197),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2197),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2167),
.B(n_1406),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2201),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2201),
.Y(n_2477)
);

INVx4_ASAP7_75t_SL g2478 ( 
.A(n_1974),
.Y(n_2478)
);

AND2x4_ASAP7_75t_L g2479 ( 
.A(n_2191),
.B(n_1698),
.Y(n_2479)
);

NOR2xp33_ASAP7_75t_L g2480 ( 
.A(n_2084),
.B(n_1216),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2203),
.Y(n_2481)
);

HB1xp67_ASAP7_75t_L g2482 ( 
.A(n_2300),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2203),
.Y(n_2483)
);

XOR2xp5_ASAP7_75t_L g2484 ( 
.A(n_2285),
.B(n_1287),
.Y(n_2484)
);

XNOR2x2_ASAP7_75t_L g2485 ( 
.A(n_2221),
.B(n_1464),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2204),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2204),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2206),
.Y(n_2488)
);

INVx1_ASAP7_75t_SL g2489 ( 
.A(n_2167),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2206),
.Y(n_2490)
);

AND2x4_ASAP7_75t_L g2491 ( 
.A(n_2251),
.B(n_1698),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2207),
.Y(n_2492)
);

INVxp33_ASAP7_75t_L g2493 ( 
.A(n_2215),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2207),
.Y(n_2494)
);

INVx2_ASAP7_75t_SL g2495 ( 
.A(n_2235),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2214),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2214),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2217),
.Y(n_2498)
);

OAI21xp5_ASAP7_75t_L g2499 ( 
.A1(n_2179),
.A2(n_1865),
.B(n_1713),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_SL g2500 ( 
.A(n_2080),
.B(n_1713),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2217),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2220),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_1967),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2220),
.Y(n_2504)
);

NOR2xp33_ASAP7_75t_L g2505 ( 
.A(n_1966),
.B(n_1192),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2227),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2227),
.Y(n_2507)
);

AND2x4_ASAP7_75t_L g2508 ( 
.A(n_2251),
.B(n_1713),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2231),
.Y(n_2509)
);

NOR2xp33_ASAP7_75t_L g2510 ( 
.A(n_2085),
.B(n_1287),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2231),
.Y(n_2511)
);

BUFx3_ASAP7_75t_L g2512 ( 
.A(n_2230),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_1967),
.Y(n_2513)
);

NAND2xp33_ASAP7_75t_R g2514 ( 
.A(n_2075),
.B(n_1327),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2252),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2252),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2257),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2257),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2242),
.B(n_1473),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_L g2520 ( 
.A(n_2009),
.B(n_1291),
.Y(n_2520)
);

AND2x2_ASAP7_75t_L g2521 ( 
.A(n_2155),
.B(n_1296),
.Y(n_2521)
);

BUFx6f_ASAP7_75t_SL g2522 ( 
.A(n_2230),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_SL g2523 ( 
.A(n_2181),
.B(n_1943),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2048),
.Y(n_2524)
);

XOR2xp5_ASAP7_75t_L g2525 ( 
.A(n_1956),
.B(n_1291),
.Y(n_2525)
);

OAI21xp5_ASAP7_75t_L g2526 ( 
.A1(n_2184),
.A2(n_1943),
.B(n_1739),
.Y(n_2526)
);

INVxp67_ASAP7_75t_L g2527 ( 
.A(n_2054),
.Y(n_2527)
);

NOR2xp33_ASAP7_75t_L g2528 ( 
.A(n_2026),
.B(n_1327),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2051),
.Y(n_2529)
);

INVx1_ASAP7_75t_SL g2530 ( 
.A(n_2193),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2247),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2158),
.B(n_1301),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2248),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2234),
.B(n_1192),
.Y(n_2534)
);

NOR2xp33_ASAP7_75t_L g2535 ( 
.A(n_2026),
.B(n_1377),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_1947),
.B(n_1943),
.Y(n_2536)
);

OAI21xp5_ASAP7_75t_L g2537 ( 
.A1(n_2184),
.A2(n_1741),
.B(n_1737),
.Y(n_2537)
);

AOI21xp5_ASAP7_75t_L g2538 ( 
.A1(n_2022),
.A2(n_1742),
.B(n_1856),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2250),
.Y(n_2539)
);

BUFx3_ASAP7_75t_L g2540 ( 
.A(n_2230),
.Y(n_2540)
);

NAND2x1p5_ASAP7_75t_L g2541 ( 
.A(n_1974),
.B(n_1843),
.Y(n_2541)
);

NAND2xp33_ASAP7_75t_SL g2542 ( 
.A(n_2002),
.B(n_831),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2255),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2256),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_1975),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_1975),
.Y(n_2546)
);

CKINVDCx20_ASAP7_75t_R g2547 ( 
.A(n_2021),
.Y(n_2547)
);

INVxp67_ASAP7_75t_SL g2548 ( 
.A(n_2071),
.Y(n_2548)
);

OR2x6_ASAP7_75t_L g2549 ( 
.A(n_2118),
.B(n_1387),
.Y(n_2549)
);

NOR2xp33_ASAP7_75t_L g2550 ( 
.A(n_2026),
.B(n_1387),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_1977),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2032),
.B(n_1843),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2129),
.B(n_1199),
.Y(n_2553)
);

AND2x2_ASAP7_75t_L g2554 ( 
.A(n_2134),
.B(n_1199),
.Y(n_2554)
);

BUFx2_ASAP7_75t_SL g2555 ( 
.A(n_2185),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_1977),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_1979),
.Y(n_2557)
);

INVxp33_ASAP7_75t_SL g2558 ( 
.A(n_1956),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_1979),
.Y(n_2559)
);

XOR2xp5_ASAP7_75t_L g2560 ( 
.A(n_1997),
.B(n_1581),
.Y(n_2560)
);

INVxp33_ASAP7_75t_L g2561 ( 
.A(n_2237),
.Y(n_2561)
);

NOR2xp33_ASAP7_75t_SL g2562 ( 
.A(n_2002),
.B(n_1715),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_1987),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_1987),
.Y(n_2564)
);

NOR2xp33_ASAP7_75t_L g2565 ( 
.A(n_2043),
.B(n_1978),
.Y(n_2565)
);

OR2x6_ASAP7_75t_L g2566 ( 
.A(n_2118),
.B(n_1401),
.Y(n_2566)
);

INVx2_ASAP7_75t_SL g2567 ( 
.A(n_2245),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_1990),
.Y(n_2568)
);

AND2x6_ASAP7_75t_L g2569 ( 
.A(n_1981),
.B(n_1856),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_1990),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_1995),
.Y(n_2571)
);

INVx2_ASAP7_75t_SL g2572 ( 
.A(n_2062),
.Y(n_2572)
);

NOR2xp33_ASAP7_75t_L g2573 ( 
.A(n_2043),
.B(n_1401),
.Y(n_2573)
);

OR2x6_ASAP7_75t_L g2574 ( 
.A(n_2118),
.B(n_1407),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_1995),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2000),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_1953),
.B(n_1202),
.Y(n_2577)
);

NOR2xp67_ASAP7_75t_L g2578 ( 
.A(n_2291),
.B(n_1328),
.Y(n_2578)
);

XOR2xp5_ASAP7_75t_L g2579 ( 
.A(n_1997),
.B(n_1594),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2000),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_L g2581 ( 
.A(n_2043),
.B(n_1407),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2001),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2001),
.Y(n_2583)
);

AND2x4_ASAP7_75t_L g2584 ( 
.A(n_2233),
.B(n_1529),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2011),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2011),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2034),
.B(n_1844),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2013),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2013),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_1957),
.B(n_1202),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2014),
.Y(n_2591)
);

XNOR2xp5_ASAP7_75t_L g2592 ( 
.A(n_2213),
.B(n_1594),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_1994),
.B(n_1205),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_L g2594 ( 
.A(n_2015),
.B(n_1490),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2014),
.Y(n_2595)
);

INVxp67_ASAP7_75t_SL g2596 ( 
.A(n_2071),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2017),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2017),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2023),
.Y(n_2599)
);

XOR2xp5_ASAP7_75t_L g2600 ( 
.A(n_2266),
.B(n_1205),
.Y(n_2600)
);

INVxp67_ASAP7_75t_L g2601 ( 
.A(n_2058),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2023),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2025),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2025),
.Y(n_2604)
);

INVxp33_ASAP7_75t_L g2605 ( 
.A(n_2270),
.Y(n_2605)
);

HB1xp67_ASAP7_75t_L g2606 ( 
.A(n_2268),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2027),
.Y(n_2607)
);

CKINVDCx20_ASAP7_75t_R g2608 ( 
.A(n_2021),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2027),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2029),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2029),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2030),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2030),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2033),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2033),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_1998),
.B(n_1844),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2035),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2035),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2036),
.Y(n_2619)
);

NOR2xp33_ASAP7_75t_L g2620 ( 
.A(n_2016),
.B(n_1490),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2036),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2040),
.Y(n_2622)
);

AND2x2_ASAP7_75t_L g2623 ( 
.A(n_2008),
.B(n_1221),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_SL g2624 ( 
.A(n_2233),
.B(n_1426),
.Y(n_2624)
);

INVx2_ASAP7_75t_SL g2625 ( 
.A(n_2063),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2040),
.Y(n_2626)
);

INVxp67_ASAP7_75t_L g2627 ( 
.A(n_2125),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2143),
.B(n_1846),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2045),
.Y(n_2629)
);

AND2x2_ASAP7_75t_L g2630 ( 
.A(n_2279),
.B(n_1221),
.Y(n_2630)
);

AND2x6_ASAP7_75t_L g2631 ( 
.A(n_1981),
.B(n_1861),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2045),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2056),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2056),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_SL g2635 ( 
.A(n_1982),
.B(n_1462),
.Y(n_2635)
);

XOR2x2_ASAP7_75t_L g2636 ( 
.A(n_2041),
.B(n_1378),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2049),
.B(n_1222),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2057),
.Y(n_2638)
);

NOR2xp67_ASAP7_75t_L g2639 ( 
.A(n_2049),
.B(n_1338),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2057),
.Y(n_2640)
);

INVxp67_ASAP7_75t_SL g2641 ( 
.A(n_2071),
.Y(n_2641)
);

NOR2xp33_ASAP7_75t_L g2642 ( 
.A(n_2019),
.B(n_1574),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_1962),
.B(n_1846),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2060),
.Y(n_2644)
);

NOR2xp33_ASAP7_75t_L g2645 ( 
.A(n_2149),
.B(n_1574),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2060),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2061),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2312),
.Y(n_2648)
);

NOR2xp33_ASAP7_75t_SL g2649 ( 
.A(n_2448),
.B(n_1715),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2313),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2314),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2340),
.Y(n_2652)
);

NOR2xp33_ASAP7_75t_L g2653 ( 
.A(n_2307),
.B(n_2138),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2315),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_SL g2655 ( 
.A(n_2387),
.B(n_2106),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2306),
.B(n_2226),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2361),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_SL g2658 ( 
.A(n_2489),
.B(n_2106),
.Y(n_2658)
);

NOR2x1p5_ASAP7_75t_L g2659 ( 
.A(n_2371),
.B(n_2141),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2316),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2422),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2306),
.B(n_2239),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2408),
.B(n_1962),
.Y(n_2663)
);

AOI22xp5_ASAP7_75t_L g2664 ( 
.A1(n_2396),
.A2(n_1964),
.B1(n_1955),
.B2(n_2138),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2319),
.Y(n_2665)
);

NOR2xp33_ASAP7_75t_L g2666 ( 
.A(n_2376),
.B(n_2138),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_SL g2667 ( 
.A(n_2489),
.B(n_2130),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2408),
.B(n_1962),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2320),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2325),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2373),
.B(n_2274),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2326),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_SL g2673 ( 
.A(n_2407),
.B(n_2130),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2327),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2459),
.Y(n_2675)
);

NOR2xp33_ASAP7_75t_L g2676 ( 
.A(n_2505),
.B(n_1955),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2329),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2334),
.Y(n_2678)
);

HB1xp67_ASAP7_75t_L g2679 ( 
.A(n_2355),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_SL g2680 ( 
.A(n_2407),
.B(n_2208),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2627),
.B(n_1973),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2627),
.B(n_1973),
.Y(n_2682)
);

INVx8_ASAP7_75t_L g2683 ( 
.A(n_2347),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2370),
.B(n_2527),
.Y(n_2684)
);

BUFx5_ASAP7_75t_L g2685 ( 
.A(n_2569),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2336),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2339),
.Y(n_2687)
);

OAI22xp33_ASAP7_75t_L g2688 ( 
.A1(n_2396),
.A2(n_2208),
.B1(n_2225),
.B2(n_2269),
.Y(n_2688)
);

INVx2_ASAP7_75t_SL g2689 ( 
.A(n_2355),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2527),
.B(n_1970),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_SL g2691 ( 
.A(n_2349),
.B(n_2225),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2601),
.B(n_2505),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2601),
.B(n_1970),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_L g2694 ( 
.A(n_2437),
.B(n_1955),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2519),
.B(n_1970),
.Y(n_2695)
);

AOI22xp5_ASAP7_75t_L g2696 ( 
.A1(n_2323),
.A2(n_1964),
.B1(n_2623),
.B2(n_2593),
.Y(n_2696)
);

AO22x1_ASAP7_75t_L g2697 ( 
.A1(n_2365),
.A2(n_1397),
.B1(n_1496),
.B2(n_1420),
.Y(n_2697)
);

NOR2xp67_ASAP7_75t_SL g2698 ( 
.A(n_2555),
.B(n_1961),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_SL g2699 ( 
.A(n_2405),
.B(n_2289),
.Y(n_2699)
);

INVxp67_ASAP7_75t_L g2700 ( 
.A(n_2482),
.Y(n_2700)
);

O2A1O1Ixp5_ASAP7_75t_L g2701 ( 
.A1(n_2635),
.A2(n_2053),
.B(n_2055),
.C(n_1986),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2475),
.B(n_2072),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2442),
.B(n_2072),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2442),
.B(n_2072),
.Y(n_2704)
);

NOR2xp33_ASAP7_75t_L g2705 ( 
.A(n_2480),
.B(n_1964),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2390),
.B(n_2072),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2400),
.B(n_2072),
.Y(n_2707)
);

AOI22xp33_ASAP7_75t_L g2708 ( 
.A1(n_2323),
.A2(n_2272),
.B1(n_2283),
.B2(n_2276),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_SL g2709 ( 
.A(n_2530),
.B(n_1961),
.Y(n_2709)
);

AOI22xp5_ASAP7_75t_L g2710 ( 
.A1(n_2510),
.A2(n_2530),
.B1(n_2630),
.B2(n_2463),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2338),
.B(n_2072),
.Y(n_2711)
);

BUFx3_ASAP7_75t_L g2712 ( 
.A(n_2304),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2338),
.B(n_2064),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2449),
.B(n_2066),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2342),
.Y(n_2715)
);

NOR2xp67_ASAP7_75t_L g2716 ( 
.A(n_2453),
.B(n_2031),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2462),
.B(n_2073),
.Y(n_2717)
);

BUFx3_ASAP7_75t_L g2718 ( 
.A(n_2337),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2346),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2536),
.B(n_2079),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2536),
.B(n_2081),
.Y(n_2721)
);

AOI22xp33_ASAP7_75t_L g2722 ( 
.A1(n_2463),
.A2(n_2298),
.B1(n_1952),
.B2(n_1949),
.Y(n_2722)
);

INVxp67_ASAP7_75t_L g2723 ( 
.A(n_2482),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2364),
.B(n_2088),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_SL g2725 ( 
.A(n_2328),
.B(n_2356),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2351),
.Y(n_2726)
);

BUFx6f_ASAP7_75t_SL g2727 ( 
.A(n_2512),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2353),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_SL g2729 ( 
.A(n_2444),
.B(n_1961),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_SL g2730 ( 
.A(n_2403),
.B(n_2469),
.Y(n_2730)
);

INVx2_ASAP7_75t_SL g2731 ( 
.A(n_2317),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2455),
.B(n_2092),
.Y(n_2732)
);

NOR2x1_ASAP7_75t_L g2733 ( 
.A(n_2639),
.B(n_2156),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2503),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2359),
.Y(n_2735)
);

NOR2xp33_ASAP7_75t_L g2736 ( 
.A(n_2341),
.B(n_2137),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2360),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_SL g2738 ( 
.A(n_2469),
.B(n_1961),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2616),
.B(n_1973),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2616),
.B(n_1968),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2428),
.B(n_1972),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2428),
.B(n_2188),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2456),
.B(n_2188),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2457),
.B(n_2236),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2513),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2363),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2366),
.Y(n_2747)
);

NOR2xp67_ASAP7_75t_SL g2748 ( 
.A(n_2345),
.B(n_1961),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2551),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2458),
.B(n_2236),
.Y(n_2750)
);

NOR2xp33_ASAP7_75t_L g2751 ( 
.A(n_2358),
.B(n_2520),
.Y(n_2751)
);

A2O1A1Ixp33_ASAP7_75t_L g2752 ( 
.A1(n_2324),
.A2(n_2523),
.B(n_2565),
.C(n_2466),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2367),
.Y(n_2753)
);

INVx8_ASAP7_75t_L g2754 ( 
.A(n_2347),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2564),
.Y(n_2755)
);

O2A1O1Ixp5_ASAP7_75t_L g2756 ( 
.A1(n_2310),
.A2(n_2161),
.B(n_1986),
.C(n_2147),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2613),
.Y(n_2757)
);

NOR2xp33_ASAP7_75t_L g2758 ( 
.A(n_2414),
.B(n_2293),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_SL g2759 ( 
.A(n_2479),
.B(n_2508),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2369),
.Y(n_2760)
);

INVx3_ASAP7_75t_L g2761 ( 
.A(n_2411),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2464),
.B(n_2238),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2467),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2614),
.Y(n_2764)
);

AND2x6_ASAP7_75t_SL g2765 ( 
.A(n_2535),
.B(n_1903),
.Y(n_2765)
);

NOR2xp33_ASAP7_75t_L g2766 ( 
.A(n_2414),
.B(n_2297),
.Y(n_2766)
);

AND2x4_ASAP7_75t_L g2767 ( 
.A(n_2479),
.B(n_2287),
.Y(n_2767)
);

INVx2_ASAP7_75t_SL g2768 ( 
.A(n_2317),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_2638),
.Y(n_2769)
);

INVxp67_ASAP7_75t_L g2770 ( 
.A(n_2303),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2471),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2473),
.B(n_2107),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2377),
.Y(n_2773)
);

INVxp67_ASAP7_75t_L g2774 ( 
.A(n_2350),
.Y(n_2774)
);

AO22x1_ASAP7_75t_L g2775 ( 
.A1(n_2528),
.A2(n_1397),
.B1(n_1496),
.B2(n_1420),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2386),
.B(n_2249),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2474),
.B(n_2249),
.Y(n_2777)
);

INVxp67_ASAP7_75t_L g2778 ( 
.A(n_2350),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_SL g2779 ( 
.A(n_2491),
.B(n_2168),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_SL g2780 ( 
.A(n_2491),
.B(n_2168),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2378),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2534),
.B(n_2249),
.Y(n_2782)
);

INVx2_ASAP7_75t_SL g2783 ( 
.A(n_2427),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2476),
.B(n_2249),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2477),
.Y(n_2785)
);

NOR2xp33_ASAP7_75t_L g2786 ( 
.A(n_2348),
.B(n_1499),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2379),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_SL g2788 ( 
.A(n_2508),
.B(n_2424),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2481),
.B(n_2238),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2380),
.Y(n_2790)
);

INVxp67_ASAP7_75t_L g2791 ( 
.A(n_2406),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2381),
.Y(n_2792)
);

OAI22xp5_ASAP7_75t_L g2793 ( 
.A1(n_2483),
.A2(n_2258),
.B1(n_2086),
.B2(n_2219),
.Y(n_2793)
);

NOR2xp33_ASAP7_75t_L g2794 ( 
.A(n_2348),
.B(n_1499),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_SL g2795 ( 
.A(n_2572),
.B(n_2168),
.Y(n_2795)
);

AND2x4_ASAP7_75t_L g2796 ( 
.A(n_2388),
.B(n_2044),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2383),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2384),
.Y(n_2798)
);

INVx3_ASAP7_75t_L g2799 ( 
.A(n_2411),
.Y(n_2799)
);

NOR2xp33_ASAP7_75t_L g2800 ( 
.A(n_2318),
.B(n_2086),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2486),
.B(n_2244),
.Y(n_2801)
);

BUFx6f_ASAP7_75t_L g2802 ( 
.A(n_2322),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2487),
.B(n_2244),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2488),
.B(n_2246),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2490),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2492),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2494),
.B(n_2246),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2496),
.Y(n_2808)
);

HB1xp67_ASAP7_75t_L g2809 ( 
.A(n_2318),
.Y(n_2809)
);

NAND3xp33_ASAP7_75t_L g2810 ( 
.A(n_2324),
.B(n_1230),
.C(n_1222),
.Y(n_2810)
);

NOR2xp33_ASAP7_75t_L g2811 ( 
.A(n_2493),
.B(n_1989),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2497),
.B(n_2254),
.Y(n_2812)
);

NAND2xp33_ASAP7_75t_L g2813 ( 
.A(n_2347),
.B(n_1981),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2385),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_SL g2815 ( 
.A(n_2625),
.B(n_2262),
.Y(n_2815)
);

AOI22xp33_ASAP7_75t_L g2816 ( 
.A1(n_2426),
.A2(n_2254),
.B1(n_2210),
.B2(n_2190),
.Y(n_2816)
);

NOR2xp33_ASAP7_75t_L g2817 ( 
.A(n_2561),
.B(n_1989),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2498),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2545),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2501),
.B(n_2112),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2502),
.Y(n_2821)
);

INVx3_ASAP7_75t_L g2822 ( 
.A(n_2335),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_SL g2823 ( 
.A(n_2322),
.B(n_2262),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2504),
.B(n_2262),
.Y(n_2824)
);

NOR2xp33_ASAP7_75t_L g2825 ( 
.A(n_2605),
.B(n_1230),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2506),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2507),
.B(n_2061),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2509),
.B(n_2511),
.Y(n_2828)
);

AND2x2_ASAP7_75t_L g2829 ( 
.A(n_2577),
.B(n_1261),
.Y(n_2829)
);

OAI22xp33_ASAP7_75t_L g2830 ( 
.A1(n_2562),
.A2(n_2141),
.B1(n_1476),
.B2(n_2258),
.Y(n_2830)
);

OR2x6_ASAP7_75t_SL g2831 ( 
.A(n_2331),
.B(n_1261),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_L g2832 ( 
.A(n_2332),
.B(n_1265),
.Y(n_2832)
);

AND2x6_ASAP7_75t_SL g2833 ( 
.A(n_2550),
.B(n_1903),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2515),
.B(n_2516),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2517),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_SL g2836 ( 
.A(n_2322),
.B(n_2258),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2518),
.B(n_2068),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2552),
.B(n_2068),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2546),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2434),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_SL g2841 ( 
.A(n_2344),
.B(n_2020),
.Y(n_2841)
);

OR2x6_ASAP7_75t_L g2842 ( 
.A(n_2436),
.B(n_2260),
.Y(n_2842)
);

NAND3xp33_ASAP7_75t_L g2843 ( 
.A(n_2433),
.B(n_1278),
.C(n_1265),
.Y(n_2843)
);

CKINVDCx11_ASAP7_75t_R g2844 ( 
.A(n_2333),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2552),
.B(n_2069),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2556),
.Y(n_2846)
);

INVxp67_ASAP7_75t_L g2847 ( 
.A(n_2553),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2587),
.B(n_2069),
.Y(n_2848)
);

BUFx6f_ASAP7_75t_L g2849 ( 
.A(n_2344),
.Y(n_2849)
);

INVx1_ASAP7_75t_SL g2850 ( 
.A(n_2554),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2435),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2438),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_SL g2853 ( 
.A(n_2344),
.B(n_2402),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2587),
.B(n_2070),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2557),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2440),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2628),
.B(n_2070),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2628),
.B(n_2074),
.Y(n_2858)
);

INVx2_ASAP7_75t_SL g2859 ( 
.A(n_2388),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2391),
.B(n_2074),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2393),
.B(n_2077),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2441),
.Y(n_2862)
);

OR2x2_ASAP7_75t_L g2863 ( 
.A(n_2357),
.B(n_1278),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2445),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2559),
.Y(n_2865)
);

AND2x6_ASAP7_75t_SL g2866 ( 
.A(n_2573),
.B(n_2038),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2447),
.Y(n_2867)
);

BUFx5_ASAP7_75t_L g2868 ( 
.A(n_2569),
.Y(n_2868)
);

AND2x2_ASAP7_75t_L g2869 ( 
.A(n_2590),
.B(n_1031),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_2397),
.B(n_2077),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2563),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2451),
.Y(n_2872)
);

AOI22xp33_ASAP7_75t_L g2873 ( 
.A1(n_2446),
.A2(n_2210),
.B1(n_2190),
.B2(n_1540),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2452),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2398),
.B(n_2078),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2568),
.Y(n_2876)
);

NAND2x1p5_ASAP7_75t_L g2877 ( 
.A(n_2402),
.B(n_1981),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2454),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_SL g2879 ( 
.A(n_2402),
.B(n_1988),
.Y(n_2879)
);

AND2x4_ASAP7_75t_SL g2880 ( 
.A(n_2461),
.B(n_2157),
.Y(n_2880)
);

AOI21xp5_ASAP7_75t_L g2881 ( 
.A1(n_2499),
.A2(n_1980),
.B(n_2299),
.Y(n_2881)
);

A2O1A1Ixp33_ASAP7_75t_L g2882 ( 
.A1(n_2500),
.A2(n_2114),
.B(n_1983),
.C(n_1980),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2399),
.B(n_2078),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2401),
.B(n_2082),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_SL g2885 ( 
.A(n_2461),
.B(n_1991),
.Y(n_2885)
);

AOI22xp5_ASAP7_75t_L g2886 ( 
.A1(n_2395),
.A2(n_2114),
.B1(n_2296),
.B2(n_2185),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_SL g2887 ( 
.A(n_2461),
.B(n_1991),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2404),
.B(n_2082),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2409),
.B(n_2083),
.Y(n_2889)
);

INVx2_ASAP7_75t_SL g2890 ( 
.A(n_2425),
.Y(n_2890)
);

O2A1O1Ixp33_ASAP7_75t_L g2891 ( 
.A1(n_2620),
.A2(n_1402),
.B(n_1983),
.C(n_1540),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2410),
.B(n_2083),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2531),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2412),
.B(n_2087),
.Y(n_2894)
);

AOI22xp33_ASAP7_75t_L g2895 ( 
.A1(n_2485),
.A2(n_1529),
.B1(n_1542),
.B2(n_2185),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2413),
.B(n_2087),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2570),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2417),
.B(n_2089),
.Y(n_2898)
);

INVx2_ASAP7_75t_L g2899 ( 
.A(n_2571),
.Y(n_2899)
);

NOR2x1_ASAP7_75t_L g2900 ( 
.A(n_2578),
.B(n_2171),
.Y(n_2900)
);

AND2x2_ASAP7_75t_L g2901 ( 
.A(n_2637),
.B(n_1058),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2418),
.B(n_2089),
.Y(n_2902)
);

BUFx6f_ASAP7_75t_L g2903 ( 
.A(n_2347),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_SL g2904 ( 
.A(n_2584),
.B(n_1988),
.Y(n_2904)
);

NOR2xp33_ASAP7_75t_L g2905 ( 
.A(n_2600),
.B(n_1338),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_SL g2906 ( 
.A(n_2584),
.B(n_1988),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2533),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2575),
.Y(n_2908)
);

BUFx6f_ASAP7_75t_L g2909 ( 
.A(n_2368),
.Y(n_2909)
);

AND2x2_ASAP7_75t_L g2910 ( 
.A(n_2521),
.B(n_1073),
.Y(n_2910)
);

OAI22xp5_ASAP7_75t_L g2911 ( 
.A1(n_2330),
.A2(n_2419),
.B1(n_2543),
.B2(n_2539),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2330),
.B(n_2090),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_L g2913 ( 
.A(n_2594),
.B(n_2495),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2544),
.B(n_2090),
.Y(n_2914)
);

AOI22xp33_ASAP7_75t_L g2915 ( 
.A1(n_2311),
.A2(n_1542),
.B1(n_2296),
.B2(n_1991),
.Y(n_2915)
);

OR2x6_ASAP7_75t_L g2916 ( 
.A(n_2436),
.B(n_2299),
.Y(n_2916)
);

NOR2xp33_ASAP7_75t_L g2917 ( 
.A(n_2567),
.B(n_1351),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_SL g2918 ( 
.A(n_2562),
.B(n_1991),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2576),
.Y(n_2919)
);

NOR2xp33_ASAP7_75t_L g2920 ( 
.A(n_2642),
.B(n_2581),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2499),
.A2(n_2299),
.B(n_2012),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_SL g2922 ( 
.A(n_2302),
.B(n_1991),
.Y(n_2922)
);

NAND2xp33_ASAP7_75t_SL g2923 ( 
.A(n_2522),
.B(n_2296),
.Y(n_2923)
);

INVxp67_ASAP7_75t_L g2924 ( 
.A(n_2532),
.Y(n_2924)
);

NOR2x1_ASAP7_75t_L g2925 ( 
.A(n_2540),
.B(n_2171),
.Y(n_2925)
);

AOI22xp33_ASAP7_75t_L g2926 ( 
.A1(n_2375),
.A2(n_2368),
.B1(n_2374),
.B2(n_2308),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2524),
.B(n_2091),
.Y(n_2927)
);

INVx2_ASAP7_75t_L g2928 ( 
.A(n_2580),
.Y(n_2928)
);

AND2x4_ASAP7_75t_L g2929 ( 
.A(n_2425),
.B(n_1988),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_2582),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2583),
.Y(n_2931)
);

HB1xp67_ASAP7_75t_L g2932 ( 
.A(n_2606),
.Y(n_2932)
);

AND2x2_ASAP7_75t_L g2933 ( 
.A(n_2606),
.B(n_1117),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_SL g2934 ( 
.A(n_2415),
.B(n_1988),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_SL g2935 ( 
.A(n_2645),
.B(n_2020),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2692),
.B(n_2529),
.Y(n_2936)
);

AND2x2_ASAP7_75t_L g2937 ( 
.A(n_2671),
.B(n_2465),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2656),
.B(n_2354),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2656),
.B(n_2309),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2662),
.B(n_2305),
.Y(n_2940)
);

AOI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2740),
.A2(n_2881),
.B(n_2299),
.Y(n_2941)
);

BUFx6f_ASAP7_75t_L g2942 ( 
.A(n_2802),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2662),
.B(n_2368),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2720),
.B(n_2368),
.Y(n_2944)
);

BUFx2_ASAP7_75t_L g2945 ( 
.A(n_2731),
.Y(n_2945)
);

NOR2xp33_ASAP7_75t_SL g2946 ( 
.A(n_2649),
.B(n_2558),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2893),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_SL g2948 ( 
.A(n_2751),
.B(n_2542),
.Y(n_2948)
);

AOI21xp5_ASAP7_75t_L g2949 ( 
.A1(n_2740),
.A2(n_2012),
.B(n_2921),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_SL g2950 ( 
.A(n_2710),
.B(n_2362),
.Y(n_2950)
);

AOI21xp5_ASAP7_75t_L g2951 ( 
.A1(n_2741),
.A2(n_2012),
.B(n_2548),
.Y(n_2951)
);

AO21x1_ASAP7_75t_L g2952 ( 
.A1(n_2911),
.A2(n_2443),
.B(n_2538),
.Y(n_2952)
);

NOR2x2_ASAP7_75t_L g2953 ( 
.A(n_2842),
.B(n_2436),
.Y(n_2953)
);

OAI22xp5_ASAP7_75t_L g2954 ( 
.A1(n_2713),
.A2(n_2548),
.B1(n_2641),
.B2(n_2596),
.Y(n_2954)
);

AOI21xp5_ASAP7_75t_L g2955 ( 
.A1(n_2741),
.A2(n_2012),
.B(n_2596),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2684),
.B(n_2308),
.Y(n_2956)
);

OAI21xp5_ASAP7_75t_L g2957 ( 
.A1(n_2752),
.A2(n_2538),
.B(n_2472),
.Y(n_2957)
);

OAI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_2701),
.A2(n_2472),
.B(n_2389),
.Y(n_2958)
);

INVx2_ASAP7_75t_L g2959 ( 
.A(n_2819),
.Y(n_2959)
);

AOI21xp5_ASAP7_75t_L g2960 ( 
.A1(n_2882),
.A2(n_2813),
.B(n_2838),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2684),
.B(n_2308),
.Y(n_2961)
);

OAI21xp5_ASAP7_75t_L g2962 ( 
.A1(n_2695),
.A2(n_2389),
.B(n_2526),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2839),
.Y(n_2963)
);

AOI21xp5_ASAP7_75t_L g2964 ( 
.A1(n_2838),
.A2(n_2848),
.B(n_2845),
.Y(n_2964)
);

AOI21xp5_ASAP7_75t_L g2965 ( 
.A1(n_2845),
.A2(n_2641),
.B(n_2526),
.Y(n_2965)
);

OAI22xp5_ASAP7_75t_L g2966 ( 
.A1(n_2834),
.A2(n_2321),
.B1(n_2382),
.B2(n_2335),
.Y(n_2966)
);

BUFx6f_ASAP7_75t_L g2967 ( 
.A(n_2802),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_SL g2968 ( 
.A(n_2850),
.B(n_2768),
.Y(n_2968)
);

AOI21x1_ASAP7_75t_L g2969 ( 
.A1(n_2703),
.A2(n_2443),
.B(n_2343),
.Y(n_2969)
);

INVx3_ASAP7_75t_L g2970 ( 
.A(n_2683),
.Y(n_2970)
);

AOI21x1_ASAP7_75t_L g2971 ( 
.A1(n_2704),
.A2(n_2343),
.B(n_2161),
.Y(n_2971)
);

BUFx2_ASAP7_75t_L g2972 ( 
.A(n_2774),
.Y(n_2972)
);

OAI21xp5_ASAP7_75t_L g2973 ( 
.A1(n_2756),
.A2(n_2537),
.B(n_2421),
.Y(n_2973)
);

INVx2_ASAP7_75t_SL g2974 ( 
.A(n_2712),
.Y(n_2974)
);

OAI21xp5_ASAP7_75t_L g2975 ( 
.A1(n_2711),
.A2(n_2537),
.B(n_2423),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2846),
.Y(n_2976)
);

AND2x4_ASAP7_75t_L g2977 ( 
.A(n_2796),
.B(n_2478),
.Y(n_2977)
);

AOI21xp5_ASAP7_75t_L g2978 ( 
.A1(n_2848),
.A2(n_2624),
.B(n_2076),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2721),
.B(n_2308),
.Y(n_2979)
);

OAI22xp5_ASAP7_75t_L g2980 ( 
.A1(n_2834),
.A2(n_2321),
.B1(n_2382),
.B2(n_2420),
.Y(n_2980)
);

NOR2xp67_ASAP7_75t_L g2981 ( 
.A(n_2917),
.B(n_1351),
.Y(n_2981)
);

NOR2xp33_ASAP7_75t_L g2982 ( 
.A(n_2920),
.B(n_2416),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2724),
.B(n_2430),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2653),
.B(n_2431),
.Y(n_2984)
);

AOI21xp5_ASAP7_75t_L g2985 ( 
.A1(n_2854),
.A2(n_2076),
.B(n_2071),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2676),
.B(n_2432),
.Y(n_2986)
);

OAI21xp5_ASAP7_75t_L g2987 ( 
.A1(n_2706),
.A2(n_2643),
.B(n_2586),
.Y(n_2987)
);

AOI21xp5_ASAP7_75t_L g2988 ( 
.A1(n_2854),
.A2(n_2076),
.B(n_2071),
.Y(n_2988)
);

AOI33xp33_ASAP7_75t_L g2989 ( 
.A1(n_2869),
.A2(n_1212),
.A3(n_1207),
.B1(n_1217),
.B2(n_1215),
.B3(n_1211),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_SL g2990 ( 
.A(n_2913),
.B(n_2429),
.Y(n_2990)
);

AOI21xp5_ASAP7_75t_L g2991 ( 
.A1(n_2739),
.A2(n_2095),
.B(n_2076),
.Y(n_2991)
);

NOR2xp33_ASAP7_75t_L g2992 ( 
.A(n_2832),
.B(n_2439),
.Y(n_2992)
);

INVxp67_ASAP7_75t_L g2993 ( 
.A(n_2679),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_SL g2994 ( 
.A(n_2778),
.B(n_2636),
.Y(n_2994)
);

AOI22xp5_ASAP7_75t_L g2995 ( 
.A1(n_2694),
.A2(n_2352),
.B1(n_2514),
.B2(n_2484),
.Y(n_2995)
);

O2A1O1Ixp33_ASAP7_75t_L g2996 ( 
.A1(n_2847),
.A2(n_2691),
.B(n_2699),
.C(n_2791),
.Y(n_2996)
);

AND2x4_ASAP7_75t_L g2997 ( 
.A(n_2796),
.B(n_2478),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2714),
.B(n_2643),
.Y(n_2998)
);

OAI21xp5_ASAP7_75t_L g2999 ( 
.A1(n_2707),
.A2(n_2588),
.B(n_2585),
.Y(n_2999)
);

NOR2xp33_ASAP7_75t_L g3000 ( 
.A(n_2705),
.B(n_2450),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2717),
.B(n_2589),
.Y(n_3001)
);

AOI21xp5_ASAP7_75t_L g3002 ( 
.A1(n_2739),
.A2(n_2095),
.B(n_2076),
.Y(n_3002)
);

A2O1A1Ixp33_ASAP7_75t_L g3003 ( 
.A1(n_2891),
.A2(n_2618),
.B(n_2619),
.C(n_2617),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_SL g3004 ( 
.A(n_2825),
.B(n_1378),
.Y(n_3004)
);

AOI21xp5_ASAP7_75t_L g3005 ( 
.A1(n_2857),
.A2(n_2103),
.B(n_2095),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_SL g3006 ( 
.A(n_2783),
.B(n_1378),
.Y(n_3006)
);

A2O1A1Ixp33_ASAP7_75t_L g3007 ( 
.A1(n_2696),
.A2(n_2626),
.B(n_2629),
.C(n_2622),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_SL g3008 ( 
.A(n_2829),
.B(n_2157),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2907),
.Y(n_3009)
);

OAI21xp5_ASAP7_75t_L g3010 ( 
.A1(n_2702),
.A2(n_2595),
.B(n_2591),
.Y(n_3010)
);

OAI21xp5_ASAP7_75t_L g3011 ( 
.A1(n_2673),
.A2(n_2598),
.B(n_2597),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2855),
.Y(n_3012)
);

NOR2x1_ASAP7_75t_L g3013 ( 
.A(n_2718),
.B(n_2394),
.Y(n_3013)
);

OR2x6_ASAP7_75t_L g3014 ( 
.A(n_2683),
.B(n_2754),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_SL g3015 ( 
.A(n_2758),
.B(n_2157),
.Y(n_3015)
);

INVx1_ASAP7_75t_SL g3016 ( 
.A(n_2809),
.Y(n_3016)
);

AND2x4_ASAP7_75t_L g3017 ( 
.A(n_2929),
.B(n_2478),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2725),
.B(n_2599),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2690),
.B(n_2602),
.Y(n_3019)
);

INVx2_ASAP7_75t_SL g3020 ( 
.A(n_2880),
.Y(n_3020)
);

AOI22xp33_ASAP7_75t_L g3021 ( 
.A1(n_2776),
.A2(n_2566),
.B1(n_2574),
.B2(n_2549),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2648),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2865),
.Y(n_3023)
);

OAI21xp5_ASAP7_75t_L g3024 ( 
.A1(n_2680),
.A2(n_2604),
.B(n_2603),
.Y(n_3024)
);

OAI22xp5_ASAP7_75t_L g3025 ( 
.A1(n_2828),
.A2(n_2541),
.B1(n_2609),
.B2(n_2607),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_SL g3026 ( 
.A(n_2766),
.B(n_2003),
.Y(n_3026)
);

INVx1_ASAP7_75t_SL g3027 ( 
.A(n_2689),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2871),
.Y(n_3028)
);

AOI21xp5_ASAP7_75t_L g3029 ( 
.A1(n_2857),
.A2(n_2103),
.B(n_2095),
.Y(n_3029)
);

AOI21xp5_ASAP7_75t_L g3030 ( 
.A1(n_2858),
.A2(n_2668),
.B(n_2663),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2693),
.B(n_2610),
.Y(n_3031)
);

A2O1A1Ixp33_ASAP7_75t_L g3032 ( 
.A1(n_2810),
.A2(n_2621),
.B(n_2632),
.C(n_2615),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2782),
.B(n_2611),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_2901),
.B(n_2612),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2650),
.Y(n_3035)
);

CKINVDCx10_ASAP7_75t_R g3036 ( 
.A(n_2727),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_SL g3037 ( 
.A(n_2736),
.B(n_2003),
.Y(n_3037)
);

AOI21xp5_ASAP7_75t_L g3038 ( 
.A1(n_2858),
.A2(n_2103),
.B(n_2095),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2732),
.B(n_2633),
.Y(n_3039)
);

AOI21xp5_ASAP7_75t_L g3040 ( 
.A1(n_2663),
.A2(n_2109),
.B(n_2103),
.Y(n_3040)
);

AOI21xp5_ASAP7_75t_L g3041 ( 
.A1(n_2668),
.A2(n_2109),
.B(n_2103),
.Y(n_3041)
);

NOR2xp67_ASAP7_75t_L g3042 ( 
.A(n_2770),
.B(n_1373),
.Y(n_3042)
);

NOR2xp33_ASAP7_75t_L g3043 ( 
.A(n_2843),
.B(n_2525),
.Y(n_3043)
);

OAI21xp5_ASAP7_75t_L g3044 ( 
.A1(n_2824),
.A2(n_2640),
.B(n_2634),
.Y(n_3044)
);

AOI21xp5_ASAP7_75t_L g3045 ( 
.A1(n_2742),
.A2(n_2192),
.B(n_2109),
.Y(n_3045)
);

OAI21xp5_ASAP7_75t_L g3046 ( 
.A1(n_2742),
.A2(n_2646),
.B(n_2644),
.Y(n_3046)
);

NOR2x1_ASAP7_75t_L g3047 ( 
.A(n_2733),
.B(n_2460),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2772),
.B(n_2647),
.Y(n_3048)
);

INVx3_ASAP7_75t_L g3049 ( 
.A(n_2683),
.Y(n_3049)
);

AOI21xp5_ASAP7_75t_L g3050 ( 
.A1(n_2912),
.A2(n_2192),
.B(n_2109),
.Y(n_3050)
);

AOI21xp5_ASAP7_75t_L g3051 ( 
.A1(n_2912),
.A2(n_2192),
.B(n_2109),
.Y(n_3051)
);

AOI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_2935),
.A2(n_2195),
.B(n_2192),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2924),
.B(n_2091),
.Y(n_3053)
);

AND2x4_ASAP7_75t_L g3054 ( 
.A(n_2929),
.B(n_2549),
.Y(n_3054)
);

OAI21xp5_ASAP7_75t_L g3055 ( 
.A1(n_2911),
.A2(n_2655),
.B(n_2816),
.Y(n_3055)
);

AOI21xp5_ASAP7_75t_L g3056 ( 
.A1(n_2793),
.A2(n_2195),
.B(n_2192),
.Y(n_3056)
);

AOI22xp33_ASAP7_75t_L g3057 ( 
.A1(n_2817),
.A2(n_2566),
.B1(n_2574),
.B2(n_2549),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_2910),
.B(n_2094),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2651),
.Y(n_3059)
);

A2O1A1Ixp33_ASAP7_75t_L g3060 ( 
.A1(n_2873),
.A2(n_2094),
.B(n_2104),
.C(n_2099),
.Y(n_3060)
);

INVx3_ASAP7_75t_L g3061 ( 
.A(n_2754),
.Y(n_3061)
);

AOI21xp5_ASAP7_75t_L g3062 ( 
.A1(n_2793),
.A2(n_2196),
.B(n_2195),
.Y(n_3062)
);

HB1xp67_ASAP7_75t_L g3063 ( 
.A(n_2700),
.Y(n_3063)
);

AOI21xp5_ASAP7_75t_L g3064 ( 
.A1(n_2918),
.A2(n_2196),
.B(n_2195),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2933),
.B(n_2099),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2767),
.B(n_2104),
.Y(n_3066)
);

AOI21xp5_ASAP7_75t_L g3067 ( 
.A1(n_2836),
.A2(n_2196),
.B(n_2195),
.Y(n_3067)
);

HB1xp67_ASAP7_75t_L g3068 ( 
.A(n_2723),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2767),
.B(n_2108),
.Y(n_3069)
);

AOI21xp5_ASAP7_75t_L g3070 ( 
.A1(n_2681),
.A2(n_2205),
.B(n_2196),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2654),
.B(n_2108),
.Y(n_3071)
);

HB1xp67_ASAP7_75t_L g3072 ( 
.A(n_2932),
.Y(n_3072)
);

O2A1O1Ixp33_ASAP7_75t_L g3073 ( 
.A1(n_2688),
.A2(n_1124),
.B(n_1560),
.C(n_1497),
.Y(n_3073)
);

AOI21xp5_ASAP7_75t_L g3074 ( 
.A1(n_2681),
.A2(n_2205),
.B(n_2196),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_2876),
.Y(n_3075)
);

AOI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_2682),
.A2(n_2216),
.B(n_2205),
.Y(n_3076)
);

HB1xp67_ASAP7_75t_L g3077 ( 
.A(n_2802),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2660),
.B(n_2111),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2897),
.Y(n_3079)
);

CKINVDCx10_ASAP7_75t_R g3080 ( 
.A(n_2727),
.Y(n_3080)
);

INVx1_ASAP7_75t_SL g3081 ( 
.A(n_2863),
.Y(n_3081)
);

AOI21xp5_ASAP7_75t_L g3082 ( 
.A1(n_2682),
.A2(n_2216),
.B(n_2205),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2665),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_SL g3084 ( 
.A(n_2716),
.B(n_2003),
.Y(n_3084)
);

AO21x1_ASAP7_75t_L g3085 ( 
.A1(n_2777),
.A2(n_2541),
.B(n_1849),
.Y(n_3085)
);

AND2x2_ASAP7_75t_L g3086 ( 
.A(n_2666),
.B(n_1025),
.Y(n_3086)
);

BUFx4f_ASAP7_75t_L g3087 ( 
.A(n_2903),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_SL g3088 ( 
.A(n_2800),
.B(n_2003),
.Y(n_3088)
);

OAI21xp5_ASAP7_75t_L g3089 ( 
.A1(n_2784),
.A2(n_2159),
.B(n_2144),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2669),
.B(n_2111),
.Y(n_3090)
);

AOI21xp5_ASAP7_75t_L g3091 ( 
.A1(n_2779),
.A2(n_2216),
.B(n_2205),
.Y(n_3091)
);

OAI21xp5_ASAP7_75t_L g3092 ( 
.A1(n_2729),
.A2(n_2243),
.B(n_2263),
.Y(n_3092)
);

AOI21xp5_ASAP7_75t_L g3093 ( 
.A1(n_2780),
.A2(n_2216),
.B(n_2020),
.Y(n_3093)
);

AOI21xp5_ASAP7_75t_L g3094 ( 
.A1(n_2904),
.A2(n_2216),
.B(n_2020),
.Y(n_3094)
);

O2A1O1Ixp33_ASAP7_75t_L g3095 ( 
.A1(n_2730),
.A2(n_1497),
.B(n_1530),
.C(n_1487),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_2744),
.B(n_2750),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2670),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2672),
.Y(n_3098)
);

INVxp33_ASAP7_75t_L g3099 ( 
.A(n_2811),
.Y(n_3099)
);

AOI21xp5_ASAP7_75t_L g3100 ( 
.A1(n_2906),
.A2(n_2020),
.B(n_2003),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_2744),
.B(n_2113),
.Y(n_3101)
);

CKINVDCx5p33_ASAP7_75t_R g3102 ( 
.A(n_2844),
.Y(n_3102)
);

AOI21x1_ASAP7_75t_L g3103 ( 
.A1(n_2795),
.A2(n_2264),
.B(n_2263),
.Y(n_3103)
);

AOI21xp5_ASAP7_75t_L g3104 ( 
.A1(n_2743),
.A2(n_2209),
.B(n_2264),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2750),
.B(n_2113),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2762),
.B(n_2115),
.Y(n_3106)
);

NOR2xp67_ASAP7_75t_L g3107 ( 
.A(n_2859),
.B(n_1373),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2762),
.B(n_2115),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2789),
.B(n_2116),
.Y(n_3109)
);

AOI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_2743),
.A2(n_2209),
.B(n_2265),
.Y(n_3110)
);

OAI21xp5_ASAP7_75t_L g3111 ( 
.A1(n_2708),
.A2(n_2267),
.B(n_2265),
.Y(n_3111)
);

NOR2xp33_ASAP7_75t_L g3112 ( 
.A(n_2788),
.B(n_2468),
.Y(n_3112)
);

AOI21xp5_ASAP7_75t_L g3113 ( 
.A1(n_2922),
.A2(n_2209),
.B(n_2267),
.Y(n_3113)
);

INVx4_ASAP7_75t_L g3114 ( 
.A(n_2754),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2674),
.Y(n_3115)
);

AND2x2_ASAP7_75t_L g3116 ( 
.A(n_2890),
.B(n_1065),
.Y(n_3116)
);

AOI21xp5_ASAP7_75t_L g3117 ( 
.A1(n_2934),
.A2(n_2277),
.B(n_2273),
.Y(n_3117)
);

AOI21xp5_ASAP7_75t_L g3118 ( 
.A1(n_2815),
.A2(n_2277),
.B(n_2273),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_2899),
.Y(n_3119)
);

NOR2xp33_ASAP7_75t_L g3120 ( 
.A(n_2905),
.B(n_2470),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2908),
.Y(n_3121)
);

AOI21xp5_ASAP7_75t_L g3122 ( 
.A1(n_2789),
.A2(n_2281),
.B(n_2280),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_SL g3123 ( 
.A(n_2664),
.B(n_2849),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2801),
.B(n_2116),
.Y(n_3124)
);

NOR2xp67_ASAP7_75t_L g3125 ( 
.A(n_2786),
.B(n_1374),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2677),
.Y(n_3126)
);

A2O1A1Ixp33_ASAP7_75t_L g3127 ( 
.A1(n_2895),
.A2(n_2119),
.B(n_2126),
.C(n_2117),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2801),
.B(n_2117),
.Y(n_3128)
);

AOI21xp5_ASAP7_75t_L g3129 ( 
.A1(n_2803),
.A2(n_2281),
.B(n_2280),
.Y(n_3129)
);

BUFx8_ASAP7_75t_L g3130 ( 
.A(n_2849),
.Y(n_3130)
);

HB1xp67_ASAP7_75t_L g3131 ( 
.A(n_2849),
.Y(n_3131)
);

INVx2_ASAP7_75t_SL g3132 ( 
.A(n_2853),
.Y(n_3132)
);

AOI21xp5_ASAP7_75t_L g3133 ( 
.A1(n_2803),
.A2(n_2292),
.B(n_2284),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_SL g3134 ( 
.A(n_2830),
.B(n_2372),
.Y(n_3134)
);

NOR2xp33_ASAP7_75t_L g3135 ( 
.A(n_2794),
.B(n_1374),
.Y(n_3135)
);

OAI21xp5_ASAP7_75t_L g3136 ( 
.A1(n_2804),
.A2(n_2292),
.B(n_2284),
.Y(n_3136)
);

NOR2xp33_ASAP7_75t_L g3137 ( 
.A(n_2658),
.B(n_2560),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2678),
.B(n_2686),
.Y(n_3138)
);

AOI21xp5_ASAP7_75t_L g3139 ( 
.A1(n_2804),
.A2(n_2812),
.B(n_2807),
.Y(n_3139)
);

OAI22xp5_ASAP7_75t_L g3140 ( 
.A1(n_2936),
.A2(n_2715),
.B1(n_2719),
.B2(n_2687),
.Y(n_3140)
);

AOI21xp5_ASAP7_75t_L g3141 ( 
.A1(n_2949),
.A2(n_2941),
.B(n_2960),
.Y(n_3141)
);

AO22x1_ASAP7_75t_L g3142 ( 
.A1(n_2982),
.A2(n_2900),
.B1(n_2925),
.B2(n_2851),
.Y(n_3142)
);

BUFx12f_ASAP7_75t_L g3143 ( 
.A(n_3102),
.Y(n_3143)
);

OAI21xp5_ASAP7_75t_L g3144 ( 
.A1(n_3055),
.A2(n_2926),
.B(n_2812),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_SL g3145 ( 
.A(n_2984),
.B(n_2886),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_2937),
.B(n_2773),
.Y(n_3146)
);

OAI22xp5_ASAP7_75t_L g3147 ( 
.A1(n_2995),
.A2(n_3099),
.B1(n_2950),
.B2(n_2986),
.Y(n_3147)
);

AOI22xp33_ASAP7_75t_L g3148 ( 
.A1(n_3134),
.A2(n_2667),
.B1(n_2915),
.B2(n_2722),
.Y(n_3148)
);

NAND2x1p5_ASAP7_75t_L g3149 ( 
.A(n_2970),
.B(n_2903),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_SL g3150 ( 
.A(n_3034),
.B(n_2807),
.Y(n_3150)
);

OAI22xp5_ASAP7_75t_L g3151 ( 
.A1(n_2948),
.A2(n_2852),
.B1(n_2856),
.B2(n_2840),
.Y(n_3151)
);

BUFx2_ASAP7_75t_L g3152 ( 
.A(n_2972),
.Y(n_3152)
);

BUFx3_ASAP7_75t_L g3153 ( 
.A(n_3130),
.Y(n_3153)
);

O2A1O1Ixp33_ASAP7_75t_L g3154 ( 
.A1(n_3015),
.A2(n_2759),
.B(n_2842),
.C(n_2726),
.Y(n_3154)
);

NOR2xp67_ASAP7_75t_L g3155 ( 
.A(n_2974),
.B(n_2822),
.Y(n_3155)
);

O2A1O1Ixp5_ASAP7_75t_L g3156 ( 
.A1(n_2957),
.A2(n_2709),
.B(n_2823),
.C(n_2841),
.Y(n_3156)
);

INVx1_ASAP7_75t_SL g3157 ( 
.A(n_3016),
.Y(n_3157)
);

AOI21xp5_ASAP7_75t_L g3158 ( 
.A1(n_2964),
.A2(n_2885),
.B(n_2879),
.Y(n_3158)
);

AOI21xp5_ASAP7_75t_L g3159 ( 
.A1(n_2951),
.A2(n_2955),
.B(n_2958),
.Y(n_3159)
);

OR2x2_ASAP7_75t_L g3160 ( 
.A(n_3081),
.B(n_2781),
.Y(n_3160)
);

HB1xp67_ASAP7_75t_L g3161 ( 
.A(n_3072),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_SL g3162 ( 
.A(n_2981),
.B(n_2996),
.Y(n_3162)
);

O2A1O1Ixp33_ASAP7_75t_L g3163 ( 
.A1(n_3004),
.A2(n_3008),
.B(n_3123),
.C(n_3073),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2959),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_2946),
.B(n_2787),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_3086),
.B(n_2728),
.Y(n_3166)
);

NAND3xp33_ASAP7_75t_L g3167 ( 
.A(n_2992),
.B(n_2697),
.C(n_2775),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2939),
.B(n_2735),
.Y(n_3168)
);

AOI21xp5_ASAP7_75t_L g3169 ( 
.A1(n_3030),
.A2(n_2887),
.B(n_2738),
.Y(n_3169)
);

HB1xp67_ASAP7_75t_L g3170 ( 
.A(n_2945),
.Y(n_3170)
);

A2O1A1Ixp33_ASAP7_75t_L g3171 ( 
.A1(n_2979),
.A2(n_2864),
.B(n_2867),
.C(n_2862),
.Y(n_3171)
);

AOI21xp5_ASAP7_75t_L g3172 ( 
.A1(n_3139),
.A2(n_2837),
.B(n_2822),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_3138),
.Y(n_3173)
);

O2A1O1Ixp33_ASAP7_75t_SL g3174 ( 
.A1(n_3084),
.A2(n_2820),
.B(n_2927),
.C(n_2914),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2938),
.B(n_2737),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2940),
.B(n_2746),
.Y(n_3176)
);

INVx6_ASAP7_75t_L g3177 ( 
.A(n_3130),
.Y(n_3177)
);

AOI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_2965),
.A2(n_2837),
.B(n_2860),
.Y(n_3178)
);

OAI22xp5_ASAP7_75t_L g3179 ( 
.A1(n_2990),
.A2(n_2874),
.B1(n_2878),
.B2(n_2872),
.Y(n_3179)
);

AOI21xp5_ASAP7_75t_L g3180 ( 
.A1(n_2966),
.A2(n_2861),
.B(n_2860),
.Y(n_3180)
);

OR2x6_ASAP7_75t_SL g3181 ( 
.A(n_2956),
.B(n_782),
.Y(n_3181)
);

NAND2xp33_ASAP7_75t_L g3182 ( 
.A(n_3020),
.B(n_2685),
.Y(n_3182)
);

AOI21xp5_ASAP7_75t_L g3183 ( 
.A1(n_2966),
.A2(n_2902),
.B(n_2898),
.Y(n_3183)
);

INVx3_ASAP7_75t_L g3184 ( 
.A(n_3017),
.Y(n_3184)
);

O2A1O1Ixp33_ASAP7_75t_L g3185 ( 
.A1(n_3006),
.A2(n_2842),
.B(n_2753),
.C(n_2760),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2963),
.Y(n_3186)
);

A2O1A1Ixp33_ASAP7_75t_SL g3187 ( 
.A1(n_3135),
.A2(n_2698),
.B(n_2748),
.C(n_2761),
.Y(n_3187)
);

AOI21xp5_ASAP7_75t_L g3188 ( 
.A1(n_2962),
.A2(n_2870),
.B(n_2861),
.Y(n_3188)
);

A2O1A1Ixp33_ASAP7_75t_L g3189 ( 
.A1(n_3007),
.A2(n_2763),
.B(n_2771),
.C(n_2747),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2940),
.B(n_2785),
.Y(n_3190)
);

AND2x2_ASAP7_75t_L g3191 ( 
.A(n_3116),
.B(n_2790),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_3001),
.B(n_2805),
.Y(n_3192)
);

AOI22xp5_ASAP7_75t_L g3193 ( 
.A1(n_3000),
.A2(n_2592),
.B1(n_2392),
.B2(n_2579),
.Y(n_3193)
);

NOR2x1_ASAP7_75t_L g3194 ( 
.A(n_3107),
.B(n_3125),
.Y(n_3194)
);

NOR2xp33_ASAP7_75t_SL g3195 ( 
.A(n_3114),
.B(n_2522),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_2976),
.Y(n_3196)
);

AOI21xp5_ASAP7_75t_L g3197 ( 
.A1(n_3096),
.A2(n_2902),
.B(n_2898),
.Y(n_3197)
);

OAI21xp5_ASAP7_75t_L g3198 ( 
.A1(n_3003),
.A2(n_2875),
.B(n_2870),
.Y(n_3198)
);

NOR2xp67_ASAP7_75t_L g3199 ( 
.A(n_2993),
.B(n_2652),
.Y(n_3199)
);

AOI21xp5_ASAP7_75t_L g3200 ( 
.A1(n_3096),
.A2(n_2884),
.B(n_2875),
.Y(n_3200)
);

NOR2xp33_ASAP7_75t_L g3201 ( 
.A(n_3043),
.B(n_2831),
.Y(n_3201)
);

AOI21xp5_ASAP7_75t_L g3202 ( 
.A1(n_2954),
.A2(n_2884),
.B(n_2914),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_SL g3203 ( 
.A(n_3065),
.B(n_2792),
.Y(n_3203)
);

AOI21xp5_ASAP7_75t_L g3204 ( 
.A1(n_2954),
.A2(n_2827),
.B(n_2883),
.Y(n_3204)
);

AND2x2_ASAP7_75t_L g3205 ( 
.A(n_3112),
.B(n_2797),
.Y(n_3205)
);

NOR3xp33_ASAP7_75t_L g3206 ( 
.A(n_2994),
.B(n_2923),
.C(n_1224),
.Y(n_3206)
);

OAI22xp5_ASAP7_75t_L g3207 ( 
.A1(n_2998),
.A2(n_2808),
.B1(n_2818),
.B2(n_2806),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_SL g3208 ( 
.A(n_3058),
.B(n_2798),
.Y(n_3208)
);

AOI21xp5_ASAP7_75t_L g3209 ( 
.A1(n_3056),
.A2(n_2889),
.B(n_2888),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_2983),
.B(n_2821),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_SL g3211 ( 
.A(n_3042),
.B(n_2814),
.Y(n_3211)
);

AOI21xp5_ASAP7_75t_L g3212 ( 
.A1(n_3062),
.A2(n_2894),
.B(n_2892),
.Y(n_3212)
);

AOI21xp5_ASAP7_75t_SL g3213 ( 
.A1(n_3014),
.A2(n_2909),
.B(n_2903),
.Y(n_3213)
);

NOR2xp67_ASAP7_75t_L g3214 ( 
.A(n_3063),
.B(n_2657),
.Y(n_3214)
);

AND2x2_ASAP7_75t_SL g3215 ( 
.A(n_3021),
.B(n_2909),
.Y(n_3215)
);

AOI21x1_ASAP7_75t_L g3216 ( 
.A1(n_2971),
.A2(n_2896),
.B(n_2927),
.Y(n_3216)
);

OAI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_2978),
.A2(n_2928),
.B(n_2919),
.Y(n_3217)
);

AOI22xp5_ASAP7_75t_L g3218 ( 
.A1(n_3137),
.A2(n_2547),
.B1(n_2608),
.B2(n_2574),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2947),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_SL g3220 ( 
.A(n_3018),
.B(n_2826),
.Y(n_3220)
);

INVx2_ASAP7_75t_L g3221 ( 
.A(n_3012),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_3039),
.B(n_2835),
.Y(n_3222)
);

OAI21xp5_ASAP7_75t_L g3223 ( 
.A1(n_2987),
.A2(n_2931),
.B(n_2930),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_3023),
.Y(n_3224)
);

NOR3xp33_ASAP7_75t_L g3225 ( 
.A(n_3047),
.B(n_1225),
.C(n_1219),
.Y(n_3225)
);

NOR2xp33_ASAP7_75t_L g3226 ( 
.A(n_3027),
.B(n_2866),
.Y(n_3226)
);

INVx2_ASAP7_75t_SL g3227 ( 
.A(n_3036),
.Y(n_3227)
);

OAI21xp33_ASAP7_75t_L g3228 ( 
.A1(n_2989),
.A2(n_1083),
.B(n_1078),
.Y(n_3228)
);

AOI21xp5_ASAP7_75t_L g3229 ( 
.A1(n_2973),
.A2(n_3089),
.B(n_3051),
.Y(n_3229)
);

NOR2xp33_ASAP7_75t_L g3230 ( 
.A(n_3120),
.B(n_2765),
.Y(n_3230)
);

AOI22xp5_ASAP7_75t_L g3231 ( 
.A1(n_3013),
.A2(n_2566),
.B1(n_2659),
.B2(n_2916),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_3048),
.B(n_2661),
.Y(n_3232)
);

AND2x2_ASAP7_75t_L g3233 ( 
.A(n_3054),
.B(n_2675),
.Y(n_3233)
);

AOI21xp5_ASAP7_75t_L g3234 ( 
.A1(n_3050),
.A2(n_3046),
.B(n_2988),
.Y(n_3234)
);

AOI21xp5_ASAP7_75t_L g3235 ( 
.A1(n_2985),
.A2(n_2909),
.B(n_2916),
.Y(n_3235)
);

AOI21xp5_ASAP7_75t_L g3236 ( 
.A1(n_3005),
.A2(n_2916),
.B(n_2799),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_2968),
.B(n_2734),
.Y(n_3237)
);

AOI21xp5_ASAP7_75t_L g3238 ( 
.A1(n_3029),
.A2(n_3038),
.B(n_3044),
.Y(n_3238)
);

BUFx12f_ASAP7_75t_L g3239 ( 
.A(n_2942),
.Y(n_3239)
);

OAI21xp5_ASAP7_75t_L g3240 ( 
.A1(n_2943),
.A2(n_2294),
.B(n_2745),
.Y(n_3240)
);

AOI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_2991),
.A2(n_2799),
.B(n_2761),
.Y(n_3241)
);

OR2x6_ASAP7_75t_SL g3242 ( 
.A(n_2961),
.B(n_787),
.Y(n_3242)
);

NOR2xp33_ASAP7_75t_L g3243 ( 
.A(n_3068),
.B(n_2833),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_3009),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_3033),
.B(n_2749),
.Y(n_3245)
);

OAI21x1_ASAP7_75t_L g3246 ( 
.A1(n_3113),
.A2(n_2173),
.B(n_2171),
.Y(n_3246)
);

AOI21xp5_ASAP7_75t_L g3247 ( 
.A1(n_3002),
.A2(n_2868),
.B(n_2685),
.Y(n_3247)
);

A2O1A1Ixp33_ASAP7_75t_L g3248 ( 
.A1(n_3095),
.A2(n_2755),
.B(n_2764),
.C(n_2757),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_3022),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_3019),
.B(n_2769),
.Y(n_3250)
);

INVx3_ASAP7_75t_L g3251 ( 
.A(n_3017),
.Y(n_3251)
);

O2A1O1Ixp33_ASAP7_75t_L g3252 ( 
.A1(n_3088),
.A2(n_1530),
.B(n_1536),
.C(n_1487),
.Y(n_3252)
);

INVx2_ASAP7_75t_SL g3253 ( 
.A(n_3080),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_3031),
.B(n_2877),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3035),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_3054),
.B(n_1088),
.Y(n_3256)
);

NOR2xp33_ASAP7_75t_L g3257 ( 
.A(n_3053),
.B(n_2038),
.Y(n_3257)
);

AOI21x1_ASAP7_75t_L g3258 ( 
.A1(n_3104),
.A2(n_1849),
.B(n_1848),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3028),
.B(n_2877),
.Y(n_3259)
);

AOI21xp5_ASAP7_75t_L g3260 ( 
.A1(n_2952),
.A2(n_2868),
.B(n_2685),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3059),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_SL g3262 ( 
.A(n_2944),
.B(n_2685),
.Y(n_3262)
);

AOI21xp5_ASAP7_75t_L g3263 ( 
.A1(n_3110),
.A2(n_2868),
.B(n_2685),
.Y(n_3263)
);

CKINVDCx5p33_ASAP7_75t_R g3264 ( 
.A(n_3077),
.Y(n_3264)
);

AND2x4_ASAP7_75t_L g3265 ( 
.A(n_2977),
.B(n_2294),
.Y(n_3265)
);

OAI22xp5_ASAP7_75t_L g3266 ( 
.A1(n_3057),
.A2(n_2176),
.B1(n_2228),
.B2(n_2173),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_SL g3267 ( 
.A(n_2944),
.B(n_2685),
.Y(n_3267)
);

AOI21xp5_ASAP7_75t_L g3268 ( 
.A1(n_2980),
.A2(n_2868),
.B(n_2126),
.Y(n_3268)
);

NOR2xp67_ASAP7_75t_L g3269 ( 
.A(n_3075),
.B(n_2228),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3083),
.Y(n_3270)
);

OAI21xp5_ASAP7_75t_L g3271 ( 
.A1(n_2943),
.A2(n_1851),
.B(n_1848),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_L g3272 ( 
.A(n_3079),
.B(n_1536),
.Y(n_3272)
);

OAI22xp5_ASAP7_75t_L g3273 ( 
.A1(n_3132),
.A2(n_2240),
.B1(n_2176),
.B2(n_2228),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_3119),
.B(n_1551),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_3121),
.B(n_1551),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_SL g3276 ( 
.A(n_3066),
.B(n_2868),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_3097),
.B(n_1554),
.Y(n_3277)
);

A2O1A1Ixp33_ASAP7_75t_SL g3278 ( 
.A1(n_3010),
.A2(n_1580),
.B(n_1554),
.C(n_2173),
.Y(n_3278)
);

AO21x1_ASAP7_75t_L g3279 ( 
.A1(n_3025),
.A2(n_1854),
.B(n_1851),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_3098),
.B(n_1580),
.Y(n_3280)
);

NAND2xp33_ASAP7_75t_L g3281 ( 
.A(n_2942),
.B(n_2868),
.Y(n_3281)
);

AOI21xp5_ASAP7_75t_L g3282 ( 
.A1(n_2980),
.A2(n_2127),
.B(n_2119),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_3115),
.Y(n_3283)
);

AOI21xp5_ASAP7_75t_L g3284 ( 
.A1(n_3045),
.A2(n_2128),
.B(n_2127),
.Y(n_3284)
);

OAI22xp5_ASAP7_75t_L g3285 ( 
.A1(n_3126),
.A2(n_788),
.B1(n_791),
.B2(n_789),
.Y(n_3285)
);

OAI21x1_ASAP7_75t_L g3286 ( 
.A1(n_2969),
.A2(n_2232),
.B(n_2176),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3069),
.B(n_2128),
.Y(n_3287)
);

AOI22xp33_ASAP7_75t_L g3288 ( 
.A1(n_3026),
.A2(n_1220),
.B1(n_1228),
.B2(n_1172),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_2977),
.B(n_2132),
.Y(n_3289)
);

AND2x4_ASAP7_75t_L g3290 ( 
.A(n_2997),
.B(n_2569),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_SL g3291 ( 
.A(n_2999),
.B(n_2132),
.Y(n_3291)
);

AOI21xp5_ASAP7_75t_L g3292 ( 
.A1(n_3040),
.A2(n_2139),
.B(n_2136),
.Y(n_3292)
);

AOI21xp5_ASAP7_75t_L g3293 ( 
.A1(n_3041),
.A2(n_3025),
.B(n_3070),
.Y(n_3293)
);

OAI21xp5_ASAP7_75t_L g3294 ( 
.A1(n_3060),
.A2(n_1858),
.B(n_1854),
.Y(n_3294)
);

INVx3_ASAP7_75t_L g3295 ( 
.A(n_3014),
.Y(n_3295)
);

BUFx3_ASAP7_75t_L g3296 ( 
.A(n_2942),
.Y(n_3296)
);

NOR2xp33_ASAP7_75t_L g3297 ( 
.A(n_3131),
.B(n_1235),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_2997),
.B(n_2136),
.Y(n_3298)
);

AND2x2_ASAP7_75t_L g3299 ( 
.A(n_3087),
.B(n_2967),
.Y(n_3299)
);

AOI21xp5_ASAP7_75t_L g3300 ( 
.A1(n_3074),
.A2(n_2146),
.B(n_2139),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_SL g3301 ( 
.A(n_3087),
.B(n_2146),
.Y(n_3301)
);

NOR2xp33_ASAP7_75t_L g3302 ( 
.A(n_3037),
.B(n_1247),
.Y(n_3302)
);

AND2x2_ASAP7_75t_L g3303 ( 
.A(n_2967),
.B(n_1231),
.Y(n_3303)
);

AOI21xp5_ASAP7_75t_L g3304 ( 
.A1(n_3076),
.A2(n_2163),
.B(n_2160),
.Y(n_3304)
);

OA22x2_ASAP7_75t_L g3305 ( 
.A1(n_3014),
.A2(n_796),
.B1(n_797),
.B2(n_794),
.Y(n_3305)
);

AOI21xp5_ASAP7_75t_L g3306 ( 
.A1(n_3082),
.A2(n_2163),
.B(n_2160),
.Y(n_3306)
);

AND2x2_ASAP7_75t_L g3307 ( 
.A(n_2967),
.B(n_1232),
.Y(n_3307)
);

OAI22xp5_ASAP7_75t_L g3308 ( 
.A1(n_3032),
.A2(n_2240),
.B1(n_2275),
.B2(n_2232),
.Y(n_3308)
);

AO21x1_ASAP7_75t_L g3309 ( 
.A1(n_2975),
.A2(n_1859),
.B(n_1858),
.Y(n_3309)
);

CKINVDCx6p67_ASAP7_75t_R g3310 ( 
.A(n_3114),
.Y(n_3310)
);

AOI21xp5_ASAP7_75t_L g3311 ( 
.A1(n_3064),
.A2(n_2169),
.B(n_2165),
.Y(n_3311)
);

NOR2x1_ASAP7_75t_L g3312 ( 
.A(n_2970),
.B(n_2093),
.Y(n_3312)
);

OAI22xp5_ASAP7_75t_L g3313 ( 
.A1(n_3049),
.A2(n_2232),
.B1(n_2275),
.B2(n_2240),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_3071),
.B(n_2165),
.Y(n_3314)
);

AND2x4_ASAP7_75t_L g3315 ( 
.A(n_3049),
.B(n_2569),
.Y(n_3315)
);

OR2x6_ASAP7_75t_SL g3316 ( 
.A(n_2953),
.B(n_798),
.Y(n_3316)
);

NOR3xp33_ASAP7_75t_L g3317 ( 
.A(n_3061),
.B(n_1234),
.C(n_1233),
.Y(n_3317)
);

AOI21xp5_ASAP7_75t_L g3318 ( 
.A1(n_3101),
.A2(n_2169),
.B(n_2096),
.Y(n_3318)
);

CKINVDCx5p33_ASAP7_75t_R g3319 ( 
.A(n_3061),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3078),
.Y(n_3320)
);

OAI21xp5_ASAP7_75t_L g3321 ( 
.A1(n_3127),
.A2(n_1879),
.B(n_1859),
.Y(n_3321)
);

AOI22xp33_ASAP7_75t_L g3322 ( 
.A1(n_3085),
.A2(n_1525),
.B1(n_1907),
.B2(n_1879),
.Y(n_3322)
);

INVx1_ASAP7_75t_SL g3323 ( 
.A(n_3090),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3101),
.Y(n_3324)
);

AOI21xp5_ASAP7_75t_L g3325 ( 
.A1(n_3105),
.A2(n_2096),
.B(n_2093),
.Y(n_3325)
);

OAI22xp5_ASAP7_75t_L g3326 ( 
.A1(n_3105),
.A2(n_801),
.B1(n_805),
.B2(n_802),
.Y(n_3326)
);

AOI22xp5_ASAP7_75t_L g3327 ( 
.A1(n_3011),
.A2(n_749),
.B1(n_750),
.B2(n_743),
.Y(n_3327)
);

NOR2xp33_ASAP7_75t_L g3328 ( 
.A(n_3024),
.B(n_754),
.Y(n_3328)
);

OAI21xp5_ASAP7_75t_L g3329 ( 
.A1(n_3122),
.A2(n_1908),
.B(n_1907),
.Y(n_3329)
);

AND2x2_ASAP7_75t_SL g3330 ( 
.A(n_3106),
.B(n_1236),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_SL g3331 ( 
.A(n_3106),
.B(n_2278),
.Y(n_3331)
);

NOR2xp33_ASAP7_75t_R g3332 ( 
.A(n_3103),
.B(n_2631),
.Y(n_3332)
);

INVxp67_ASAP7_75t_L g3333 ( 
.A(n_3108),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3108),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3109),
.Y(n_3335)
);

AOI21xp5_ASAP7_75t_L g3336 ( 
.A1(n_3109),
.A2(n_3128),
.B(n_3124),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3124),
.Y(n_3337)
);

A2O1A1Ixp33_ASAP7_75t_L g3338 ( 
.A1(n_3100),
.A2(n_1911),
.B(n_1908),
.C(n_1765),
.Y(n_3338)
);

OR2x2_ASAP7_75t_L g3339 ( 
.A(n_3128),
.B(n_1238),
.Y(n_3339)
);

O2A1O1Ixp33_ASAP7_75t_SL g3340 ( 
.A1(n_3094),
.A2(n_1911),
.B(n_1770),
.C(n_1776),
.Y(n_3340)
);

AOI21xp5_ASAP7_75t_L g3341 ( 
.A1(n_3093),
.A2(n_2096),
.B(n_2093),
.Y(n_3341)
);

AOI22xp5_ASAP7_75t_L g3342 ( 
.A1(n_3111),
.A2(n_759),
.B1(n_772),
.B2(n_758),
.Y(n_3342)
);

BUFx8_ASAP7_75t_L g3343 ( 
.A(n_3227),
.Y(n_3343)
);

OAI21x1_ASAP7_75t_L g3344 ( 
.A1(n_3258),
.A2(n_3133),
.B(n_3129),
.Y(n_3344)
);

OAI21x1_ASAP7_75t_L g3345 ( 
.A1(n_3293),
.A2(n_3052),
.B(n_3118),
.Y(n_3345)
);

INVxp67_ASAP7_75t_SL g3346 ( 
.A(n_3161),
.Y(n_3346)
);

OR2x2_ASAP7_75t_L g3347 ( 
.A(n_3160),
.B(n_3136),
.Y(n_3347)
);

INVx6_ASAP7_75t_SL g3348 ( 
.A(n_3290),
.Y(n_3348)
);

OAI21x1_ASAP7_75t_L g3349 ( 
.A1(n_3159),
.A2(n_3117),
.B(n_3067),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_3173),
.B(n_809),
.Y(n_3350)
);

INVx3_ASAP7_75t_L g3351 ( 
.A(n_3184),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3219),
.Y(n_3352)
);

AOI21xp5_ASAP7_75t_L g3353 ( 
.A1(n_3229),
.A2(n_3092),
.B(n_3091),
.Y(n_3353)
);

NAND2x1p5_ASAP7_75t_L g3354 ( 
.A(n_3157),
.B(n_3152),
.Y(n_3354)
);

AOI21x1_ASAP7_75t_L g3355 ( 
.A1(n_3162),
.A2(n_3260),
.B(n_3216),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3205),
.B(n_813),
.Y(n_3356)
);

NAND3xp33_ASAP7_75t_L g3357 ( 
.A(n_3328),
.B(n_817),
.C(n_814),
.Y(n_3357)
);

OAI21x1_ASAP7_75t_L g3358 ( 
.A1(n_3141),
.A2(n_2278),
.B(n_2275),
.Y(n_3358)
);

AOI221x1_ASAP7_75t_L g3359 ( 
.A1(n_3147),
.A2(n_1244),
.B1(n_1246),
.B2(n_1243),
.C(n_1239),
.Y(n_3359)
);

BUFx12f_ASAP7_75t_L g3360 ( 
.A(n_3143),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_3283),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3244),
.Y(n_3362)
);

OAI21xp5_ASAP7_75t_L g3363 ( 
.A1(n_3163),
.A2(n_1780),
.B(n_1762),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3146),
.B(n_1249),
.Y(n_3364)
);

AOI21xp5_ASAP7_75t_L g3365 ( 
.A1(n_3238),
.A2(n_1867),
.B(n_1861),
.Y(n_3365)
);

A2O1A1Ixp33_ASAP7_75t_L g3366 ( 
.A1(n_3154),
.A2(n_1251),
.B(n_1253),
.C(n_1250),
.Y(n_3366)
);

OAI21x1_ASAP7_75t_L g3367 ( 
.A1(n_3263),
.A2(n_2278),
.B(n_2110),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_3168),
.B(n_820),
.Y(n_3368)
);

OAI21x1_ASAP7_75t_SL g3369 ( 
.A1(n_3185),
.A2(n_1255),
.B(n_1254),
.Y(n_3369)
);

INVx1_ASAP7_75t_SL g3370 ( 
.A(n_3157),
.Y(n_3370)
);

BUFx2_ASAP7_75t_L g3371 ( 
.A(n_3264),
.Y(n_3371)
);

CKINVDCx6p67_ASAP7_75t_R g3372 ( 
.A(n_3153),
.Y(n_3372)
);

INVx5_ASAP7_75t_L g3373 ( 
.A(n_3177),
.Y(n_3373)
);

OAI21xp33_ASAP7_75t_L g3374 ( 
.A1(n_3330),
.A2(n_823),
.B(n_822),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_SL g3375 ( 
.A(n_3215),
.B(n_1578),
.Y(n_3375)
);

OAI21x1_ASAP7_75t_L g3376 ( 
.A1(n_3234),
.A2(n_2110),
.B(n_2098),
.Y(n_3376)
);

INVx2_ASAP7_75t_L g3377 ( 
.A(n_3164),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3249),
.Y(n_3378)
);

BUFx6f_ASAP7_75t_L g3379 ( 
.A(n_3239),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3255),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3323),
.B(n_827),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_3323),
.B(n_832),
.Y(n_3382)
);

AOI21xp5_ASAP7_75t_L g3383 ( 
.A1(n_3182),
.A2(n_1868),
.B(n_1867),
.Y(n_3383)
);

INVx1_ASAP7_75t_SL g3384 ( 
.A(n_3170),
.Y(n_3384)
);

AOI21xp5_ASAP7_75t_SL g3385 ( 
.A1(n_3211),
.A2(n_1809),
.B(n_1798),
.Y(n_3385)
);

AND2x4_ASAP7_75t_L g3386 ( 
.A(n_3295),
.B(n_3184),
.Y(n_3386)
);

OAI21x1_ASAP7_75t_L g3387 ( 
.A1(n_3246),
.A2(n_2110),
.B(n_2098),
.Y(n_3387)
);

AND2x2_ASAP7_75t_L g3388 ( 
.A(n_3233),
.B(n_1256),
.Y(n_3388)
);

AOI21xp5_ASAP7_75t_L g3389 ( 
.A1(n_3172),
.A2(n_1869),
.B(n_1868),
.Y(n_3389)
);

OAI22xp5_ASAP7_75t_L g3390 ( 
.A1(n_3148),
.A2(n_835),
.B1(n_840),
.B2(n_833),
.Y(n_3390)
);

A2O1A1Ixp33_ASAP7_75t_L g3391 ( 
.A1(n_3302),
.A2(n_1258),
.B(n_1259),
.C(n_1257),
.Y(n_3391)
);

OAI22xp5_ASAP7_75t_L g3392 ( 
.A1(n_3167),
.A2(n_3257),
.B1(n_3231),
.B2(n_3214),
.Y(n_3392)
);

BUFx3_ASAP7_75t_L g3393 ( 
.A(n_3177),
.Y(n_3393)
);

INVx3_ASAP7_75t_L g3394 ( 
.A(n_3251),
.Y(n_3394)
);

INVx2_ASAP7_75t_L g3395 ( 
.A(n_3186),
.Y(n_3395)
);

AOI21xp5_ASAP7_75t_L g3396 ( 
.A1(n_3197),
.A2(n_1871),
.B(n_1869),
.Y(n_3396)
);

INVx4_ASAP7_75t_L g3397 ( 
.A(n_3177),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3175),
.B(n_844),
.Y(n_3398)
);

BUFx12f_ASAP7_75t_L g3399 ( 
.A(n_3253),
.Y(n_3399)
);

OAI21x1_ASAP7_75t_L g3400 ( 
.A1(n_3268),
.A2(n_2121),
.B(n_2098),
.Y(n_3400)
);

OAI21x1_ASAP7_75t_L g3401 ( 
.A1(n_3247),
.A2(n_2124),
.B(n_2121),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3192),
.B(n_845),
.Y(n_3402)
);

AOI31xp67_ASAP7_75t_L g3403 ( 
.A1(n_3145),
.A2(n_1871),
.A3(n_1875),
.B(n_1873),
.Y(n_3403)
);

INVx3_ASAP7_75t_L g3404 ( 
.A(n_3251),
.Y(n_3404)
);

AOI21xp5_ASAP7_75t_L g3405 ( 
.A1(n_3200),
.A2(n_1875),
.B(n_1873),
.Y(n_3405)
);

AOI21x1_ASAP7_75t_SL g3406 ( 
.A1(n_3166),
.A2(n_2),
.B(n_3),
.Y(n_3406)
);

AO21x2_ASAP7_75t_L g3407 ( 
.A1(n_3309),
.A2(n_1811),
.B(n_1810),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_3196),
.Y(n_3408)
);

AO31x2_ASAP7_75t_L g3409 ( 
.A1(n_3279),
.A2(n_1878),
.A3(n_1814),
.B(n_1823),
.Y(n_3409)
);

OAI22x1_ASAP7_75t_L g3410 ( 
.A1(n_3165),
.A2(n_849),
.B1(n_857),
.B2(n_847),
.Y(n_3410)
);

OAI21x1_ASAP7_75t_L g3411 ( 
.A1(n_3286),
.A2(n_2124),
.B(n_2121),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_3210),
.B(n_860),
.Y(n_3412)
);

AO31x2_ASAP7_75t_L g3413 ( 
.A1(n_3180),
.A2(n_1878),
.A3(n_1826),
.B(n_1834),
.Y(n_3413)
);

AOI21xp5_ASAP7_75t_SL g3414 ( 
.A1(n_3189),
.A2(n_1836),
.B(n_1813),
.Y(n_3414)
);

OAI21x1_ASAP7_75t_L g3415 ( 
.A1(n_3282),
.A2(n_2124),
.B(n_1886),
.Y(n_3415)
);

OAI21x1_ASAP7_75t_L g3416 ( 
.A1(n_3209),
.A2(n_1886),
.B(n_1884),
.Y(n_3416)
);

OAI22xp5_ASAP7_75t_L g3417 ( 
.A1(n_3218),
.A2(n_863),
.B1(n_865),
.B2(n_862),
.Y(n_3417)
);

AOI211x1_ASAP7_75t_L g3418 ( 
.A1(n_3142),
.A2(n_1262),
.B(n_1266),
.C(n_1260),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3261),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_3270),
.Y(n_3420)
);

BUFx6f_ASAP7_75t_L g3421 ( 
.A(n_3296),
.Y(n_3421)
);

OAI21x1_ASAP7_75t_L g3422 ( 
.A1(n_3212),
.A2(n_1887),
.B(n_1884),
.Y(n_3422)
);

BUFx6f_ASAP7_75t_L g3423 ( 
.A(n_3299),
.Y(n_3423)
);

AND2x2_ASAP7_75t_L g3424 ( 
.A(n_3191),
.B(n_1267),
.Y(n_3424)
);

AND2x2_ASAP7_75t_L g3425 ( 
.A(n_3303),
.B(n_3307),
.Y(n_3425)
);

AND2x2_ASAP7_75t_L g3426 ( 
.A(n_3221),
.B(n_1268),
.Y(n_3426)
);

HB1xp67_ASAP7_75t_L g3427 ( 
.A(n_3179),
.Y(n_3427)
);

HB1xp67_ASAP7_75t_L g3428 ( 
.A(n_3199),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3217),
.Y(n_3429)
);

OAI22x1_ASAP7_75t_L g3430 ( 
.A1(n_3194),
.A2(n_882),
.B1(n_887),
.B2(n_869),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_SL g3431 ( 
.A(n_3206),
.B(n_1583),
.Y(n_3431)
);

AND2x2_ASAP7_75t_L g3432 ( 
.A(n_3224),
.B(n_1269),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3222),
.B(n_889),
.Y(n_3433)
);

BUFx2_ASAP7_75t_L g3434 ( 
.A(n_3319),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3150),
.B(n_890),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_3237),
.Y(n_3436)
);

AOI221xp5_ASAP7_75t_L g3437 ( 
.A1(n_3326),
.A2(n_899),
.B1(n_906),
.B2(n_893),
.C(n_891),
.Y(n_3437)
);

OAI21x1_ASAP7_75t_L g3438 ( 
.A1(n_3241),
.A2(n_1890),
.B(n_1887),
.Y(n_3438)
);

BUFx3_ASAP7_75t_L g3439 ( 
.A(n_3256),
.Y(n_3439)
);

INVx1_ASAP7_75t_SL g3440 ( 
.A(n_3297),
.Y(n_3440)
);

AOI21x1_ASAP7_75t_L g3441 ( 
.A1(n_3235),
.A2(n_1863),
.B(n_1862),
.Y(n_3441)
);

AOI21xp33_ASAP7_75t_L g3442 ( 
.A1(n_3342),
.A2(n_1882),
.B(n_1870),
.Y(n_3442)
);

NOR2xp67_ASAP7_75t_L g3443 ( 
.A(n_3236),
.B(n_1885),
.Y(n_3443)
);

OAI21x1_ASAP7_75t_L g3444 ( 
.A1(n_3178),
.A2(n_1897),
.B(n_1890),
.Y(n_3444)
);

OAI21x1_ASAP7_75t_L g3445 ( 
.A1(n_3284),
.A2(n_1905),
.B(n_1897),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3176),
.B(n_907),
.Y(n_3446)
);

AOI21xp5_ASAP7_75t_L g3447 ( 
.A1(n_3174),
.A2(n_1898),
.B(n_1889),
.Y(n_3447)
);

OAI21x1_ASAP7_75t_L g3448 ( 
.A1(n_3292),
.A2(n_1910),
.B(n_1905),
.Y(n_3448)
);

OAI21x1_ASAP7_75t_L g3449 ( 
.A1(n_3329),
.A2(n_1915),
.B(n_1910),
.Y(n_3449)
);

AO31x2_ASAP7_75t_L g3450 ( 
.A1(n_3183),
.A2(n_1900),
.A3(n_1922),
.B(n_1899),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_3259),
.Y(n_3451)
);

BUFx4f_ASAP7_75t_L g3452 ( 
.A(n_3310),
.Y(n_3452)
);

BUFx6f_ASAP7_75t_L g3453 ( 
.A(n_3290),
.Y(n_3453)
);

OAI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_3181),
.A2(n_914),
.B1(n_920),
.B2(n_913),
.Y(n_3454)
);

AOI21xp5_ASAP7_75t_L g3455 ( 
.A1(n_3188),
.A2(n_1931),
.B(n_1924),
.Y(n_3455)
);

OAI21xp33_ASAP7_75t_SL g3456 ( 
.A1(n_3144),
.A2(n_3198),
.B(n_3324),
.Y(n_3456)
);

CKINVDCx16_ASAP7_75t_R g3457 ( 
.A(n_3316),
.Y(n_3457)
);

AOI21xp5_ASAP7_75t_L g3458 ( 
.A1(n_3202),
.A2(n_1941),
.B(n_1938),
.Y(n_3458)
);

A2O1A1Ixp33_ASAP7_75t_L g3459 ( 
.A1(n_3144),
.A2(n_1273),
.B(n_1274),
.C(n_1270),
.Y(n_3459)
);

AOI21xp5_ASAP7_75t_L g3460 ( 
.A1(n_3281),
.A2(n_3158),
.B(n_3204),
.Y(n_3460)
);

INVx3_ASAP7_75t_L g3461 ( 
.A(n_3149),
.Y(n_3461)
);

O2A1O1Ixp5_ASAP7_75t_L g3462 ( 
.A1(n_3156),
.A2(n_1275),
.B(n_1942),
.C(n_1917),
.Y(n_3462)
);

INVxp67_ASAP7_75t_SL g3463 ( 
.A(n_3333),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3217),
.Y(n_3464)
);

AOI21x1_ASAP7_75t_L g3465 ( 
.A1(n_3300),
.A2(n_1917),
.B(n_1915),
.Y(n_3465)
);

OAI21x1_ASAP7_75t_L g3466 ( 
.A1(n_3329),
.A2(n_1921),
.B(n_1920),
.Y(n_3466)
);

OAI21xp5_ASAP7_75t_L g3467 ( 
.A1(n_3327),
.A2(n_2631),
.B(n_779),
.Y(n_3467)
);

HB1xp67_ASAP7_75t_L g3468 ( 
.A(n_3254),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_3190),
.B(n_922),
.Y(n_3469)
);

OAI21xp33_ASAP7_75t_SL g3470 ( 
.A1(n_3198),
.A2(n_1921),
.B(n_1920),
.Y(n_3470)
);

AOI221x1_ASAP7_75t_L g3471 ( 
.A1(n_3151),
.A2(n_1598),
.B1(n_1587),
.B2(n_1597),
.C(n_1585),
.Y(n_3471)
);

AOI21xp5_ASAP7_75t_L g3472 ( 
.A1(n_3169),
.A2(n_1933),
.B(n_1929),
.Y(n_3472)
);

OAI21x1_ASAP7_75t_L g3473 ( 
.A1(n_3304),
.A2(n_1933),
.B(n_1929),
.Y(n_3473)
);

OAI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_3171),
.A2(n_2631),
.B(n_781),
.Y(n_3474)
);

OAI21x1_ASAP7_75t_L g3475 ( 
.A1(n_3306),
.A2(n_1935),
.B(n_1934),
.Y(n_3475)
);

OAI21x1_ASAP7_75t_L g3476 ( 
.A1(n_3311),
.A2(n_1935),
.B(n_1934),
.Y(n_3476)
);

INVx3_ASAP7_75t_L g3477 ( 
.A(n_3149),
.Y(n_3477)
);

AND2x4_ASAP7_75t_L g3478 ( 
.A(n_3295),
.B(n_2631),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_L g3479 ( 
.A(n_3250),
.B(n_924),
.Y(n_3479)
);

OAI21x1_ASAP7_75t_L g3480 ( 
.A1(n_3341),
.A2(n_1633),
.B(n_1621),
.Y(n_3480)
);

AO21x1_ASAP7_75t_L g3481 ( 
.A1(n_3140),
.A2(n_1598),
.B(n_3),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_3272),
.Y(n_3482)
);

AOI21xp5_ASAP7_75t_L g3483 ( 
.A1(n_3336),
.A2(n_1633),
.B(n_1621),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3334),
.Y(n_3484)
);

NOR2xp33_ASAP7_75t_L g3485 ( 
.A(n_3201),
.B(n_775),
.Y(n_3485)
);

INVx1_ASAP7_75t_SL g3486 ( 
.A(n_3226),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3232),
.B(n_926),
.Y(n_3487)
);

OAI21x1_ASAP7_75t_L g3488 ( 
.A1(n_3325),
.A2(n_1633),
.B(n_1621),
.Y(n_3488)
);

OR2x2_ASAP7_75t_L g3489 ( 
.A(n_3335),
.B(n_3337),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_3320),
.B(n_1583),
.Y(n_3490)
);

INVx3_ASAP7_75t_L g3491 ( 
.A(n_3265),
.Y(n_3491)
);

OAI21x1_ASAP7_75t_L g3492 ( 
.A1(n_3318),
.A2(n_1671),
.B(n_1658),
.Y(n_3492)
);

AO32x2_ASAP7_75t_L g3493 ( 
.A1(n_3140),
.A2(n_6),
.A3(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_3493)
);

OAI22x1_ASAP7_75t_L g3494 ( 
.A1(n_3243),
.A2(n_790),
.B1(n_792),
.B2(n_785),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3245),
.B(n_1583),
.Y(n_3495)
);

AO31x2_ASAP7_75t_L g3496 ( 
.A1(n_3338),
.A2(n_1743),
.A3(n_1385),
.B(n_1367),
.Y(n_3496)
);

INVx5_ASAP7_75t_L g3497 ( 
.A(n_3315),
.Y(n_3497)
);

BUFx6f_ASAP7_75t_L g3498 ( 
.A(n_3265),
.Y(n_3498)
);

AOI21xp5_ASAP7_75t_L g3499 ( 
.A1(n_3187),
.A2(n_1671),
.B(n_1658),
.Y(n_3499)
);

OAI21xp5_ASAP7_75t_L g3500 ( 
.A1(n_3271),
.A2(n_804),
.B(n_795),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3203),
.B(n_1583),
.Y(n_3501)
);

OAI21xp5_ASAP7_75t_L g3502 ( 
.A1(n_3271),
.A2(n_825),
.B(n_808),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3262),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3220),
.B(n_1585),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_SL g3505 ( 
.A(n_3305),
.B(n_1585),
.Y(n_3505)
);

OAI21xp5_ASAP7_75t_L g3506 ( 
.A1(n_3225),
.A2(n_828),
.B(n_826),
.Y(n_3506)
);

OAI21x1_ASAP7_75t_L g3507 ( 
.A1(n_3294),
.A2(n_1671),
.B(n_1658),
.Y(n_3507)
);

AO31x2_ASAP7_75t_L g3508 ( 
.A1(n_3308),
.A2(n_1743),
.A3(n_1385),
.B(n_1367),
.Y(n_3508)
);

AND2x2_ASAP7_75t_L g3509 ( 
.A(n_3242),
.B(n_829),
.Y(n_3509)
);

OAI21x1_ASAP7_75t_L g3510 ( 
.A1(n_3294),
.A2(n_1735),
.B(n_1723),
.Y(n_3510)
);

OAI21x1_ASAP7_75t_L g3511 ( 
.A1(n_3321),
.A2(n_1735),
.B(n_1723),
.Y(n_3511)
);

HB1xp67_ASAP7_75t_L g3512 ( 
.A(n_3267),
.Y(n_3512)
);

AOI21xp5_ASAP7_75t_L g3513 ( 
.A1(n_3291),
.A2(n_1735),
.B(n_1723),
.Y(n_3513)
);

AO31x2_ASAP7_75t_L g3514 ( 
.A1(n_3248),
.A2(n_3313),
.A3(n_3207),
.B(n_3266),
.Y(n_3514)
);

BUFx6f_ASAP7_75t_L g3515 ( 
.A(n_3315),
.Y(n_3515)
);

AND2x4_ASAP7_75t_L g3516 ( 
.A(n_3155),
.B(n_283),
.Y(n_3516)
);

AO31x2_ASAP7_75t_L g3517 ( 
.A1(n_3273),
.A2(n_3314),
.A3(n_3278),
.B(n_3287),
.Y(n_3517)
);

AOI22xp5_ASAP7_75t_L g3518 ( 
.A1(n_3317),
.A2(n_843),
.B1(n_848),
.B2(n_841),
.Y(n_3518)
);

AOI21xp5_ASAP7_75t_L g3519 ( 
.A1(n_3223),
.A2(n_1773),
.B(n_1748),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3208),
.B(n_1585),
.Y(n_3520)
);

AOI21x1_ASAP7_75t_L g3521 ( 
.A1(n_3331),
.A2(n_1773),
.B(n_1748),
.Y(n_3521)
);

INVx3_ASAP7_75t_L g3522 ( 
.A(n_3289),
.Y(n_3522)
);

O2A1O1Ixp5_ASAP7_75t_L g3523 ( 
.A1(n_3276),
.A2(n_1773),
.B(n_1806),
.C(n_1748),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_L g3524 ( 
.A(n_3339),
.B(n_1587),
.Y(n_3524)
);

AO31x2_ASAP7_75t_L g3525 ( 
.A1(n_3277),
.A2(n_1743),
.A3(n_1385),
.B(n_1367),
.Y(n_3525)
);

CKINVDCx5p33_ASAP7_75t_R g3526 ( 
.A(n_3230),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_3326),
.B(n_1587),
.Y(n_3527)
);

BUFx3_ASAP7_75t_L g3528 ( 
.A(n_3193),
.Y(n_3528)
);

NOR2x1_ASAP7_75t_SL g3529 ( 
.A(n_3301),
.B(n_1587),
.Y(n_3529)
);

INVx1_ASAP7_75t_SL g3530 ( 
.A(n_3298),
.Y(n_3530)
);

OAI21x1_ASAP7_75t_L g3531 ( 
.A1(n_3321),
.A2(n_1828),
.B(n_1806),
.Y(n_3531)
);

CKINVDCx5p33_ASAP7_75t_R g3532 ( 
.A(n_3213),
.Y(n_3532)
);

INVx2_ASAP7_75t_SL g3533 ( 
.A(n_3305),
.Y(n_3533)
);

OR2x2_ASAP7_75t_L g3534 ( 
.A(n_3280),
.B(n_1597),
.Y(n_3534)
);

INVx4_ASAP7_75t_L g3535 ( 
.A(n_3195),
.Y(n_3535)
);

OAI21xp5_ASAP7_75t_L g3536 ( 
.A1(n_3223),
.A2(n_853),
.B(n_851),
.Y(n_3536)
);

OAI21x1_ASAP7_75t_L g3537 ( 
.A1(n_3240),
.A2(n_1828),
.B(n_1806),
.Y(n_3537)
);

A2O1A1Ixp33_ASAP7_75t_L g3538 ( 
.A1(n_3228),
.A2(n_859),
.B(n_861),
.C(n_856),
.Y(n_3538)
);

AOI21xp5_ASAP7_75t_L g3539 ( 
.A1(n_3340),
.A2(n_1835),
.B(n_1828),
.Y(n_3539)
);

INVxp67_ASAP7_75t_L g3540 ( 
.A(n_3274),
.Y(n_3540)
);

OA21x2_ASAP7_75t_L g3541 ( 
.A1(n_3240),
.A2(n_3322),
.B(n_3275),
.Y(n_3541)
);

AOI21xp5_ASAP7_75t_L g3542 ( 
.A1(n_3252),
.A2(n_1864),
.B(n_1835),
.Y(n_3542)
);

NOR2x1_ASAP7_75t_L g3543 ( 
.A(n_3312),
.B(n_1835),
.Y(n_3543)
);

OAI21xp5_ASAP7_75t_L g3544 ( 
.A1(n_3288),
.A2(n_874),
.B(n_873),
.Y(n_3544)
);

AO21x2_ASAP7_75t_L g3545 ( 
.A1(n_3332),
.A2(n_878),
.B(n_876),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3269),
.Y(n_3546)
);

NOR2xp33_ASAP7_75t_L g3547 ( 
.A(n_3195),
.B(n_881),
.Y(n_3547)
);

OAI21x1_ASAP7_75t_L g3548 ( 
.A1(n_3285),
.A2(n_1866),
.B(n_1864),
.Y(n_3548)
);

A2O1A1Ixp33_ASAP7_75t_L g3549 ( 
.A1(n_3285),
.A2(n_896),
.B(n_900),
.C(n_885),
.Y(n_3549)
);

INVx3_ASAP7_75t_L g3550 ( 
.A(n_3184),
.Y(n_3550)
);

AND2x2_ASAP7_75t_L g3551 ( 
.A(n_3205),
.B(n_902),
.Y(n_3551)
);

OAI21x1_ASAP7_75t_L g3552 ( 
.A1(n_3258),
.A2(n_1866),
.B(n_1864),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3173),
.B(n_1597),
.Y(n_3553)
);

OR2x6_ASAP7_75t_L g3554 ( 
.A(n_3535),
.B(n_1597),
.Y(n_3554)
);

BUFx6f_ASAP7_75t_L g3555 ( 
.A(n_3421),
.Y(n_3555)
);

AOI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_3460),
.A2(n_911),
.B(n_903),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_3468),
.B(n_916),
.Y(n_3557)
);

A2O1A1Ixp33_ASAP7_75t_SL g3558 ( 
.A1(n_3547),
.A2(n_1872),
.B(n_1883),
.C(n_1866),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3463),
.B(n_4),
.Y(n_3559)
);

AOI222xp33_ASAP7_75t_L g3560 ( 
.A1(n_3357),
.A2(n_11),
.B1(n_15),
.B2(n_9),
.C1(n_10),
.C2(n_14),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3352),
.Y(n_3561)
);

OR2x2_ASAP7_75t_L g3562 ( 
.A(n_3346),
.B(n_11),
.Y(n_3562)
);

OAI221xp5_ASAP7_75t_L g3563 ( 
.A1(n_3485),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.C(n_18),
.Y(n_3563)
);

BUFx3_ASAP7_75t_L g3564 ( 
.A(n_3434),
.Y(n_3564)
);

INVx3_ASAP7_75t_L g3565 ( 
.A(n_3386),
.Y(n_3565)
);

CKINVDCx8_ASAP7_75t_R g3566 ( 
.A(n_3373),
.Y(n_3566)
);

AOI22xp33_ASAP7_75t_L g3567 ( 
.A1(n_3533),
.A2(n_1385),
.B1(n_1367),
.B2(n_1872),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3352),
.Y(n_3568)
);

AND2x4_ASAP7_75t_L g3569 ( 
.A(n_3373),
.B(n_285),
.Y(n_3569)
);

INVx2_ASAP7_75t_L g3570 ( 
.A(n_3361),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3362),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3362),
.Y(n_3572)
);

INVx3_ASAP7_75t_L g3573 ( 
.A(n_3386),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3378),
.Y(n_3574)
);

AND2x2_ASAP7_75t_L g3575 ( 
.A(n_3425),
.B(n_16),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3378),
.Y(n_3576)
);

A2O1A1Ixp33_ASAP7_75t_L g3577 ( 
.A1(n_3456),
.A2(n_22),
.B(n_19),
.C(n_21),
.Y(n_3577)
);

INVx2_ASAP7_75t_SL g3578 ( 
.A(n_3421),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3451),
.B(n_19),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3380),
.Y(n_3580)
);

OAI321xp33_ASAP7_75t_L g3581 ( 
.A1(n_3505),
.A2(n_23),
.A3(n_26),
.B1(n_21),
.B2(n_22),
.C(n_24),
.Y(n_3581)
);

NOR2xp33_ASAP7_75t_R g3582 ( 
.A(n_3532),
.B(n_3526),
.Y(n_3582)
);

O2A1O1Ixp5_ASAP7_75t_SL g3583 ( 
.A1(n_3392),
.A2(n_1883),
.B(n_1891),
.C(n_1872),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3380),
.Y(n_3584)
);

AOI22xp33_ASAP7_75t_L g3585 ( 
.A1(n_3528),
.A2(n_1385),
.B1(n_1367),
.B2(n_1883),
.Y(n_3585)
);

OA21x2_ASAP7_75t_L g3586 ( 
.A1(n_3471),
.A2(n_23),
.B(n_26),
.Y(n_3586)
);

BUFx12f_ASAP7_75t_L g3587 ( 
.A(n_3360),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3419),
.Y(n_3588)
);

AND2x2_ASAP7_75t_L g3589 ( 
.A(n_3423),
.B(n_27),
.Y(n_3589)
);

OR2x2_ASAP7_75t_L g3590 ( 
.A(n_3419),
.B(n_27),
.Y(n_3590)
);

AND2x2_ASAP7_75t_L g3591 ( 
.A(n_3423),
.B(n_29),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3436),
.B(n_3530),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3370),
.B(n_29),
.Y(n_3593)
);

INVx3_ASAP7_75t_L g3594 ( 
.A(n_3423),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_3384),
.B(n_3522),
.Y(n_3595)
);

INVx1_ASAP7_75t_SL g3596 ( 
.A(n_3371),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3414),
.A2(n_1939),
.B(n_1912),
.Y(n_3597)
);

INVx2_ASAP7_75t_L g3598 ( 
.A(n_3420),
.Y(n_3598)
);

BUFx6f_ASAP7_75t_L g3599 ( 
.A(n_3421),
.Y(n_3599)
);

AND2x4_ASAP7_75t_L g3600 ( 
.A(n_3373),
.B(n_290),
.Y(n_3600)
);

INVx2_ASAP7_75t_L g3601 ( 
.A(n_3420),
.Y(n_3601)
);

OR2x6_ASAP7_75t_L g3602 ( 
.A(n_3535),
.B(n_1419),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3522),
.B(n_30),
.Y(n_3603)
);

OAI22xp5_ASAP7_75t_L g3604 ( 
.A1(n_3375),
.A2(n_1939),
.B1(n_1912),
.B2(n_1932),
.Y(n_3604)
);

BUFx3_ASAP7_75t_L g3605 ( 
.A(n_3354),
.Y(n_3605)
);

O2A1O1Ixp33_ASAP7_75t_L g3606 ( 
.A1(n_3431),
.A2(n_35),
.B(n_31),
.C(n_33),
.Y(n_3606)
);

AOI221x1_ASAP7_75t_L g3607 ( 
.A1(n_3410),
.A2(n_37),
.B1(n_31),
.B2(n_35),
.C(n_40),
.Y(n_3607)
);

INVx2_ASAP7_75t_L g3608 ( 
.A(n_3377),
.Y(n_3608)
);

INVx8_ASAP7_75t_L g3609 ( 
.A(n_3399),
.Y(n_3609)
);

INVx2_ASAP7_75t_L g3610 ( 
.A(n_3395),
.Y(n_3610)
);

AND2x2_ASAP7_75t_L g3611 ( 
.A(n_3512),
.B(n_37),
.Y(n_3611)
);

NOR2xp67_ASAP7_75t_L g3612 ( 
.A(n_3428),
.B(n_41),
.Y(n_3612)
);

AOI21xp5_ASAP7_75t_L g3613 ( 
.A1(n_3353),
.A2(n_1939),
.B(n_1912),
.Y(n_3613)
);

AOI22xp33_ASAP7_75t_L g3614 ( 
.A1(n_3427),
.A2(n_1891),
.B1(n_1932),
.B2(n_1414),
.Y(n_3614)
);

AOI22xp33_ASAP7_75t_L g3615 ( 
.A1(n_3440),
.A2(n_1891),
.B1(n_1932),
.B2(n_1414),
.Y(n_3615)
);

NOR2xp33_ASAP7_75t_SL g3616 ( 
.A(n_3486),
.B(n_3397),
.Y(n_3616)
);

BUFx12f_ASAP7_75t_L g3617 ( 
.A(n_3343),
.Y(n_3617)
);

OR2x2_ASAP7_75t_L g3618 ( 
.A(n_3347),
.B(n_42),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_3503),
.B(n_44),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3484),
.Y(n_3620)
);

OA21x2_ASAP7_75t_L g3621 ( 
.A1(n_3349),
.A2(n_44),
.B(n_45),
.Y(n_3621)
);

OR2x2_ASAP7_75t_L g3622 ( 
.A(n_3503),
.B(n_3429),
.Y(n_3622)
);

A2O1A1Ixp33_ASAP7_75t_L g3623 ( 
.A1(n_3456),
.A2(n_3374),
.B(n_3518),
.C(n_3474),
.Y(n_3623)
);

CKINVDCx11_ASAP7_75t_R g3624 ( 
.A(n_3372),
.Y(n_3624)
);

AND2x6_ASAP7_75t_L g3625 ( 
.A(n_3478),
.B(n_1673),
.Y(n_3625)
);

AND2x4_ASAP7_75t_L g3626 ( 
.A(n_3484),
.B(n_292),
.Y(n_3626)
);

AOI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_3458),
.A2(n_3443),
.B(n_3470),
.Y(n_3627)
);

AOI21xp5_ASAP7_75t_L g3628 ( 
.A1(n_3443),
.A2(n_1685),
.B(n_1673),
.Y(n_3628)
);

INVx2_ASAP7_75t_L g3629 ( 
.A(n_3408),
.Y(n_3629)
);

INVx2_ASAP7_75t_SL g3630 ( 
.A(n_3393),
.Y(n_3630)
);

INVx2_ASAP7_75t_L g3631 ( 
.A(n_3489),
.Y(n_3631)
);

AND2x4_ASAP7_75t_L g3632 ( 
.A(n_3397),
.B(n_293),
.Y(n_3632)
);

NOR2xp33_ASAP7_75t_L g3633 ( 
.A(n_3439),
.B(n_45),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3388),
.B(n_46),
.Y(n_3634)
);

AND2x2_ASAP7_75t_L g3635 ( 
.A(n_3364),
.B(n_46),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3540),
.B(n_47),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3429),
.Y(n_3637)
);

A2O1A1Ixp33_ASAP7_75t_L g3638 ( 
.A1(n_3374),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_3638)
);

OAI22xp5_ASAP7_75t_SL g3639 ( 
.A1(n_3457),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_3639)
);

OR2x2_ASAP7_75t_L g3640 ( 
.A(n_3464),
.B(n_51),
.Y(n_3640)
);

AOI21xp5_ASAP7_75t_L g3641 ( 
.A1(n_3470),
.A2(n_1685),
.B(n_1673),
.Y(n_3641)
);

INVx1_ASAP7_75t_SL g3642 ( 
.A(n_3551),
.Y(n_3642)
);

INVxp67_ASAP7_75t_L g3643 ( 
.A(n_3356),
.Y(n_3643)
);

INVx3_ASAP7_75t_L g3644 ( 
.A(n_3351),
.Y(n_3644)
);

AND2x2_ASAP7_75t_L g3645 ( 
.A(n_3491),
.B(n_52),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3464),
.Y(n_3646)
);

INVx2_ASAP7_75t_L g3647 ( 
.A(n_3482),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3450),
.Y(n_3648)
);

AOI21xp33_ASAP7_75t_SL g3649 ( 
.A1(n_3457),
.A2(n_52),
.B(n_53),
.Y(n_3649)
);

OAI22xp5_ASAP7_75t_L g3650 ( 
.A1(n_3518),
.A2(n_3452),
.B1(n_3549),
.B2(n_3390),
.Y(n_3650)
);

OAI22xp5_ASAP7_75t_L g3651 ( 
.A1(n_3452),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_3651)
);

INVx2_ASAP7_75t_SL g3652 ( 
.A(n_3379),
.Y(n_3652)
);

AND2x4_ASAP7_75t_L g3653 ( 
.A(n_3497),
.B(n_296),
.Y(n_3653)
);

HB1xp67_ASAP7_75t_L g3654 ( 
.A(n_3351),
.Y(n_3654)
);

BUFx2_ASAP7_75t_L g3655 ( 
.A(n_3491),
.Y(n_3655)
);

BUFx6f_ASAP7_75t_L g3656 ( 
.A(n_3379),
.Y(n_3656)
);

AOI21xp5_ASAP7_75t_L g3657 ( 
.A1(n_3442),
.A2(n_1685),
.B(n_1673),
.Y(n_3657)
);

NOR2xp67_ASAP7_75t_L g3658 ( 
.A(n_3381),
.B(n_3382),
.Y(n_3658)
);

OAI22xp5_ASAP7_75t_L g3659 ( 
.A1(n_3398),
.A2(n_59),
.B1(n_55),
.B2(n_57),
.Y(n_3659)
);

A2O1A1Ixp33_ASAP7_75t_L g3660 ( 
.A1(n_3544),
.A2(n_60),
.B(n_57),
.C(n_59),
.Y(n_3660)
);

AOI22xp33_ASAP7_75t_L g3661 ( 
.A1(n_3481),
.A2(n_1414),
.B1(n_1455),
.B2(n_1452),
.Y(n_3661)
);

INVx2_ASAP7_75t_L g3662 ( 
.A(n_3546),
.Y(n_3662)
);

OAI21xp5_ASAP7_75t_L g3663 ( 
.A1(n_3536),
.A2(n_1414),
.B(n_1309),
.Y(n_3663)
);

AND2x4_ASAP7_75t_L g3664 ( 
.A(n_3497),
.B(n_300),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3426),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_3424),
.B(n_61),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3432),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3446),
.B(n_62),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3546),
.Y(n_3669)
);

BUFx6f_ASAP7_75t_L g3670 ( 
.A(n_3379),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3493),
.Y(n_3671)
);

BUFx6f_ASAP7_75t_L g3672 ( 
.A(n_3498),
.Y(n_3672)
);

CKINVDCx20_ASAP7_75t_R g3673 ( 
.A(n_3343),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_3394),
.Y(n_3674)
);

BUFx10_ASAP7_75t_L g3675 ( 
.A(n_3516),
.Y(n_3675)
);

AND2x2_ASAP7_75t_L g3676 ( 
.A(n_3394),
.B(n_62),
.Y(n_3676)
);

AND2x4_ASAP7_75t_L g3677 ( 
.A(n_3497),
.B(n_307),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3493),
.Y(n_3678)
);

CKINVDCx16_ASAP7_75t_R g3679 ( 
.A(n_3453),
.Y(n_3679)
);

AOI21xp33_ASAP7_75t_L g3680 ( 
.A1(n_3527),
.A2(n_64),
.B(n_65),
.Y(n_3680)
);

OR2x2_ASAP7_75t_L g3681 ( 
.A(n_3553),
.B(n_64),
.Y(n_3681)
);

INVx2_ASAP7_75t_L g3682 ( 
.A(n_3404),
.Y(n_3682)
);

AND2x6_ASAP7_75t_L g3683 ( 
.A(n_3478),
.B(n_1673),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3404),
.Y(n_3684)
);

AO22x1_ASAP7_75t_L g3685 ( 
.A1(n_3516),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_3685)
);

OR2x6_ASAP7_75t_L g3686 ( 
.A(n_3385),
.B(n_1419),
.Y(n_3686)
);

OAI21xp5_ASAP7_75t_L g3687 ( 
.A1(n_3359),
.A2(n_1414),
.B(n_1309),
.Y(n_3687)
);

OAI22xp5_ASAP7_75t_SL g3688 ( 
.A1(n_3494),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_3688)
);

INVx2_ASAP7_75t_SL g3689 ( 
.A(n_3498),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3493),
.Y(n_3690)
);

CKINVDCx5p33_ASAP7_75t_R g3691 ( 
.A(n_3348),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_3550),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3355),
.Y(n_3693)
);

OR2x2_ASAP7_75t_L g3694 ( 
.A(n_3495),
.B(n_69),
.Y(n_3694)
);

AND2x2_ASAP7_75t_L g3695 ( 
.A(n_3550),
.B(n_3498),
.Y(n_3695)
);

INVx4_ASAP7_75t_L g3696 ( 
.A(n_3461),
.Y(n_3696)
);

CKINVDCx5p33_ASAP7_75t_R g3697 ( 
.A(n_3348),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3450),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3450),
.Y(n_3699)
);

OR2x2_ASAP7_75t_L g3700 ( 
.A(n_3490),
.B(n_70),
.Y(n_3700)
);

OAI211xp5_ASAP7_75t_L g3701 ( 
.A1(n_3437),
.A2(n_75),
.B(n_72),
.C(n_74),
.Y(n_3701)
);

AND2x2_ASAP7_75t_L g3702 ( 
.A(n_3453),
.B(n_72),
.Y(n_3702)
);

AND2x2_ASAP7_75t_L g3703 ( 
.A(n_3453),
.B(n_76),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3413),
.Y(n_3704)
);

NAND2xp33_ASAP7_75t_L g3705 ( 
.A(n_3430),
.B(n_1685),
.Y(n_3705)
);

INVx3_ASAP7_75t_L g3706 ( 
.A(n_3461),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3413),
.Y(n_3707)
);

A2O1A1Ixp33_ASAP7_75t_L g3708 ( 
.A1(n_3506),
.A2(n_79),
.B(n_76),
.C(n_78),
.Y(n_3708)
);

A2O1A1Ixp33_ASAP7_75t_L g3709 ( 
.A1(n_3467),
.A2(n_82),
.B(n_78),
.C(n_80),
.Y(n_3709)
);

AOI21xp5_ASAP7_75t_L g3710 ( 
.A1(n_3455),
.A2(n_1729),
.B(n_1685),
.Y(n_3710)
);

O2A1O1Ixp33_ASAP7_75t_L g3711 ( 
.A1(n_3454),
.A2(n_85),
.B(n_80),
.C(n_84),
.Y(n_3711)
);

AOI22xp33_ASAP7_75t_L g3712 ( 
.A1(n_3509),
.A2(n_3369),
.B1(n_3417),
.B2(n_3500),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3469),
.B(n_85),
.Y(n_3713)
);

AOI21xp5_ASAP7_75t_L g3714 ( 
.A1(n_3502),
.A2(n_1731),
.B(n_1729),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3368),
.B(n_3479),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3487),
.B(n_86),
.Y(n_3716)
);

AND2x4_ASAP7_75t_L g3717 ( 
.A(n_3477),
.B(n_308),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3402),
.B(n_87),
.Y(n_3718)
);

CKINVDCx5p33_ASAP7_75t_R g3719 ( 
.A(n_3515),
.Y(n_3719)
);

BUFx3_ASAP7_75t_L g3720 ( 
.A(n_3515),
.Y(n_3720)
);

HB1xp67_ASAP7_75t_L g3721 ( 
.A(n_3541),
.Y(n_3721)
);

OA21x2_ASAP7_75t_L g3722 ( 
.A1(n_3345),
.A2(n_87),
.B(n_88),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3412),
.B(n_88),
.Y(n_3723)
);

BUFx2_ASAP7_75t_L g3724 ( 
.A(n_3477),
.Y(n_3724)
);

OAI21x1_ASAP7_75t_L g3725 ( 
.A1(n_3465),
.A2(n_1333),
.B(n_1304),
.Y(n_3725)
);

BUFx2_ASAP7_75t_L g3726 ( 
.A(n_3515),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3541),
.B(n_89),
.Y(n_3727)
);

AND2x4_ASAP7_75t_L g3728 ( 
.A(n_3543),
.B(n_312),
.Y(n_3728)
);

BUFx6f_ASAP7_75t_L g3729 ( 
.A(n_3534),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3413),
.Y(n_3730)
);

AOI22xp33_ASAP7_75t_SL g3731 ( 
.A1(n_3545),
.A2(n_93),
.B1(n_90),
.B2(n_92),
.Y(n_3731)
);

BUFx4f_ASAP7_75t_SL g3732 ( 
.A(n_3350),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3433),
.B(n_90),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3409),
.Y(n_3734)
);

BUFx2_ASAP7_75t_L g3735 ( 
.A(n_3545),
.Y(n_3735)
);

AND2x2_ASAP7_75t_L g3736 ( 
.A(n_3517),
.B(n_3435),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3409),
.Y(n_3737)
);

A2O1A1Ixp33_ASAP7_75t_L g3738 ( 
.A1(n_3538),
.A2(n_95),
.B(n_92),
.C(n_94),
.Y(n_3738)
);

AOI21xp5_ASAP7_75t_L g3739 ( 
.A1(n_3462),
.A2(n_1731),
.B(n_1729),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3409),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3524),
.B(n_94),
.Y(n_3741)
);

NAND3xp33_ASAP7_75t_L g3742 ( 
.A(n_3418),
.B(n_1455),
.C(n_1452),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3504),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3407),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3407),
.Y(n_3745)
);

AND2x4_ASAP7_75t_L g3746 ( 
.A(n_3543),
.B(n_315),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3501),
.Y(n_3747)
);

AND2x4_ASAP7_75t_L g3748 ( 
.A(n_3441),
.B(n_322),
.Y(n_3748)
);

AND2x2_ASAP7_75t_L g3749 ( 
.A(n_3517),
.B(n_96),
.Y(n_3749)
);

CKINVDCx5p33_ASAP7_75t_R g3750 ( 
.A(n_3520),
.Y(n_3750)
);

AND2x2_ASAP7_75t_L g3751 ( 
.A(n_3517),
.B(n_96),
.Y(n_3751)
);

AND2x2_ASAP7_75t_L g3752 ( 
.A(n_3514),
.B(n_98),
.Y(n_3752)
);

AO21x1_ASAP7_75t_L g3753 ( 
.A1(n_3363),
.A2(n_98),
.B(n_99),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_L g3754 ( 
.A(n_3418),
.B(n_100),
.Y(n_3754)
);

INVx4_ASAP7_75t_L g3755 ( 
.A(n_3406),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3514),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3514),
.Y(n_3757)
);

AND2x4_ASAP7_75t_L g3758 ( 
.A(n_3548),
.B(n_327),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3376),
.Y(n_3759)
);

AND2x2_ASAP7_75t_L g3760 ( 
.A(n_3537),
.B(n_100),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3459),
.B(n_101),
.Y(n_3761)
);

AOI22xp33_ASAP7_75t_L g3762 ( 
.A1(n_3519),
.A2(n_1455),
.B1(n_1459),
.B2(n_1452),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_SL g3763 ( 
.A(n_3366),
.B(n_3391),
.Y(n_3763)
);

BUFx2_ASAP7_75t_L g3764 ( 
.A(n_3507),
.Y(n_3764)
);

CKINVDCx5p33_ASAP7_75t_R g3765 ( 
.A(n_3513),
.Y(n_3765)
);

OR2x2_ASAP7_75t_L g3766 ( 
.A(n_3510),
.B(n_101),
.Y(n_3766)
);

AND2x2_ASAP7_75t_SL g3767 ( 
.A(n_3529),
.B(n_102),
.Y(n_3767)
);

A2O1A1Ixp33_ASAP7_75t_L g3768 ( 
.A1(n_3523),
.A2(n_106),
.B(n_103),
.C(n_105),
.Y(n_3768)
);

BUFx3_ASAP7_75t_L g3769 ( 
.A(n_3449),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3365),
.B(n_106),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_L g3771 ( 
.A(n_3396),
.B(n_108),
.Y(n_3771)
);

AOI21xp5_ASAP7_75t_L g3772 ( 
.A1(n_3483),
.A2(n_1731),
.B(n_1729),
.Y(n_3772)
);

OAI22xp5_ASAP7_75t_L g3773 ( 
.A1(n_3447),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_3773)
);

AOI22xp33_ASAP7_75t_SL g3774 ( 
.A1(n_3650),
.A2(n_3531),
.B1(n_3511),
.B2(n_3499),
.Y(n_3774)
);

INVx6_ASAP7_75t_L g3775 ( 
.A(n_3617),
.Y(n_3775)
);

INVx11_ASAP7_75t_L g3776 ( 
.A(n_3587),
.Y(n_3776)
);

AOI22xp33_ASAP7_75t_L g3777 ( 
.A1(n_3560),
.A2(n_3542),
.B1(n_3472),
.B2(n_3405),
.Y(n_3777)
);

BUFx6f_ASAP7_75t_L g3778 ( 
.A(n_3555),
.Y(n_3778)
);

BUFx10_ASAP7_75t_L g3779 ( 
.A(n_3656),
.Y(n_3779)
);

OAI21xp5_ASAP7_75t_L g3780 ( 
.A1(n_3623),
.A2(n_3383),
.B(n_3389),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3561),
.Y(n_3781)
);

BUFx6f_ASAP7_75t_L g3782 ( 
.A(n_3555),
.Y(n_3782)
);

AOI22xp33_ASAP7_75t_L g3783 ( 
.A1(n_3688),
.A2(n_3763),
.B1(n_3563),
.B2(n_3639),
.Y(n_3783)
);

OAI22xp33_ASAP7_75t_L g3784 ( 
.A1(n_3607),
.A2(n_3539),
.B1(n_3521),
.B2(n_3496),
.Y(n_3784)
);

AOI22xp33_ASAP7_75t_L g3785 ( 
.A1(n_3755),
.A2(n_3466),
.B1(n_3416),
.B2(n_3422),
.Y(n_3785)
);

BUFx3_ASAP7_75t_L g3786 ( 
.A(n_3609),
.Y(n_3786)
);

INVx8_ASAP7_75t_L g3787 ( 
.A(n_3609),
.Y(n_3787)
);

CKINVDCx5p33_ASAP7_75t_R g3788 ( 
.A(n_3624),
.Y(n_3788)
);

CKINVDCx6p67_ASAP7_75t_R g3789 ( 
.A(n_3673),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3561),
.Y(n_3790)
);

CKINVDCx20_ASAP7_75t_R g3791 ( 
.A(n_3582),
.Y(n_3791)
);

INVx1_ASAP7_75t_SL g3792 ( 
.A(n_3724),
.Y(n_3792)
);

AOI22xp33_ASAP7_75t_L g3793 ( 
.A1(n_3755),
.A2(n_3444),
.B1(n_3438),
.B2(n_3488),
.Y(n_3793)
);

OR2x2_ASAP7_75t_L g3794 ( 
.A(n_3631),
.B(n_3344),
.Y(n_3794)
);

BUFx6f_ASAP7_75t_L g3795 ( 
.A(n_3555),
.Y(n_3795)
);

INVx2_ASAP7_75t_L g3796 ( 
.A(n_3662),
.Y(n_3796)
);

AOI22xp33_ASAP7_75t_L g3797 ( 
.A1(n_3753),
.A2(n_3492),
.B1(n_3445),
.B2(n_3473),
.Y(n_3797)
);

AOI22xp33_ASAP7_75t_SL g3798 ( 
.A1(n_3701),
.A2(n_3552),
.B1(n_3358),
.B2(n_3480),
.Y(n_3798)
);

AOI22xp33_ASAP7_75t_L g3799 ( 
.A1(n_3732),
.A2(n_3448),
.B1(n_3475),
.B2(n_3476),
.Y(n_3799)
);

INVx2_ASAP7_75t_L g3800 ( 
.A(n_3669),
.Y(n_3800)
);

AOI22xp33_ASAP7_75t_L g3801 ( 
.A1(n_3651),
.A2(n_3712),
.B1(n_3658),
.B2(n_3731),
.Y(n_3801)
);

AOI22xp33_ASAP7_75t_L g3802 ( 
.A1(n_3752),
.A2(n_3415),
.B1(n_3400),
.B2(n_3401),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3595),
.B(n_109),
.Y(n_3803)
);

OAI21xp5_ASAP7_75t_SL g3804 ( 
.A1(n_3711),
.A2(n_110),
.B(n_112),
.Y(n_3804)
);

INVx2_ASAP7_75t_SL g3805 ( 
.A(n_3599),
.Y(n_3805)
);

BUFx4f_ASAP7_75t_SL g3806 ( 
.A(n_3596),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3568),
.Y(n_3807)
);

OAI21xp5_ASAP7_75t_L g3808 ( 
.A1(n_3709),
.A2(n_3367),
.B(n_3403),
.Y(n_3808)
);

BUFx8_ASAP7_75t_SL g3809 ( 
.A(n_3691),
.Y(n_3809)
);

AOI22xp33_ASAP7_75t_L g3810 ( 
.A1(n_3659),
.A2(n_3387),
.B1(n_3411),
.B2(n_1455),
.Y(n_3810)
);

INVx5_ASAP7_75t_L g3811 ( 
.A(n_3554),
.Y(n_3811)
);

INVx2_ASAP7_75t_L g3812 ( 
.A(n_3576),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3571),
.Y(n_3813)
);

CKINVDCx11_ASAP7_75t_R g3814 ( 
.A(n_3566),
.Y(n_3814)
);

AOI22xp33_ASAP7_75t_L g3815 ( 
.A1(n_3680),
.A2(n_1459),
.B1(n_1452),
.B2(n_1333),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_L g3816 ( 
.A(n_3592),
.B(n_112),
.Y(n_3816)
);

OR2x2_ASAP7_75t_L g3817 ( 
.A(n_3622),
.B(n_3496),
.Y(n_3817)
);

CKINVDCx11_ASAP7_75t_R g3818 ( 
.A(n_3656),
.Y(n_3818)
);

AOI22xp5_ASAP7_75t_L g3819 ( 
.A1(n_3708),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3647),
.B(n_114),
.Y(n_3820)
);

AOI22xp33_ASAP7_75t_L g3821 ( 
.A1(n_3761),
.A2(n_1459),
.B1(n_1362),
.B2(n_1390),
.Y(n_3821)
);

OAI22xp5_ASAP7_75t_SL g3822 ( 
.A1(n_3642),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_3822)
);

AOI22xp33_ASAP7_75t_L g3823 ( 
.A1(n_3705),
.A2(n_1459),
.B1(n_1362),
.B2(n_1390),
.Y(n_3823)
);

CKINVDCx11_ASAP7_75t_R g3824 ( 
.A(n_3656),
.Y(n_3824)
);

AOI22xp33_ASAP7_75t_SL g3825 ( 
.A1(n_3616),
.A2(n_119),
.B1(n_116),
.B2(n_118),
.Y(n_3825)
);

INVx1_ASAP7_75t_SL g3826 ( 
.A(n_3654),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3572),
.Y(n_3827)
);

INVx2_ASAP7_75t_L g3828 ( 
.A(n_3598),
.Y(n_3828)
);

OAI21xp5_ASAP7_75t_SL g3829 ( 
.A1(n_3649),
.A2(n_118),
.B(n_121),
.Y(n_3829)
);

CKINVDCx11_ASAP7_75t_R g3830 ( 
.A(n_3670),
.Y(n_3830)
);

AOI22xp33_ASAP7_75t_L g3831 ( 
.A1(n_3736),
.A2(n_1304),
.B1(n_126),
.B2(n_122),
.Y(n_3831)
);

AOI22xp33_ASAP7_75t_L g3832 ( 
.A1(n_3735),
.A2(n_127),
.B1(n_123),
.B2(n_126),
.Y(n_3832)
);

CKINVDCx5p33_ASAP7_75t_R g3833 ( 
.A(n_3599),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_L g3834 ( 
.A(n_3743),
.B(n_127),
.Y(n_3834)
);

CKINVDCx11_ASAP7_75t_R g3835 ( 
.A(n_3670),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3574),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3580),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3584),
.Y(n_3838)
);

INVx3_ASAP7_75t_L g3839 ( 
.A(n_3605),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3601),
.Y(n_3840)
);

INVx4_ASAP7_75t_SL g3841 ( 
.A(n_3670),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_3747),
.B(n_128),
.Y(n_3842)
);

INVx8_ASAP7_75t_L g3843 ( 
.A(n_3569),
.Y(n_3843)
);

BUFx12f_ASAP7_75t_L g3844 ( 
.A(n_3652),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3588),
.Y(n_3845)
);

OAI22xp33_ASAP7_75t_L g3846 ( 
.A1(n_3581),
.A2(n_3496),
.B1(n_3508),
.B2(n_3525),
.Y(n_3846)
);

AOI22xp33_ASAP7_75t_SL g3847 ( 
.A1(n_3749),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_3847)
);

BUFx2_ASAP7_75t_L g3848 ( 
.A(n_3565),
.Y(n_3848)
);

INVx2_ASAP7_75t_SL g3849 ( 
.A(n_3599),
.Y(n_3849)
);

INVx2_ASAP7_75t_L g3850 ( 
.A(n_3620),
.Y(n_3850)
);

OAI22xp5_ASAP7_75t_L g3851 ( 
.A1(n_3638),
.A2(n_3525),
.B1(n_3508),
.B2(n_133),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3637),
.Y(n_3852)
);

BUFx6f_ASAP7_75t_L g3853 ( 
.A(n_3672),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3570),
.Y(n_3854)
);

OAI22xp33_ASAP7_75t_L g3855 ( 
.A1(n_3754),
.A2(n_3508),
.B1(n_3525),
.B2(n_133),
.Y(n_3855)
);

INVx4_ASAP7_75t_L g3856 ( 
.A(n_3729),
.Y(n_3856)
);

INVx2_ASAP7_75t_L g3857 ( 
.A(n_3608),
.Y(n_3857)
);

INVx4_ASAP7_75t_L g3858 ( 
.A(n_3729),
.Y(n_3858)
);

INVx6_ASAP7_75t_L g3859 ( 
.A(n_3675),
.Y(n_3859)
);

BUFx12f_ASAP7_75t_L g3860 ( 
.A(n_3697),
.Y(n_3860)
);

AOI22xp33_ASAP7_75t_SL g3861 ( 
.A1(n_3751),
.A2(n_134),
.B1(n_131),
.B2(n_132),
.Y(n_3861)
);

AOI21xp5_ASAP7_75t_L g3862 ( 
.A1(n_3714),
.A2(n_1731),
.B(n_1729),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3637),
.Y(n_3863)
);

AND2x2_ASAP7_75t_L g3864 ( 
.A(n_3565),
.B(n_135),
.Y(n_3864)
);

AOI22xp33_ASAP7_75t_L g3865 ( 
.A1(n_3643),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3646),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3646),
.Y(n_3867)
);

OAI22xp5_ASAP7_75t_L g3868 ( 
.A1(n_3660),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3610),
.Y(n_3869)
);

INVx1_ASAP7_75t_SL g3870 ( 
.A(n_3655),
.Y(n_3870)
);

AOI22xp33_ASAP7_75t_L g3871 ( 
.A1(n_3729),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_3871)
);

AOI22xp5_ASAP7_75t_L g3872 ( 
.A1(n_3715),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_3872)
);

INVx2_ASAP7_75t_R g3873 ( 
.A(n_3693),
.Y(n_3873)
);

INVx1_ASAP7_75t_SL g3874 ( 
.A(n_3750),
.Y(n_3874)
);

INVx4_ASAP7_75t_SL g3875 ( 
.A(n_3625),
.Y(n_3875)
);

AOI22xp33_ASAP7_75t_L g3876 ( 
.A1(n_3773),
.A2(n_147),
.B1(n_143),
.B2(n_146),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3629),
.Y(n_3877)
);

OAI22xp5_ASAP7_75t_L g3878 ( 
.A1(n_3577),
.A2(n_150),
.B1(n_146),
.B2(n_149),
.Y(n_3878)
);

AOI22xp33_ASAP7_75t_L g3879 ( 
.A1(n_3665),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_3879)
);

OAI22xp5_ASAP7_75t_L g3880 ( 
.A1(n_3738),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3667),
.Y(n_3881)
);

OAI22xp5_ASAP7_75t_L g3882 ( 
.A1(n_3767),
.A2(n_156),
.B1(n_153),
.B2(n_154),
.Y(n_3882)
);

BUFx3_ASAP7_75t_L g3883 ( 
.A(n_3564),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3727),
.Y(n_3884)
);

AND2x2_ASAP7_75t_L g3885 ( 
.A(n_3573),
.B(n_156),
.Y(n_3885)
);

BUFx2_ASAP7_75t_L g3886 ( 
.A(n_3573),
.Y(n_3886)
);

AOI22xp33_ASAP7_75t_SL g3887 ( 
.A1(n_3586),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_3887)
);

INVx2_ASAP7_75t_L g3888 ( 
.A(n_3674),
.Y(n_3888)
);

BUFx4f_ASAP7_75t_SL g3889 ( 
.A(n_3630),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3682),
.Y(n_3890)
);

AOI22xp33_ASAP7_75t_L g3891 ( 
.A1(n_3765),
.A2(n_3748),
.B1(n_3626),
.B2(n_3633),
.Y(n_3891)
);

AOI22xp33_ASAP7_75t_SL g3892 ( 
.A1(n_3586),
.A2(n_3678),
.B1(n_3690),
.B2(n_3671),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_3684),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3692),
.Y(n_3894)
);

AND2x2_ASAP7_75t_L g3895 ( 
.A(n_3695),
.B(n_157),
.Y(n_3895)
);

INVx6_ASAP7_75t_L g3896 ( 
.A(n_3675),
.Y(n_3896)
);

BUFx6f_ASAP7_75t_L g3897 ( 
.A(n_3672),
.Y(n_3897)
);

AOI22xp33_ASAP7_75t_L g3898 ( 
.A1(n_3748),
.A2(n_162),
.B1(n_159),
.B2(n_161),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3648),
.Y(n_3899)
);

AOI22xp33_ASAP7_75t_L g3900 ( 
.A1(n_3626),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_L g3901 ( 
.A(n_3618),
.B(n_166),
.Y(n_3901)
);

AOI22xp5_ASAP7_75t_L g3902 ( 
.A1(n_3685),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.Y(n_3902)
);

AND2x4_ASAP7_75t_L g3903 ( 
.A(n_3706),
.B(n_168),
.Y(n_3903)
);

INVx2_ASAP7_75t_L g3904 ( 
.A(n_3706),
.Y(n_3904)
);

INVx1_ASAP7_75t_SL g3905 ( 
.A(n_3644),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3644),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_3559),
.B(n_170),
.Y(n_3907)
);

BUFx2_ASAP7_75t_L g3908 ( 
.A(n_3594),
.Y(n_3908)
);

OAI22xp5_ASAP7_75t_L g3909 ( 
.A1(n_3606),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_3909)
);

CKINVDCx20_ASAP7_75t_R g3910 ( 
.A(n_3679),
.Y(n_3910)
);

AND2x2_ASAP7_75t_L g3911 ( 
.A(n_3594),
.B(n_171),
.Y(n_3911)
);

NAND2x1p5_ASAP7_75t_L g3912 ( 
.A(n_3653),
.B(n_1419),
.Y(n_3912)
);

AOI21xp5_ASAP7_75t_L g3913 ( 
.A1(n_3663),
.A2(n_1757),
.B(n_1731),
.Y(n_3913)
);

AOI22xp33_ASAP7_75t_SL g3914 ( 
.A1(n_3770),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3648),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3698),
.Y(n_3916)
);

HB1xp67_ASAP7_75t_L g3917 ( 
.A(n_3721),
.Y(n_3917)
);

CKINVDCx20_ASAP7_75t_R g3918 ( 
.A(n_3719),
.Y(n_3918)
);

BUFx4f_ASAP7_75t_SL g3919 ( 
.A(n_3578),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3696),
.Y(n_3920)
);

HB1xp67_ASAP7_75t_L g3921 ( 
.A(n_3756),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3698),
.Y(n_3922)
);

BUFx12f_ASAP7_75t_L g3923 ( 
.A(n_3589),
.Y(n_3923)
);

BUFx12f_ASAP7_75t_L g3924 ( 
.A(n_3591),
.Y(n_3924)
);

AOI22xp33_ASAP7_75t_L g3925 ( 
.A1(n_3634),
.A2(n_3635),
.B1(n_3713),
.B2(n_3668),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3699),
.Y(n_3926)
);

AOI22xp33_ASAP7_75t_L g3927 ( 
.A1(n_3718),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_3927)
);

AOI22xp33_ASAP7_75t_L g3928 ( 
.A1(n_3723),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_3928)
);

INVx6_ASAP7_75t_L g3929 ( 
.A(n_3672),
.Y(n_3929)
);

AOI22xp33_ASAP7_75t_L g3930 ( 
.A1(n_3733),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_3930)
);

CKINVDCx11_ASAP7_75t_R g3931 ( 
.A(n_3720),
.Y(n_3931)
);

AND2x4_ASAP7_75t_L g3932 ( 
.A(n_3696),
.B(n_181),
.Y(n_3932)
);

CKINVDCx11_ASAP7_75t_R g3933 ( 
.A(n_3726),
.Y(n_3933)
);

BUFx3_ASAP7_75t_L g3934 ( 
.A(n_3689),
.Y(n_3934)
);

INVxp67_ASAP7_75t_L g3935 ( 
.A(n_3636),
.Y(n_3935)
);

INVx2_ASAP7_75t_L g3936 ( 
.A(n_3590),
.Y(n_3936)
);

AOI22xp33_ASAP7_75t_SL g3937 ( 
.A1(n_3771),
.A2(n_182),
.B1(n_184),
.B2(n_186),
.Y(n_3937)
);

AOI22xp33_ASAP7_75t_SL g3938 ( 
.A1(n_3556),
.A2(n_184),
.B1(n_187),
.B2(n_188),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_3603),
.B(n_3611),
.Y(n_3939)
);

CKINVDCx5p33_ASAP7_75t_R g3940 ( 
.A(n_3575),
.Y(n_3940)
);

CKINVDCx5p33_ASAP7_75t_R g3941 ( 
.A(n_3702),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3699),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_L g3943 ( 
.A(n_3619),
.B(n_187),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3704),
.Y(n_3944)
);

BUFx2_ASAP7_75t_L g3945 ( 
.A(n_3602),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3884),
.B(n_3757),
.Y(n_3946)
);

NOR3xp33_ASAP7_75t_L g3947 ( 
.A(n_3804),
.B(n_3716),
.C(n_3666),
.Y(n_3947)
);

OA21x2_ASAP7_75t_L g3948 ( 
.A1(n_3899),
.A2(n_3707),
.B(n_3704),
.Y(n_3948)
);

INVx2_ASAP7_75t_SL g3949 ( 
.A(n_3883),
.Y(n_3949)
);

O2A1O1Ixp33_ASAP7_75t_L g3950 ( 
.A1(n_3804),
.A2(n_3640),
.B(n_3741),
.C(n_3593),
.Y(n_3950)
);

O2A1O1Ixp33_ASAP7_75t_L g3951 ( 
.A1(n_3829),
.A2(n_3768),
.B(n_3694),
.C(n_3579),
.Y(n_3951)
);

AND2x2_ASAP7_75t_L g3952 ( 
.A(n_3848),
.B(n_3764),
.Y(n_3952)
);

AOI21xp5_ASAP7_75t_SL g3953 ( 
.A1(n_3780),
.A2(n_3664),
.B(n_3653),
.Y(n_3953)
);

A2O1A1Ixp33_ASAP7_75t_L g3954 ( 
.A1(n_3829),
.A2(n_3612),
.B(n_3562),
.C(n_3627),
.Y(n_3954)
);

HB1xp67_ASAP7_75t_L g3955 ( 
.A(n_3917),
.Y(n_3955)
);

O2A1O1Ixp33_ASAP7_75t_L g3956 ( 
.A1(n_3868),
.A2(n_3878),
.B(n_3882),
.C(n_3880),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3781),
.Y(n_3957)
);

AND2x2_ASAP7_75t_L g3958 ( 
.A(n_3886),
.B(n_3769),
.Y(n_3958)
);

OA21x2_ASAP7_75t_L g3959 ( 
.A1(n_3915),
.A2(n_3707),
.B(n_3730),
.Y(n_3959)
);

O2A1O1Ixp33_ASAP7_75t_L g3960 ( 
.A1(n_3783),
.A2(n_3909),
.B(n_3801),
.C(n_3907),
.Y(n_3960)
);

NOR2xp67_ASAP7_75t_L g3961 ( 
.A(n_3856),
.B(n_3734),
.Y(n_3961)
);

CKINVDCx20_ASAP7_75t_R g3962 ( 
.A(n_3791),
.Y(n_3962)
);

INVx3_ASAP7_75t_L g3963 ( 
.A(n_3859),
.Y(n_3963)
);

OR2x2_ASAP7_75t_L g3964 ( 
.A(n_3826),
.B(n_3744),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3790),
.Y(n_3965)
);

AOI21xp5_ASAP7_75t_SL g3966 ( 
.A1(n_3902),
.A2(n_3677),
.B(n_3664),
.Y(n_3966)
);

OA21x2_ASAP7_75t_L g3967 ( 
.A1(n_3916),
.A2(n_3740),
.B(n_3737),
.Y(n_3967)
);

OR2x2_ASAP7_75t_L g3968 ( 
.A(n_3826),
.B(n_3745),
.Y(n_3968)
);

INVx2_ASAP7_75t_L g3969 ( 
.A(n_3796),
.Y(n_3969)
);

O2A1O1Ixp5_ASAP7_75t_L g3970 ( 
.A1(n_3851),
.A2(n_3557),
.B(n_3758),
.C(n_3760),
.Y(n_3970)
);

AND2x2_ASAP7_75t_L g3971 ( 
.A(n_3870),
.B(n_3703),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_L g3972 ( 
.A(n_3936),
.B(n_3766),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3807),
.Y(n_3973)
);

AND2x4_ASAP7_75t_L g3974 ( 
.A(n_3920),
.B(n_3856),
.Y(n_3974)
);

OA21x2_ASAP7_75t_L g3975 ( 
.A1(n_3922),
.A2(n_3772),
.B(n_3641),
.Y(n_3975)
);

AOI31xp33_ASAP7_75t_L g3976 ( 
.A1(n_3847),
.A2(n_3700),
.A3(n_3681),
.B(n_3600),
.Y(n_3976)
);

OAI22xp5_ASAP7_75t_L g3977 ( 
.A1(n_3819),
.A2(n_3554),
.B1(n_3686),
.B2(n_3602),
.Y(n_3977)
);

A2O1A1Ixp33_ASAP7_75t_L g3978 ( 
.A1(n_3819),
.A2(n_3569),
.B(n_3600),
.C(n_3632),
.Y(n_3978)
);

AND2x2_ASAP7_75t_L g3979 ( 
.A(n_3870),
.B(n_3621),
.Y(n_3979)
);

AND2x6_ASAP7_75t_L g3980 ( 
.A(n_3902),
.B(n_3677),
.Y(n_3980)
);

OAI22xp5_ASAP7_75t_L g3981 ( 
.A1(n_3872),
.A2(n_3661),
.B1(n_3621),
.B2(n_3722),
.Y(n_3981)
);

OAI22xp5_ASAP7_75t_L g3982 ( 
.A1(n_3872),
.A2(n_3722),
.B1(n_3686),
.B2(n_3742),
.Y(n_3982)
);

AOI21xp5_ASAP7_75t_L g3983 ( 
.A1(n_3913),
.A2(n_3558),
.B(n_3710),
.Y(n_3983)
);

INVx2_ASAP7_75t_L g3984 ( 
.A(n_3800),
.Y(n_3984)
);

AOI21xp5_ASAP7_75t_L g3985 ( 
.A1(n_3777),
.A2(n_3657),
.B(n_3628),
.Y(n_3985)
);

AND2x2_ASAP7_75t_L g3986 ( 
.A(n_3792),
.B(n_3676),
.Y(n_3986)
);

OAI22xp5_ASAP7_75t_L g3987 ( 
.A1(n_3887),
.A2(n_3728),
.B1(n_3746),
.B2(n_3758),
.Y(n_3987)
);

AND2x2_ASAP7_75t_L g3988 ( 
.A(n_3792),
.B(n_3645),
.Y(n_3988)
);

AND2x2_ASAP7_75t_L g3989 ( 
.A(n_3839),
.B(n_3759),
.Y(n_3989)
);

OA21x2_ASAP7_75t_L g3990 ( 
.A1(n_3926),
.A2(n_3725),
.B(n_3613),
.Y(n_3990)
);

NOR2x1_ASAP7_75t_SL g3991 ( 
.A(n_3858),
.B(n_3604),
.Y(n_3991)
);

OR2x2_ASAP7_75t_L g3992 ( 
.A(n_3794),
.B(n_3845),
.Y(n_3992)
);

O2A1O1Ixp5_ASAP7_75t_L g3993 ( 
.A1(n_3855),
.A2(n_3728),
.B(n_3746),
.C(n_3632),
.Y(n_3993)
);

INVx6_ASAP7_75t_L g3994 ( 
.A(n_3860),
.Y(n_3994)
);

OA21x2_ASAP7_75t_L g3995 ( 
.A1(n_3942),
.A2(n_3739),
.B(n_3687),
.Y(n_3995)
);

OA21x2_ASAP7_75t_L g3996 ( 
.A1(n_3944),
.A2(n_3597),
.B(n_3762),
.Y(n_3996)
);

BUFx8_ASAP7_75t_SL g3997 ( 
.A(n_3809),
.Y(n_3997)
);

AOI21xp5_ASAP7_75t_L g3998 ( 
.A1(n_3862),
.A2(n_3784),
.B(n_3808),
.Y(n_3998)
);

BUFx6f_ASAP7_75t_L g3999 ( 
.A(n_3818),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3869),
.B(n_3583),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_3877),
.B(n_3717),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3890),
.B(n_3717),
.Y(n_4002)
);

BUFx12f_ASAP7_75t_L g4003 ( 
.A(n_3788),
.Y(n_4003)
);

BUFx3_ASAP7_75t_L g4004 ( 
.A(n_3918),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_3893),
.B(n_3894),
.Y(n_4005)
);

HB1xp67_ASAP7_75t_L g4006 ( 
.A(n_3905),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3813),
.Y(n_4007)
);

CKINVDCx20_ASAP7_75t_R g4008 ( 
.A(n_3789),
.Y(n_4008)
);

OA21x2_ASAP7_75t_L g4009 ( 
.A1(n_3852),
.A2(n_3614),
.B(n_3567),
.Y(n_4009)
);

OAI22xp5_ASAP7_75t_L g4010 ( 
.A1(n_3891),
.A2(n_3615),
.B1(n_3585),
.B2(n_3683),
.Y(n_4010)
);

O2A1O1Ixp5_ASAP7_75t_L g4011 ( 
.A1(n_3932),
.A2(n_189),
.B(n_190),
.C(n_191),
.Y(n_4011)
);

OR2x2_ASAP7_75t_L g4012 ( 
.A(n_3850),
.B(n_189),
.Y(n_4012)
);

AND2x2_ASAP7_75t_L g4013 ( 
.A(n_3839),
.B(n_3625),
.Y(n_4013)
);

AOI21x1_ASAP7_75t_SL g4014 ( 
.A1(n_3932),
.A2(n_191),
.B(n_194),
.Y(n_4014)
);

AOI21xp5_ASAP7_75t_SL g4015 ( 
.A1(n_3912),
.A2(n_3683),
.B(n_3625),
.Y(n_4015)
);

AND2x2_ASAP7_75t_L g4016 ( 
.A(n_3908),
.B(n_3625),
.Y(n_4016)
);

OR2x2_ASAP7_75t_L g4017 ( 
.A(n_3812),
.B(n_194),
.Y(n_4017)
);

OR2x2_ASAP7_75t_L g4018 ( 
.A(n_3828),
.B(n_195),
.Y(n_4018)
);

INVx3_ASAP7_75t_L g4019 ( 
.A(n_3859),
.Y(n_4019)
);

O2A1O1Ixp33_ASAP7_75t_L g4020 ( 
.A1(n_3935),
.A2(n_195),
.B(n_196),
.C(n_197),
.Y(n_4020)
);

OA21x2_ASAP7_75t_L g4021 ( 
.A1(n_3863),
.A2(n_3683),
.B(n_198),
.Y(n_4021)
);

AND2x2_ASAP7_75t_L g4022 ( 
.A(n_3858),
.B(n_3683),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_3854),
.B(n_3857),
.Y(n_4023)
);

AOI21xp5_ASAP7_75t_SL g4024 ( 
.A1(n_3903),
.A2(n_198),
.B(n_199),
.Y(n_4024)
);

AND2x2_ASAP7_75t_L g4025 ( 
.A(n_3905),
.B(n_199),
.Y(n_4025)
);

CKINVDCx20_ASAP7_75t_R g4026 ( 
.A(n_3806),
.Y(n_4026)
);

O2A1O1Ixp33_ASAP7_75t_L g4027 ( 
.A1(n_3834),
.A2(n_202),
.B(n_207),
.C(n_208),
.Y(n_4027)
);

OAI22xp5_ASAP7_75t_L g4028 ( 
.A1(n_3831),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_4028)
);

AOI211xp5_ASAP7_75t_L g4029 ( 
.A1(n_3822),
.A2(n_209),
.B(n_214),
.C(n_215),
.Y(n_4029)
);

OA21x2_ASAP7_75t_L g4030 ( 
.A1(n_3866),
.A2(n_214),
.B(n_215),
.Y(n_4030)
);

O2A1O1Ixp33_ASAP7_75t_L g4031 ( 
.A1(n_3842),
.A2(n_216),
.B(n_220),
.C(n_224),
.Y(n_4031)
);

OAI22xp5_ASAP7_75t_L g4032 ( 
.A1(n_3861),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_3881),
.B(n_225),
.Y(n_4033)
);

OAI22xp5_ASAP7_75t_L g4034 ( 
.A1(n_3832),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_4034)
);

AOI21xp5_ASAP7_75t_SL g4035 ( 
.A1(n_3903),
.A2(n_227),
.B(n_229),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3906),
.B(n_232),
.Y(n_4036)
);

AND2x2_ASAP7_75t_L g4037 ( 
.A(n_3904),
.B(n_234),
.Y(n_4037)
);

INVx2_ASAP7_75t_L g4038 ( 
.A(n_3888),
.Y(n_4038)
);

AND2x2_ASAP7_75t_L g4039 ( 
.A(n_3933),
.B(n_234),
.Y(n_4039)
);

AOI21xp5_ASAP7_75t_L g4040 ( 
.A1(n_3808),
.A2(n_3846),
.B(n_3798),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_3827),
.B(n_235),
.Y(n_4041)
);

OAI22xp5_ASAP7_75t_L g4042 ( 
.A1(n_3898),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_3836),
.B(n_239),
.Y(n_4043)
);

O2A1O1Ixp33_ASAP7_75t_L g4044 ( 
.A1(n_3803),
.A2(n_240),
.B(n_241),
.C(n_242),
.Y(n_4044)
);

O2A1O1Ixp5_ASAP7_75t_L g4045 ( 
.A1(n_3901),
.A2(n_241),
.B(n_243),
.C(n_244),
.Y(n_4045)
);

AOI21xp5_ASAP7_75t_SL g4046 ( 
.A1(n_3786),
.A2(n_243),
.B(n_244),
.Y(n_4046)
);

O2A1O1Ixp33_ASAP7_75t_L g4047 ( 
.A1(n_3927),
.A2(n_245),
.B(n_246),
.C(n_247),
.Y(n_4047)
);

AND2x2_ASAP7_75t_L g4048 ( 
.A(n_3874),
.B(n_246),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_L g4049 ( 
.A(n_3837),
.B(n_248),
.Y(n_4049)
);

AOI21xp5_ASAP7_75t_L g4050 ( 
.A1(n_3843),
.A2(n_1767),
.B(n_1757),
.Y(n_4050)
);

AND2x2_ASAP7_75t_L g4051 ( 
.A(n_3874),
.B(n_248),
.Y(n_4051)
);

AND2x2_ASAP7_75t_L g4052 ( 
.A(n_3840),
.B(n_249),
.Y(n_4052)
);

INVx8_ASAP7_75t_L g4053 ( 
.A(n_3787),
.Y(n_4053)
);

BUFx6f_ASAP7_75t_L g4054 ( 
.A(n_3824),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3838),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3867),
.Y(n_4056)
);

INVx2_ASAP7_75t_L g4057 ( 
.A(n_3921),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_L g4058 ( 
.A(n_3939),
.B(n_249),
.Y(n_4058)
);

OAI22xp5_ASAP7_75t_L g4059 ( 
.A1(n_3900),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3892),
.B(n_252),
.Y(n_4060)
);

AND2x2_ASAP7_75t_L g4061 ( 
.A(n_3934),
.B(n_254),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3817),
.Y(n_4062)
);

HB1xp67_ASAP7_75t_L g4063 ( 
.A(n_3873),
.Y(n_4063)
);

AOI221x1_ASAP7_75t_SL g4064 ( 
.A1(n_3943),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.C(n_259),
.Y(n_4064)
);

CKINVDCx5p33_ASAP7_75t_R g4065 ( 
.A(n_3776),
.Y(n_4065)
);

OAI22xp5_ASAP7_75t_L g4066 ( 
.A1(n_3876),
.A2(n_256),
.B1(n_257),
.B2(n_259),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_3820),
.Y(n_4067)
);

NOR2xp33_ASAP7_75t_L g4068 ( 
.A(n_3775),
.B(n_3814),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_3816),
.B(n_261),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3945),
.Y(n_4070)
);

NOR2xp33_ASAP7_75t_L g4071 ( 
.A(n_3775),
.B(n_261),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_3805),
.Y(n_4072)
);

CKINVDCx5p33_ASAP7_75t_R g4073 ( 
.A(n_3830),
.Y(n_4073)
);

INVx3_ASAP7_75t_L g4074 ( 
.A(n_3896),
.Y(n_4074)
);

OAI22xp5_ASAP7_75t_L g4075 ( 
.A1(n_3938),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3849),
.Y(n_4076)
);

INVx2_ASAP7_75t_L g4077 ( 
.A(n_3896),
.Y(n_4077)
);

A2O1A1Ixp33_ASAP7_75t_L g4078 ( 
.A1(n_3825),
.A2(n_264),
.B(n_266),
.C(n_267),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_L g4079 ( 
.A(n_4067),
.B(n_3925),
.Y(n_4079)
);

CKINVDCx5p33_ASAP7_75t_R g4080 ( 
.A(n_3997),
.Y(n_4080)
);

BUFx3_ASAP7_75t_L g4081 ( 
.A(n_4003),
.Y(n_4081)
);

BUFx10_ASAP7_75t_L g4082 ( 
.A(n_3994),
.Y(n_4082)
);

AND2x2_ASAP7_75t_SL g4083 ( 
.A(n_3999),
.B(n_3864),
.Y(n_4083)
);

INVx2_ASAP7_75t_L g4084 ( 
.A(n_3992),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_3964),
.Y(n_4085)
);

AOI22xp33_ASAP7_75t_L g4086 ( 
.A1(n_3980),
.A2(n_3937),
.B1(n_3914),
.B2(n_3822),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3957),
.Y(n_4087)
);

NAND2xp33_ASAP7_75t_R g4088 ( 
.A(n_4073),
.B(n_3940),
.Y(n_4088)
);

INVx2_ASAP7_75t_L g4089 ( 
.A(n_3968),
.Y(n_4089)
);

AND2x4_ASAP7_75t_L g4090 ( 
.A(n_3963),
.B(n_3841),
.Y(n_4090)
);

CKINVDCx5p33_ASAP7_75t_R g4091 ( 
.A(n_4026),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_L g4092 ( 
.A(n_3972),
.B(n_3885),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_3955),
.B(n_3979),
.Y(n_4093)
);

OR2x2_ASAP7_75t_L g4094 ( 
.A(n_4062),
.B(n_3895),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_3946),
.B(n_3911),
.Y(n_4095)
);

NAND2xp33_ASAP7_75t_SL g4096 ( 
.A(n_3999),
.B(n_3910),
.Y(n_4096)
);

NOR2x1_ASAP7_75t_L g4097 ( 
.A(n_4021),
.B(n_3778),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_4006),
.B(n_3774),
.Y(n_4098)
);

AND2x2_ASAP7_75t_L g4099 ( 
.A(n_3986),
.B(n_3931),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_3965),
.Y(n_4100)
);

CKINVDCx5p33_ASAP7_75t_R g4101 ( 
.A(n_3962),
.Y(n_4101)
);

A2O1A1Ixp33_ASAP7_75t_L g4102 ( 
.A1(n_4064),
.A2(n_3930),
.B(n_3928),
.C(n_3865),
.Y(n_4102)
);

INVx2_ASAP7_75t_L g4103 ( 
.A(n_3952),
.Y(n_4103)
);

AND2x2_ASAP7_75t_L g4104 ( 
.A(n_3988),
.B(n_4077),
.Y(n_4104)
);

AND2x2_ASAP7_75t_L g4105 ( 
.A(n_3974),
.B(n_3833),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_L g4106 ( 
.A(n_4070),
.B(n_3778),
.Y(n_4106)
);

CKINVDCx5p33_ASAP7_75t_R g4107 ( 
.A(n_4065),
.Y(n_4107)
);

AOI22xp33_ASAP7_75t_L g4108 ( 
.A1(n_3980),
.A2(n_3924),
.B1(n_3923),
.B2(n_3843),
.Y(n_4108)
);

AND2x2_ASAP7_75t_L g4109 ( 
.A(n_3974),
.B(n_3835),
.Y(n_4109)
);

OR2x2_ASAP7_75t_L g4110 ( 
.A(n_4057),
.B(n_3853),
.Y(n_4110)
);

AND2x2_ASAP7_75t_L g4111 ( 
.A(n_3971),
.B(n_3941),
.Y(n_4111)
);

O2A1O1Ixp33_ASAP7_75t_L g4112 ( 
.A1(n_4060),
.A2(n_3871),
.B(n_3879),
.C(n_3823),
.Y(n_4112)
);

INVx2_ASAP7_75t_L g4113 ( 
.A(n_3989),
.Y(n_4113)
);

INVx1_ASAP7_75t_SL g4114 ( 
.A(n_4021),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_4056),
.Y(n_4115)
);

NOR2xp33_ASAP7_75t_L g4116 ( 
.A(n_4068),
.B(n_3787),
.Y(n_4116)
);

AND2x4_ASAP7_75t_L g4117 ( 
.A(n_3963),
.B(n_3841),
.Y(n_4117)
);

INVx2_ASAP7_75t_L g4118 ( 
.A(n_3973),
.Y(n_4118)
);

AND2x2_ASAP7_75t_L g4119 ( 
.A(n_4019),
.B(n_3929),
.Y(n_4119)
);

HB1xp67_ASAP7_75t_L g4120 ( 
.A(n_3969),
.Y(n_4120)
);

INVx2_ASAP7_75t_L g4121 ( 
.A(n_4007),
.Y(n_4121)
);

OR2x6_ASAP7_75t_L g4122 ( 
.A(n_3953),
.B(n_3787),
.Y(n_4122)
);

OAI21xp5_ASAP7_75t_L g4123 ( 
.A1(n_4040),
.A2(n_3815),
.B(n_3821),
.Y(n_4123)
);

AND2x2_ASAP7_75t_L g4124 ( 
.A(n_4019),
.B(n_3929),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_4055),
.B(n_3778),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_SL g4126 ( 
.A(n_3999),
.B(n_3782),
.Y(n_4126)
);

AOI22xp33_ASAP7_75t_L g4127 ( 
.A1(n_3980),
.A2(n_3843),
.B1(n_3811),
.B2(n_3889),
.Y(n_4127)
);

INVx2_ASAP7_75t_SL g4128 ( 
.A(n_4054),
.Y(n_4128)
);

OAI22xp5_ASAP7_75t_L g4129 ( 
.A1(n_4029),
.A2(n_3811),
.B1(n_3919),
.B2(n_3782),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_4005),
.Y(n_4130)
);

BUFx12f_ASAP7_75t_L g4131 ( 
.A(n_4054),
.Y(n_4131)
);

CKINVDCx16_ASAP7_75t_R g4132 ( 
.A(n_4008),
.Y(n_4132)
);

OR2x6_ASAP7_75t_L g4133 ( 
.A(n_3966),
.B(n_3844),
.Y(n_4133)
);

OAI22xp5_ASAP7_75t_L g4134 ( 
.A1(n_4029),
.A2(n_3811),
.B1(n_3782),
.B2(n_3795),
.Y(n_4134)
);

OR2x2_ASAP7_75t_L g4135 ( 
.A(n_4023),
.B(n_3853),
.Y(n_4135)
);

INVx2_ASAP7_75t_L g4136 ( 
.A(n_3984),
.Y(n_4136)
);

AND2x2_ASAP7_75t_L g4137 ( 
.A(n_4074),
.B(n_3853),
.Y(n_4137)
);

INVx2_ASAP7_75t_L g4138 ( 
.A(n_4038),
.Y(n_4138)
);

AO31x2_ASAP7_75t_L g4139 ( 
.A1(n_3998),
.A2(n_3875),
.A3(n_3779),
.B(n_3897),
.Y(n_4139)
);

OR2x2_ASAP7_75t_L g4140 ( 
.A(n_4001),
.B(n_3897),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_3959),
.Y(n_4141)
);

NOR3xp33_ASAP7_75t_SL g4142 ( 
.A(n_3954),
.B(n_3779),
.C(n_3875),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_3959),
.Y(n_4143)
);

NOR2xp33_ASAP7_75t_R g4144 ( 
.A(n_4054),
.B(n_3795),
.Y(n_4144)
);

AND2x2_ASAP7_75t_L g4145 ( 
.A(n_4074),
.B(n_3897),
.Y(n_4145)
);

OAI22xp5_ASAP7_75t_L g4146 ( 
.A1(n_3976),
.A2(n_3978),
.B1(n_4078),
.B2(n_3987),
.Y(n_4146)
);

BUFx2_ASAP7_75t_L g4147 ( 
.A(n_3958),
.Y(n_4147)
);

CKINVDCx20_ASAP7_75t_R g4148 ( 
.A(n_4004),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_3948),
.Y(n_4149)
);

NOR2xp33_ASAP7_75t_R g4150 ( 
.A(n_3994),
.B(n_3795),
.Y(n_4150)
);

A2O1A1Ixp33_ASAP7_75t_L g4151 ( 
.A1(n_4064),
.A2(n_3810),
.B(n_3797),
.C(n_3799),
.Y(n_4151)
);

CKINVDCx5p33_ASAP7_75t_R g4152 ( 
.A(n_4053),
.Y(n_4152)
);

INVxp67_ASAP7_75t_L g4153 ( 
.A(n_4012),
.Y(n_4153)
);

HB1xp67_ASAP7_75t_L g4154 ( 
.A(n_4063),
.Y(n_4154)
);

BUFx4f_ASAP7_75t_L g4155 ( 
.A(n_4053),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_4025),
.B(n_3802),
.Y(n_4156)
);

NAND3xp33_ASAP7_75t_L g4157 ( 
.A(n_4044),
.B(n_3785),
.C(n_3793),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_3948),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3967),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_3967),
.Y(n_4160)
);

CKINVDCx5p33_ASAP7_75t_R g4161 ( 
.A(n_4053),
.Y(n_4161)
);

OAI22xp5_ASAP7_75t_L g4162 ( 
.A1(n_3976),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_4030),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_SL g4164 ( 
.A(n_3949),
.B(n_1419),
.Y(n_4164)
);

CKINVDCx5p33_ASAP7_75t_R g4165 ( 
.A(n_4071),
.Y(n_4165)
);

HB1xp67_ASAP7_75t_L g4166 ( 
.A(n_4030),
.Y(n_4166)
);

AO31x2_ASAP7_75t_L g4167 ( 
.A1(n_3981),
.A2(n_269),
.A3(n_270),
.B(n_271),
.Y(n_4167)
);

INVx2_ASAP7_75t_L g4168 ( 
.A(n_4072),
.Y(n_4168)
);

AOI22xp33_ASAP7_75t_L g4169 ( 
.A1(n_3980),
.A2(n_1936),
.B1(n_1923),
.B2(n_1902),
.Y(n_4169)
);

HB1xp67_ASAP7_75t_L g4170 ( 
.A(n_4017),
.Y(n_4170)
);

NAND3xp33_ASAP7_75t_L g4171 ( 
.A(n_4027),
.B(n_4031),
.C(n_4020),
.Y(n_4171)
);

AND2x4_ASAP7_75t_L g4172 ( 
.A(n_4013),
.B(n_269),
.Y(n_4172)
);

AND2x2_ASAP7_75t_L g4173 ( 
.A(n_4076),
.B(n_270),
.Y(n_4173)
);

AND2x2_ASAP7_75t_L g4174 ( 
.A(n_4016),
.B(n_272),
.Y(n_4174)
);

BUFx12f_ASAP7_75t_L g4175 ( 
.A(n_4039),
.Y(n_4175)
);

INVx3_ASAP7_75t_L g4176 ( 
.A(n_4018),
.Y(n_4176)
);

OR2x2_ASAP7_75t_L g4177 ( 
.A(n_4002),
.B(n_273),
.Y(n_4177)
);

CKINVDCx5p33_ASAP7_75t_R g4178 ( 
.A(n_4048),
.Y(n_4178)
);

AND2x2_ASAP7_75t_L g4179 ( 
.A(n_4022),
.B(n_274),
.Y(n_4179)
);

OAI22xp33_ASAP7_75t_L g4180 ( 
.A1(n_3977),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_4180)
);

NAND2xp33_ASAP7_75t_R g4181 ( 
.A(n_4051),
.B(n_4061),
.Y(n_4181)
);

AND2x2_ASAP7_75t_L g4182 ( 
.A(n_3961),
.B(n_275),
.Y(n_4182)
);

INVx4_ASAP7_75t_L g4183 ( 
.A(n_4052),
.Y(n_4183)
);

CKINVDCx5p33_ASAP7_75t_R g4184 ( 
.A(n_4046),
.Y(n_4184)
);

NAND2xp33_ASAP7_75t_R g4185 ( 
.A(n_4036),
.B(n_277),
.Y(n_4185)
);

AO31x2_ASAP7_75t_L g4186 ( 
.A1(n_3981),
.A2(n_277),
.A3(n_279),
.B(n_280),
.Y(n_4186)
);

AND2x4_ASAP7_75t_L g4187 ( 
.A(n_3961),
.B(n_279),
.Y(n_4187)
);

NOR2xp33_ASAP7_75t_R g4188 ( 
.A(n_4058),
.B(n_4069),
.Y(n_4188)
);

NOR2xp33_ASAP7_75t_R g4189 ( 
.A(n_4037),
.B(n_280),
.Y(n_4189)
);

AND2x4_ASAP7_75t_L g4190 ( 
.A(n_3991),
.B(n_329),
.Y(n_4190)
);

BUFx6f_ASAP7_75t_L g4191 ( 
.A(n_4041),
.Y(n_4191)
);

INVx2_ASAP7_75t_L g4192 ( 
.A(n_4033),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_3947),
.B(n_330),
.Y(n_4193)
);

INVx2_ASAP7_75t_L g4194 ( 
.A(n_4043),
.Y(n_4194)
);

BUFx3_ASAP7_75t_L g4195 ( 
.A(n_4049),
.Y(n_4195)
);

INVxp67_ASAP7_75t_SL g4196 ( 
.A(n_4000),
.Y(n_4196)
);

OR2x2_ASAP7_75t_L g4197 ( 
.A(n_3982),
.B(n_331),
.Y(n_4197)
);

BUFx3_ASAP7_75t_L g4198 ( 
.A(n_4009),
.Y(n_4198)
);

BUFx6f_ASAP7_75t_L g4199 ( 
.A(n_4009),
.Y(n_4199)
);

AO31x2_ASAP7_75t_L g4200 ( 
.A1(n_3982),
.A2(n_335),
.A3(n_342),
.B(n_343),
.Y(n_4200)
);

AND2x2_ASAP7_75t_L g4201 ( 
.A(n_3993),
.B(n_3970),
.Y(n_4201)
);

OR2x2_ASAP7_75t_L g4202 ( 
.A(n_3975),
.B(n_344),
.Y(n_4202)
);

AND2x2_ASAP7_75t_L g4203 ( 
.A(n_3996),
.B(n_345),
.Y(n_4203)
);

INVx2_ASAP7_75t_L g4204 ( 
.A(n_4149),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4087),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_4100),
.Y(n_4206)
);

INVx2_ASAP7_75t_L g4207 ( 
.A(n_4158),
.Y(n_4207)
);

AND2x2_ASAP7_75t_L g4208 ( 
.A(n_4201),
.B(n_3996),
.Y(n_4208)
);

INVx2_ASAP7_75t_L g4209 ( 
.A(n_4141),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_4115),
.Y(n_4210)
);

INVx2_ASAP7_75t_L g4211 ( 
.A(n_4143),
.Y(n_4211)
);

OR2x2_ASAP7_75t_L g4212 ( 
.A(n_4114),
.B(n_3975),
.Y(n_4212)
);

AND2x2_ASAP7_75t_L g4213 ( 
.A(n_4133),
.B(n_3995),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_4118),
.Y(n_4214)
);

INVx2_ASAP7_75t_L g4215 ( 
.A(n_4159),
.Y(n_4215)
);

INVx2_ASAP7_75t_L g4216 ( 
.A(n_4160),
.Y(n_4216)
);

AO21x2_ASAP7_75t_L g4217 ( 
.A1(n_4166),
.A2(n_3983),
.B(n_3985),
.Y(n_4217)
);

OAI321xp33_ASAP7_75t_L g4218 ( 
.A1(n_4146),
.A2(n_4162),
.A3(n_4134),
.B1(n_4171),
.B2(n_4129),
.C(n_4157),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_4121),
.Y(n_4219)
);

AND2x2_ASAP7_75t_L g4220 ( 
.A(n_4133),
.B(n_3995),
.Y(n_4220)
);

OR2x6_ASAP7_75t_L g4221 ( 
.A(n_4133),
.B(n_4024),
.Y(n_4221)
);

AND2x2_ASAP7_75t_L g4222 ( 
.A(n_4198),
.B(n_4015),
.Y(n_4222)
);

OAI21x1_ASAP7_75t_L g4223 ( 
.A1(n_4097),
.A2(n_3990),
.B(n_4050),
.Y(n_4223)
);

AND2x2_ASAP7_75t_L g4224 ( 
.A(n_4147),
.B(n_3990),
.Y(n_4224)
);

OAI22xp5_ASAP7_75t_L g4225 ( 
.A1(n_4146),
.A2(n_3956),
.B1(n_3960),
.B2(n_3951),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_4085),
.B(n_4035),
.Y(n_4226)
);

AND2x2_ASAP7_75t_L g4227 ( 
.A(n_4089),
.B(n_3950),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_4163),
.Y(n_4228)
);

AND2x2_ASAP7_75t_L g4229 ( 
.A(n_4084),
.B(n_4011),
.Y(n_4229)
);

AND2x2_ASAP7_75t_L g4230 ( 
.A(n_4154),
.B(n_4045),
.Y(n_4230)
);

INVx2_ASAP7_75t_L g4231 ( 
.A(n_4199),
.Y(n_4231)
);

INVx4_ASAP7_75t_L g4232 ( 
.A(n_4131),
.Y(n_4232)
);

AOI22xp33_ASAP7_75t_L g4233 ( 
.A1(n_4171),
.A2(n_4075),
.B1(n_4032),
.B2(n_4042),
.Y(n_4233)
);

INVx2_ASAP7_75t_L g4234 ( 
.A(n_4199),
.Y(n_4234)
);

AO21x2_ASAP7_75t_L g4235 ( 
.A1(n_4162),
.A2(n_4028),
.B(n_4034),
.Y(n_4235)
);

OA21x2_ASAP7_75t_L g4236 ( 
.A1(n_4114),
.A2(n_4010),
.B(n_4059),
.Y(n_4236)
);

AND2x2_ASAP7_75t_L g4237 ( 
.A(n_4137),
.B(n_4066),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_4130),
.Y(n_4238)
);

INVx4_ASAP7_75t_L g4239 ( 
.A(n_4082),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4120),
.Y(n_4240)
);

AND2x2_ASAP7_75t_L g4241 ( 
.A(n_4145),
.B(n_4047),
.Y(n_4241)
);

AND2x2_ASAP7_75t_L g4242 ( 
.A(n_4139),
.B(n_4014),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_4136),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_4138),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4170),
.Y(n_4245)
);

AOI21xp5_ASAP7_75t_L g4246 ( 
.A1(n_4134),
.A2(n_346),
.B(n_348),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4167),
.Y(n_4247)
);

INVx2_ASAP7_75t_L g4248 ( 
.A(n_4199),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_4167),
.Y(n_4249)
);

INVx6_ASAP7_75t_L g4250 ( 
.A(n_4082),
.Y(n_4250)
);

OAI211xp5_ASAP7_75t_SL g4251 ( 
.A1(n_4086),
.A2(n_350),
.B(n_353),
.C(n_356),
.Y(n_4251)
);

OR2x2_ASAP7_75t_L g4252 ( 
.A(n_4196),
.B(n_360),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4167),
.Y(n_4253)
);

AO21x2_ASAP7_75t_L g4254 ( 
.A1(n_4202),
.A2(n_362),
.B(n_368),
.Y(n_4254)
);

INVxp67_ASAP7_75t_R g4255 ( 
.A(n_4129),
.Y(n_4255)
);

BUFx3_ASAP7_75t_L g4256 ( 
.A(n_4080),
.Y(n_4256)
);

INVx2_ASAP7_75t_L g4257 ( 
.A(n_4097),
.Y(n_4257)
);

OR2x2_ASAP7_75t_L g4258 ( 
.A(n_4093),
.B(n_370),
.Y(n_4258)
);

INVx2_ASAP7_75t_L g4259 ( 
.A(n_4176),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_4186),
.Y(n_4260)
);

INVx3_ASAP7_75t_L g4261 ( 
.A(n_4139),
.Y(n_4261)
);

INVxp67_ASAP7_75t_L g4262 ( 
.A(n_4185),
.Y(n_4262)
);

AO21x2_ASAP7_75t_L g4263 ( 
.A1(n_4203),
.A2(n_372),
.B(n_373),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4186),
.Y(n_4264)
);

HB1xp67_ASAP7_75t_L g4265 ( 
.A(n_4186),
.Y(n_4265)
);

INVx2_ASAP7_75t_L g4266 ( 
.A(n_4176),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_4153),
.Y(n_4267)
);

OA21x2_ASAP7_75t_L g4268 ( 
.A1(n_4157),
.A2(n_376),
.B(n_381),
.Y(n_4268)
);

INVx2_ASAP7_75t_SL g4269 ( 
.A(n_4090),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_4168),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_4113),
.Y(n_4271)
);

HB1xp67_ASAP7_75t_L g4272 ( 
.A(n_4191),
.Y(n_4272)
);

AND2x2_ASAP7_75t_L g4273 ( 
.A(n_4139),
.B(n_391),
.Y(n_4273)
);

OA21x2_ASAP7_75t_L g4274 ( 
.A1(n_4098),
.A2(n_392),
.B(n_393),
.Y(n_4274)
);

AOI21x1_ASAP7_75t_L g4275 ( 
.A1(n_4126),
.A2(n_394),
.B(n_409),
.Y(n_4275)
);

AND2x2_ASAP7_75t_L g4276 ( 
.A(n_4103),
.B(n_410),
.Y(n_4276)
);

AOI22xp33_ASAP7_75t_L g4277 ( 
.A1(n_4123),
.A2(n_1425),
.B1(n_1433),
.B2(n_1440),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_4192),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_SL g4279 ( 
.A(n_4142),
.B(n_1425),
.Y(n_4279)
);

AO21x2_ASAP7_75t_L g4280 ( 
.A1(n_4182),
.A2(n_411),
.B(n_415),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_4194),
.B(n_419),
.Y(n_4281)
);

INVx5_ASAP7_75t_L g4282 ( 
.A(n_4122),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_4135),
.Y(n_4283)
);

INVx2_ASAP7_75t_L g4284 ( 
.A(n_4110),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_4187),
.Y(n_4285)
);

INVx2_ASAP7_75t_L g4286 ( 
.A(n_4187),
.Y(n_4286)
);

OR2x2_ASAP7_75t_L g4287 ( 
.A(n_4079),
.B(n_428),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_4094),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_4125),
.Y(n_4289)
);

AO21x2_ASAP7_75t_L g4290 ( 
.A1(n_4193),
.A2(n_429),
.B(n_430),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4140),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_4191),
.Y(n_4292)
);

INVx3_ASAP7_75t_L g4293 ( 
.A(n_4122),
.Y(n_4293)
);

NAND3xp33_ASAP7_75t_L g4294 ( 
.A(n_4151),
.B(n_1425),
.C(n_1433),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_4104),
.Y(n_4295)
);

BUFx2_ASAP7_75t_L g4296 ( 
.A(n_4122),
.Y(n_4296)
);

AO21x2_ASAP7_75t_L g4297 ( 
.A1(n_4180),
.A2(n_434),
.B(n_436),
.Y(n_4297)
);

HB1xp67_ASAP7_75t_L g4298 ( 
.A(n_4191),
.Y(n_4298)
);

INVxp67_ASAP7_75t_SL g4299 ( 
.A(n_4181),
.Y(n_4299)
);

AO21x2_ASAP7_75t_L g4300 ( 
.A1(n_4123),
.A2(n_437),
.B(n_443),
.Y(n_4300)
);

INVx2_ASAP7_75t_L g4301 ( 
.A(n_4190),
.Y(n_4301)
);

INVxp67_ASAP7_75t_L g4302 ( 
.A(n_4156),
.Y(n_4302)
);

AO21x2_ASAP7_75t_L g4303 ( 
.A1(n_4197),
.A2(n_446),
.B(n_450),
.Y(n_4303)
);

INVx2_ASAP7_75t_SL g4304 ( 
.A(n_4250),
.Y(n_4304)
);

AND2x2_ASAP7_75t_L g4305 ( 
.A(n_4299),
.B(n_4090),
.Y(n_4305)
);

HB1xp67_ASAP7_75t_L g4306 ( 
.A(n_4272),
.Y(n_4306)
);

INVx2_ASAP7_75t_L g4307 ( 
.A(n_4231),
.Y(n_4307)
);

AND2x2_ASAP7_75t_L g4308 ( 
.A(n_4282),
.B(n_4117),
.Y(n_4308)
);

INVx2_ASAP7_75t_L g4309 ( 
.A(n_4231),
.Y(n_4309)
);

OR2x2_ASAP7_75t_L g4310 ( 
.A(n_4245),
.B(n_4247),
.Y(n_4310)
);

AND2x4_ASAP7_75t_SL g4311 ( 
.A(n_4221),
.B(n_4117),
.Y(n_4311)
);

CKINVDCx14_ASAP7_75t_R g4312 ( 
.A(n_4232),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_L g4313 ( 
.A(n_4241),
.B(n_4195),
.Y(n_4313)
);

OR2x2_ASAP7_75t_L g4314 ( 
.A(n_4245),
.B(n_4095),
.Y(n_4314)
);

INVx2_ASAP7_75t_L g4315 ( 
.A(n_4234),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4228),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4228),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_4241),
.B(n_4188),
.Y(n_4318)
);

AND2x2_ASAP7_75t_L g4319 ( 
.A(n_4282),
.B(n_4109),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4205),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_4205),
.Y(n_4321)
);

INVx2_ASAP7_75t_L g4322 ( 
.A(n_4234),
.Y(n_4322)
);

AND2x2_ASAP7_75t_L g4323 ( 
.A(n_4282),
.B(n_4119),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4206),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_4206),
.Y(n_4325)
);

INVx2_ASAP7_75t_L g4326 ( 
.A(n_4248),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4210),
.Y(n_4327)
);

INVxp67_ASAP7_75t_L g4328 ( 
.A(n_4262),
.Y(n_4328)
);

AND2x2_ASAP7_75t_L g4329 ( 
.A(n_4282),
.B(n_4124),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4210),
.Y(n_4330)
);

AOI22xp33_ASAP7_75t_L g4331 ( 
.A1(n_4225),
.A2(n_4184),
.B1(n_4096),
.B2(n_4127),
.Y(n_4331)
);

AND2x2_ASAP7_75t_L g4332 ( 
.A(n_4282),
.B(n_4105),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4278),
.Y(n_4333)
);

AND2x4_ASAP7_75t_L g4334 ( 
.A(n_4282),
.B(n_4190),
.Y(n_4334)
);

AND2x2_ASAP7_75t_L g4335 ( 
.A(n_4269),
.B(n_4083),
.Y(n_4335)
);

INVx2_ASAP7_75t_L g4336 ( 
.A(n_4248),
.Y(n_4336)
);

HB1xp67_ASAP7_75t_L g4337 ( 
.A(n_4298),
.Y(n_4337)
);

AND2x2_ASAP7_75t_L g4338 ( 
.A(n_4269),
.B(n_4099),
.Y(n_4338)
);

NOR2xp33_ASAP7_75t_L g4339 ( 
.A(n_4232),
.B(n_4239),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_4302),
.B(n_4173),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_4278),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_4267),
.Y(n_4342)
);

OAI22xp5_ASAP7_75t_L g4343 ( 
.A1(n_4221),
.A2(n_4108),
.B1(n_4169),
.B2(n_4102),
.Y(n_4343)
);

AND2x2_ASAP7_75t_L g4344 ( 
.A(n_4296),
.B(n_4150),
.Y(n_4344)
);

AND2x2_ASAP7_75t_L g4345 ( 
.A(n_4296),
.B(n_4183),
.Y(n_4345)
);

AND2x2_ASAP7_75t_L g4346 ( 
.A(n_4222),
.B(n_4183),
.Y(n_4346)
);

INVx4_ASAP7_75t_L g4347 ( 
.A(n_4232),
.Y(n_4347)
);

INVx1_ASAP7_75t_L g4348 ( 
.A(n_4267),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_L g4349 ( 
.A(n_4227),
.B(n_4177),
.Y(n_4349)
);

OR2x2_ASAP7_75t_L g4350 ( 
.A(n_4247),
.B(n_4249),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4214),
.Y(n_4351)
);

OR2x2_ASAP7_75t_L g4352 ( 
.A(n_4249),
.B(n_4092),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4214),
.Y(n_4353)
);

BUFx2_ASAP7_75t_L g4354 ( 
.A(n_4239),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_4219),
.Y(n_4355)
);

HB1xp67_ASAP7_75t_L g4356 ( 
.A(n_4259),
.Y(n_4356)
);

NAND2xp5_ASAP7_75t_L g4357 ( 
.A(n_4227),
.B(n_4174),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4219),
.Y(n_4358)
);

AND2x2_ASAP7_75t_L g4359 ( 
.A(n_4222),
.B(n_4293),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4215),
.Y(n_4360)
);

AND2x2_ASAP7_75t_L g4361 ( 
.A(n_4293),
.B(n_4132),
.Y(n_4361)
);

AND2x2_ASAP7_75t_L g4362 ( 
.A(n_4293),
.B(n_4128),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4288),
.Y(n_4363)
);

INVx2_ASAP7_75t_L g4364 ( 
.A(n_4204),
.Y(n_4364)
);

INVxp67_ASAP7_75t_L g4365 ( 
.A(n_4265),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_4292),
.B(n_4172),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4215),
.Y(n_4367)
);

BUFx2_ASAP7_75t_L g4368 ( 
.A(n_4239),
.Y(n_4368)
);

INVxp67_ASAP7_75t_SL g4369 ( 
.A(n_4257),
.Y(n_4369)
);

OAI22xp33_ASAP7_75t_L g4370 ( 
.A1(n_4343),
.A2(n_4255),
.B1(n_4221),
.B2(n_4218),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4350),
.Y(n_4371)
);

AOI22xp33_ASAP7_75t_L g4372 ( 
.A1(n_4361),
.A2(n_4217),
.B1(n_4268),
.B2(n_4235),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_4328),
.B(n_4365),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_4350),
.Y(n_4374)
);

INVxp67_ASAP7_75t_L g4375 ( 
.A(n_4354),
.Y(n_4375)
);

AND2x2_ASAP7_75t_L g4376 ( 
.A(n_4361),
.B(n_4255),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_4310),
.Y(n_4377)
);

HB1xp67_ASAP7_75t_L g4378 ( 
.A(n_4306),
.Y(n_4378)
);

INVx2_ASAP7_75t_L g4379 ( 
.A(n_4305),
.Y(n_4379)
);

AND2x4_ASAP7_75t_L g4380 ( 
.A(n_4305),
.B(n_4292),
.Y(n_4380)
);

INVx2_ASAP7_75t_L g4381 ( 
.A(n_4338),
.Y(n_4381)
);

INVx4_ASAP7_75t_SL g4382 ( 
.A(n_4354),
.Y(n_4382)
);

OR2x6_ASAP7_75t_L g4383 ( 
.A(n_4368),
.B(n_4250),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_4338),
.Y(n_4384)
);

OAI33xp33_ASAP7_75t_L g4385 ( 
.A1(n_4342),
.A2(n_4264),
.A3(n_4253),
.B1(n_4260),
.B2(n_4294),
.B3(n_4212),
.Y(n_4385)
);

AOI221xp5_ASAP7_75t_L g4386 ( 
.A1(n_4348),
.A2(n_4217),
.B1(n_4253),
.B2(n_4264),
.C(n_4260),
.Y(n_4386)
);

AND2x4_ASAP7_75t_SL g4387 ( 
.A(n_4319),
.B(n_4221),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_L g4388 ( 
.A(n_4337),
.B(n_4229),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_4310),
.Y(n_4389)
);

OAI221xp5_ASAP7_75t_L g4390 ( 
.A1(n_4331),
.A2(n_4233),
.B1(n_4236),
.B2(n_4268),
.C(n_4208),
.Y(n_4390)
);

OR2x2_ASAP7_75t_L g4391 ( 
.A(n_4349),
.B(n_4288),
.Y(n_4391)
);

OAI31xp33_ASAP7_75t_L g4392 ( 
.A1(n_4311),
.A2(n_4230),
.A3(n_4242),
.B(n_4208),
.Y(n_4392)
);

HB1xp67_ASAP7_75t_L g4393 ( 
.A(n_4356),
.Y(n_4393)
);

NAND4xp25_ASAP7_75t_SL g4394 ( 
.A(n_4318),
.B(n_4242),
.C(n_4246),
.D(n_4230),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4321),
.Y(n_4395)
);

AOI22xp33_ASAP7_75t_SL g4396 ( 
.A1(n_4335),
.A2(n_4217),
.B1(n_4236),
.B2(n_4235),
.Y(n_4396)
);

INVx1_ASAP7_75t_SL g4397 ( 
.A(n_4344),
.Y(n_4397)
);

OA222x2_ASAP7_75t_L g4398 ( 
.A1(n_4313),
.A2(n_4212),
.B1(n_4257),
.B2(n_4261),
.C1(n_4266),
.C2(n_4259),
.Y(n_4398)
);

NOR2xp33_ASAP7_75t_R g4399 ( 
.A(n_4312),
.B(n_4256),
.Y(n_4399)
);

BUFx3_ASAP7_75t_L g4400 ( 
.A(n_4319),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_4321),
.Y(n_4401)
);

NOR2xp33_ASAP7_75t_L g4402 ( 
.A(n_4347),
.B(n_4250),
.Y(n_4402)
);

OAI211xp5_ASAP7_75t_SL g4403 ( 
.A1(n_4339),
.A2(n_4287),
.B(n_4301),
.C(n_4286),
.Y(n_4403)
);

AOI22xp33_ASAP7_75t_L g4404 ( 
.A1(n_4332),
.A2(n_4268),
.B1(n_4235),
.B2(n_4236),
.Y(n_4404)
);

INVxp67_ASAP7_75t_L g4405 ( 
.A(n_4368),
.Y(n_4405)
);

AND2x2_ASAP7_75t_L g4406 ( 
.A(n_4344),
.B(n_4250),
.Y(n_4406)
);

INVx1_ASAP7_75t_SL g4407 ( 
.A(n_4345),
.Y(n_4407)
);

NOR2x2_ASAP7_75t_L g4408 ( 
.A(n_4307),
.B(n_4285),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4324),
.Y(n_4409)
);

OAI211xp5_ASAP7_75t_L g4410 ( 
.A1(n_4345),
.A2(n_4268),
.B(n_4236),
.C(n_4189),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_4393),
.Y(n_4411)
);

NAND2x1p5_ASAP7_75t_L g4412 ( 
.A(n_4397),
.B(n_4347),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4378),
.Y(n_4413)
);

INVxp67_ASAP7_75t_SL g4414 ( 
.A(n_4388),
.Y(n_4414)
);

AND2x2_ASAP7_75t_L g4415 ( 
.A(n_4376),
.B(n_4308),
.Y(n_4415)
);

NOR2xp33_ASAP7_75t_L g4416 ( 
.A(n_4402),
.B(n_4347),
.Y(n_4416)
);

BUFx2_ASAP7_75t_L g4417 ( 
.A(n_4399),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4377),
.Y(n_4418)
);

OR2x2_ASAP7_75t_L g4419 ( 
.A(n_4388),
.B(n_4397),
.Y(n_4419)
);

AND2x2_ASAP7_75t_L g4420 ( 
.A(n_4406),
.B(n_4308),
.Y(n_4420)
);

AND2x2_ASAP7_75t_L g4421 ( 
.A(n_4400),
.B(n_4335),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_4389),
.Y(n_4422)
);

AND2x4_ASAP7_75t_L g4423 ( 
.A(n_4382),
.B(n_4311),
.Y(n_4423)
);

INVx2_ASAP7_75t_L g4424 ( 
.A(n_4382),
.Y(n_4424)
);

OR2x2_ASAP7_75t_L g4425 ( 
.A(n_4379),
.B(n_4314),
.Y(n_4425)
);

INVx1_ASAP7_75t_SL g4426 ( 
.A(n_4408),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_4382),
.Y(n_4427)
);

INVx2_ASAP7_75t_L g4428 ( 
.A(n_4383),
.Y(n_4428)
);

OR2x2_ASAP7_75t_L g4429 ( 
.A(n_4407),
.B(n_4314),
.Y(n_4429)
);

INVx2_ASAP7_75t_L g4430 ( 
.A(n_4383),
.Y(n_4430)
);

AND2x2_ASAP7_75t_L g4431 ( 
.A(n_4407),
.B(n_4362),
.Y(n_4431)
);

AND2x2_ASAP7_75t_L g4432 ( 
.A(n_4380),
.B(n_4362),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_4371),
.Y(n_4433)
);

INVx2_ASAP7_75t_L g4434 ( 
.A(n_4383),
.Y(n_4434)
);

AND2x2_ASAP7_75t_L g4435 ( 
.A(n_4380),
.B(n_4332),
.Y(n_4435)
);

INVx2_ASAP7_75t_L g4436 ( 
.A(n_4381),
.Y(n_4436)
);

AND2x2_ASAP7_75t_L g4437 ( 
.A(n_4384),
.B(n_4323),
.Y(n_4437)
);

NOR2xp33_ASAP7_75t_L g4438 ( 
.A(n_4417),
.B(n_4413),
.Y(n_4438)
);

AND2x2_ASAP7_75t_L g4439 ( 
.A(n_4417),
.B(n_4346),
.Y(n_4439)
);

HB1xp67_ASAP7_75t_L g4440 ( 
.A(n_4431),
.Y(n_4440)
);

AND2x2_ASAP7_75t_L g4441 ( 
.A(n_4415),
.B(n_4346),
.Y(n_4441)
);

OR2x2_ASAP7_75t_L g4442 ( 
.A(n_4426),
.B(n_4373),
.Y(n_4442)
);

INVx1_ASAP7_75t_L g4443 ( 
.A(n_4429),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_L g4444 ( 
.A(n_4431),
.B(n_4375),
.Y(n_4444)
);

OR2x2_ASAP7_75t_L g4445 ( 
.A(n_4419),
.B(n_4373),
.Y(n_4445)
);

AND2x2_ASAP7_75t_L g4446 ( 
.A(n_4415),
.B(n_4359),
.Y(n_4446)
);

INVx2_ASAP7_75t_L g4447 ( 
.A(n_4412),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_4429),
.Y(n_4448)
);

INVx1_ASAP7_75t_L g4449 ( 
.A(n_4413),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_L g4450 ( 
.A(n_4432),
.B(n_4405),
.Y(n_4450)
);

AND2x2_ASAP7_75t_L g4451 ( 
.A(n_4420),
.B(n_4387),
.Y(n_4451)
);

INVx2_ASAP7_75t_L g4452 ( 
.A(n_4412),
.Y(n_4452)
);

NAND3xp33_ASAP7_75t_L g4453 ( 
.A(n_4428),
.B(n_4396),
.C(n_4372),
.Y(n_4453)
);

AND2x2_ASAP7_75t_L g4454 ( 
.A(n_4420),
.B(n_4304),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_4412),
.Y(n_4455)
);

NAND2xp5_ASAP7_75t_L g4456 ( 
.A(n_4446),
.B(n_4428),
.Y(n_4456)
);

OR2x2_ASAP7_75t_L g4457 ( 
.A(n_4442),
.B(n_4419),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_4446),
.B(n_4430),
.Y(n_4458)
);

OR2x2_ASAP7_75t_L g4459 ( 
.A(n_4440),
.B(n_4444),
.Y(n_4459)
);

AOI22xp5_ASAP7_75t_L g4460 ( 
.A1(n_4439),
.A2(n_4370),
.B1(n_4394),
.B2(n_4410),
.Y(n_4460)
);

BUFx2_ASAP7_75t_L g4461 ( 
.A(n_4440),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_L g4462 ( 
.A(n_4438),
.B(n_4443),
.Y(n_4462)
);

OAI22xp33_ASAP7_75t_SL g4463 ( 
.A1(n_4445),
.A2(n_4390),
.B1(n_4414),
.B2(n_4398),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_L g4464 ( 
.A(n_4438),
.B(n_4441),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_4448),
.Y(n_4465)
);

AND2x2_ASAP7_75t_L g4466 ( 
.A(n_4441),
.B(n_4432),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_4454),
.B(n_4430),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_4450),
.Y(n_4468)
);

AND2x2_ASAP7_75t_L g4469 ( 
.A(n_4451),
.B(n_4421),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4449),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_4447),
.Y(n_4471)
);

AND2x2_ASAP7_75t_L g4472 ( 
.A(n_4447),
.B(n_4421),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_4452),
.Y(n_4473)
);

OAI22xp5_ASAP7_75t_L g4474 ( 
.A1(n_4460),
.A2(n_4404),
.B1(n_4453),
.B2(n_4304),
.Y(n_4474)
);

OR2x2_ASAP7_75t_L g4475 ( 
.A(n_4464),
.B(n_4425),
.Y(n_4475)
);

OAI22xp5_ASAP7_75t_L g4476 ( 
.A1(n_4457),
.A2(n_4357),
.B1(n_4423),
.B2(n_4434),
.Y(n_4476)
);

NOR2x1_ASAP7_75t_L g4477 ( 
.A(n_4461),
.B(n_4427),
.Y(n_4477)
);

HB1xp67_ASAP7_75t_L g4478 ( 
.A(n_4466),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_4472),
.B(n_4434),
.Y(n_4479)
);

BUFx2_ASAP7_75t_L g4480 ( 
.A(n_4469),
.Y(n_4480)
);

NAND2xp5_ASAP7_75t_L g4481 ( 
.A(n_4465),
.B(n_4411),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_4456),
.Y(n_4482)
);

NOR2xp67_ASAP7_75t_SL g4483 ( 
.A(n_4459),
.B(n_4427),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_L g4484 ( 
.A(n_4467),
.B(n_4411),
.Y(n_4484)
);

INVx2_ASAP7_75t_SL g4485 ( 
.A(n_4458),
.Y(n_4485)
);

INVx1_ASAP7_75t_L g4486 ( 
.A(n_4478),
.Y(n_4486)
);

AND2x2_ASAP7_75t_L g4487 ( 
.A(n_4480),
.B(n_4435),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_4477),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4479),
.Y(n_4489)
);

INVx2_ASAP7_75t_L g4490 ( 
.A(n_4485),
.Y(n_4490)
);

AND2x2_ASAP7_75t_L g4491 ( 
.A(n_4482),
.B(n_4435),
.Y(n_4491)
);

NOR2xp33_ASAP7_75t_L g4492 ( 
.A(n_4476),
.B(n_4462),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_L g4493 ( 
.A(n_4483),
.B(n_4424),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_L g4494 ( 
.A(n_4484),
.B(n_4463),
.Y(n_4494)
);

OAI221xp5_ASAP7_75t_L g4495 ( 
.A1(n_4494),
.A2(n_4463),
.B1(n_4474),
.B2(n_4462),
.C(n_4416),
.Y(n_4495)
);

INVx1_ASAP7_75t_SL g4496 ( 
.A(n_4487),
.Y(n_4496)
);

NAND2xp5_ASAP7_75t_L g4497 ( 
.A(n_4486),
.B(n_4424),
.Y(n_4497)
);

OAI22xp33_ASAP7_75t_L g4498 ( 
.A1(n_4494),
.A2(n_4475),
.B1(n_4425),
.B2(n_4386),
.Y(n_4498)
);

BUFx2_ASAP7_75t_L g4499 ( 
.A(n_4488),
.Y(n_4499)
);

BUFx2_ASAP7_75t_L g4500 ( 
.A(n_4493),
.Y(n_4500)
);

AOI221xp5_ASAP7_75t_L g4501 ( 
.A1(n_4492),
.A2(n_4385),
.B1(n_4481),
.B2(n_4468),
.C(n_4394),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_L g4502 ( 
.A(n_4491),
.B(n_4471),
.Y(n_4502)
);

AND2x2_ASAP7_75t_L g4503 ( 
.A(n_4490),
.B(n_4437),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4489),
.Y(n_4504)
);

OAI22xp33_ASAP7_75t_SL g4505 ( 
.A1(n_4494),
.A2(n_4423),
.B1(n_4455),
.B2(n_4452),
.Y(n_4505)
);

AND2x2_ASAP7_75t_L g4506 ( 
.A(n_4487),
.B(n_4437),
.Y(n_4506)
);

OR2x2_ASAP7_75t_L g4507 ( 
.A(n_4496),
.B(n_4436),
.Y(n_4507)
);

HB1xp67_ASAP7_75t_L g4508 ( 
.A(n_4506),
.Y(n_4508)
);

INVxp33_ASAP7_75t_L g4509 ( 
.A(n_4503),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4502),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_4497),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_L g4512 ( 
.A(n_4505),
.B(n_4473),
.Y(n_4512)
);

OAI21xp33_ASAP7_75t_L g4513 ( 
.A1(n_4495),
.A2(n_4423),
.B(n_4501),
.Y(n_4513)
);

AOI22xp5_ASAP7_75t_L g4514 ( 
.A1(n_4498),
.A2(n_4423),
.B1(n_4436),
.B2(n_4403),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4500),
.Y(n_4515)
);

NAND2xp5_ASAP7_75t_L g4516 ( 
.A(n_4508),
.B(n_4499),
.Y(n_4516)
);

AOI22xp33_ASAP7_75t_L g4517 ( 
.A1(n_4513),
.A2(n_4455),
.B1(n_4392),
.B2(n_4418),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_4512),
.Y(n_4518)
);

INVxp67_ASAP7_75t_L g4519 ( 
.A(n_4507),
.Y(n_4519)
);

NOR2xp33_ASAP7_75t_L g4520 ( 
.A(n_4509),
.B(n_4504),
.Y(n_4520)
);

OR2x2_ASAP7_75t_L g4521 ( 
.A(n_4514),
.B(n_4418),
.Y(n_4521)
);

NOR2xp33_ASAP7_75t_L g4522 ( 
.A(n_4515),
.B(n_4470),
.Y(n_4522)
);

INVx1_ASAP7_75t_L g4523 ( 
.A(n_4511),
.Y(n_4523)
);

NOR2xp33_ASAP7_75t_L g4524 ( 
.A(n_4510),
.B(n_4256),
.Y(n_4524)
);

NAND2xp5_ASAP7_75t_L g4525 ( 
.A(n_4517),
.B(n_4422),
.Y(n_4525)
);

NOR3x1_ASAP7_75t_L g4526 ( 
.A(n_4516),
.B(n_4518),
.C(n_4521),
.Y(n_4526)
);

NOR2xp33_ASAP7_75t_L g4527 ( 
.A(n_4519),
.B(n_4422),
.Y(n_4527)
);

INVx1_ASAP7_75t_L g4528 ( 
.A(n_4520),
.Y(n_4528)
);

NAND3xp33_ASAP7_75t_L g4529 ( 
.A(n_4524),
.B(n_4433),
.C(n_4374),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_SL g4530 ( 
.A(n_4522),
.B(n_4433),
.Y(n_4530)
);

AND4x1_ASAP7_75t_L g4531 ( 
.A(n_4523),
.B(n_4359),
.C(n_4116),
.D(n_4273),
.Y(n_4531)
);

NOR2x1_ASAP7_75t_L g4532 ( 
.A(n_4516),
.B(n_4395),
.Y(n_4532)
);

HB1xp67_ASAP7_75t_L g4533 ( 
.A(n_4516),
.Y(n_4533)
);

AOI211x1_ASAP7_75t_L g4534 ( 
.A1(n_4516),
.A2(n_4401),
.B(n_4409),
.C(n_4317),
.Y(n_4534)
);

HB1xp67_ASAP7_75t_L g4535 ( 
.A(n_4516),
.Y(n_4535)
);

INVx2_ASAP7_75t_L g4536 ( 
.A(n_4521),
.Y(n_4536)
);

NOR2xp33_ASAP7_75t_L g4537 ( 
.A(n_4516),
.B(n_4081),
.Y(n_4537)
);

AOI21xp5_ASAP7_75t_L g4538 ( 
.A1(n_4516),
.A2(n_4391),
.B(n_4369),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_4516),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4516),
.Y(n_4540)
);

NOR2xp67_ASAP7_75t_L g4541 ( 
.A(n_4529),
.B(n_4307),
.Y(n_4541)
);

NAND4xp25_ASAP7_75t_L g4542 ( 
.A(n_4537),
.B(n_4287),
.C(n_4329),
.D(n_4323),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_L g4543 ( 
.A(n_4531),
.B(n_4309),
.Y(n_4543)
);

AOI22xp33_ASAP7_75t_L g4544 ( 
.A1(n_4533),
.A2(n_4309),
.B1(n_4336),
.B2(n_4326),
.Y(n_4544)
);

NAND2xp5_ASAP7_75t_L g4545 ( 
.A(n_4538),
.B(n_4315),
.Y(n_4545)
);

NOR3xp33_ASAP7_75t_L g4546 ( 
.A(n_4539),
.B(n_4091),
.C(n_4107),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_4525),
.Y(n_4547)
);

AOI211xp5_ASAP7_75t_L g4548 ( 
.A1(n_4527),
.A2(n_4315),
.B(n_4326),
.C(n_4322),
.Y(n_4548)
);

INVx2_ASAP7_75t_L g4549 ( 
.A(n_4526),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_4535),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_4532),
.Y(n_4551)
);

NAND4xp25_ASAP7_75t_L g4552 ( 
.A(n_4528),
.B(n_4329),
.C(n_4336),
.D(n_4322),
.Y(n_4552)
);

NOR2xp33_ASAP7_75t_L g4553 ( 
.A(n_4536),
.B(n_4175),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_L g4554 ( 
.A(n_4534),
.B(n_4363),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_4530),
.Y(n_4555)
);

NOR2xp33_ASAP7_75t_L g4556 ( 
.A(n_4540),
.B(n_4101),
.Y(n_4556)
);

O2A1O1Ixp33_ASAP7_75t_L g4557 ( 
.A1(n_4530),
.A2(n_4261),
.B(n_4364),
.C(n_4316),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4525),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_4525),
.Y(n_4559)
);

INVx1_ASAP7_75t_SL g4560 ( 
.A(n_4525),
.Y(n_4560)
);

NOR3xp33_ASAP7_75t_L g4561 ( 
.A(n_4537),
.B(n_4340),
.C(n_4165),
.Y(n_4561)
);

NAND3xp33_ASAP7_75t_L g4562 ( 
.A(n_4537),
.B(n_4364),
.C(n_4360),
.Y(n_4562)
);

NAND2xp5_ASAP7_75t_SL g4563 ( 
.A(n_4538),
.B(n_4261),
.Y(n_4563)
);

NOR3xp33_ASAP7_75t_L g4564 ( 
.A(n_4537),
.B(n_4281),
.C(n_4366),
.Y(n_4564)
);

NAND5xp2_ASAP7_75t_L g4565 ( 
.A(n_4553),
.B(n_4273),
.C(n_4112),
.D(n_4275),
.E(n_4213),
.Y(n_4565)
);

NAND4xp75_ASAP7_75t_L g4566 ( 
.A(n_4550),
.B(n_4274),
.C(n_4360),
.D(n_4367),
.Y(n_4566)
);

NOR3xp33_ASAP7_75t_L g4567 ( 
.A(n_4556),
.B(n_4549),
.C(n_4547),
.Y(n_4567)
);

NAND2xp5_ASAP7_75t_L g4568 ( 
.A(n_4546),
.B(n_4320),
.Y(n_4568)
);

NOR2xp33_ASAP7_75t_L g4569 ( 
.A(n_4552),
.B(n_4148),
.Y(n_4569)
);

AND2x2_ASAP7_75t_L g4570 ( 
.A(n_4561),
.B(n_4266),
.Y(n_4570)
);

NOR3xp33_ASAP7_75t_L g4571 ( 
.A(n_4558),
.B(n_4161),
.C(n_4152),
.Y(n_4571)
);

AOI21xp33_ASAP7_75t_L g4572 ( 
.A1(n_4551),
.A2(n_4088),
.B(n_4252),
.Y(n_4572)
);

NAND3xp33_ASAP7_75t_L g4573 ( 
.A(n_4555),
.B(n_4367),
.C(n_4325),
.Y(n_4573)
);

NOR2xp33_ASAP7_75t_SL g4574 ( 
.A(n_4560),
.B(n_4155),
.Y(n_4574)
);

AOI211xp5_ASAP7_75t_L g4575 ( 
.A1(n_4541),
.A2(n_4252),
.B(n_4279),
.C(n_4324),
.Y(n_4575)
);

NOR3x1_ASAP7_75t_L g4576 ( 
.A(n_4545),
.B(n_4327),
.C(n_4325),
.Y(n_4576)
);

AOI211xp5_ASAP7_75t_L g4577 ( 
.A1(n_4563),
.A2(n_4559),
.B(n_4543),
.C(n_4562),
.Y(n_4577)
);

NAND3xp33_ASAP7_75t_L g4578 ( 
.A(n_4544),
.B(n_4548),
.C(n_4557),
.Y(n_4578)
);

NAND3xp33_ASAP7_75t_SL g4579 ( 
.A(n_4554),
.B(n_4144),
.C(n_4178),
.Y(n_4579)
);

NOR4xp25_ASAP7_75t_L g4580 ( 
.A(n_4542),
.B(n_4327),
.C(n_4330),
.D(n_4353),
.Y(n_4580)
);

NAND3xp33_ASAP7_75t_L g4581 ( 
.A(n_4564),
.B(n_4330),
.C(n_4355),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_4553),
.B(n_4351),
.Y(n_4582)
);

NOR3xp33_ASAP7_75t_L g4583 ( 
.A(n_4550),
.B(n_4258),
.C(n_4352),
.Y(n_4583)
);

OAI21xp5_ASAP7_75t_SL g4584 ( 
.A1(n_4546),
.A2(n_4334),
.B(n_4220),
.Y(n_4584)
);

NOR4xp25_ASAP7_75t_L g4585 ( 
.A(n_4560),
.B(n_4358),
.C(n_4341),
.D(n_4333),
.Y(n_4585)
);

OAI211xp5_ASAP7_75t_L g4586 ( 
.A1(n_4553),
.A2(n_4274),
.B(n_4352),
.C(n_4220),
.Y(n_4586)
);

NOR4xp25_ASAP7_75t_L g4587 ( 
.A(n_4560),
.B(n_4216),
.C(n_4209),
.D(n_4211),
.Y(n_4587)
);

AOI21xp5_ASAP7_75t_L g4588 ( 
.A1(n_4553),
.A2(n_4155),
.B(n_4216),
.Y(n_4588)
);

OAI21xp5_ASAP7_75t_L g4589 ( 
.A1(n_4553),
.A2(n_4229),
.B(n_4226),
.Y(n_4589)
);

NAND3xp33_ASAP7_75t_L g4590 ( 
.A(n_4556),
.B(n_4334),
.C(n_4274),
.Y(n_4590)
);

INVx2_ASAP7_75t_SL g4591 ( 
.A(n_4551),
.Y(n_4591)
);

NAND2xp5_ASAP7_75t_L g4592 ( 
.A(n_4553),
.B(n_4285),
.Y(n_4592)
);

OAI21xp5_ASAP7_75t_L g4593 ( 
.A1(n_4571),
.A2(n_4226),
.B(n_4334),
.Y(n_4593)
);

NAND2xp5_ASAP7_75t_L g4594 ( 
.A(n_4584),
.B(n_4286),
.Y(n_4594)
);

NOR2x1_ASAP7_75t_L g4595 ( 
.A(n_4578),
.B(n_4274),
.Y(n_4595)
);

AOI22xp5_ASAP7_75t_L g4596 ( 
.A1(n_4574),
.A2(n_4579),
.B1(n_4569),
.B2(n_4583),
.Y(n_4596)
);

NOR2xp33_ASAP7_75t_L g4597 ( 
.A(n_4572),
.B(n_4591),
.Y(n_4597)
);

NAND4xp75_ASAP7_75t_L g4598 ( 
.A(n_4576),
.B(n_4213),
.C(n_4179),
.D(n_4276),
.Y(n_4598)
);

AOI221xp5_ASAP7_75t_L g4599 ( 
.A1(n_4585),
.A2(n_4209),
.B1(n_4211),
.B2(n_4204),
.C(n_4207),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4592),
.Y(n_4600)
);

NOR2x1_ASAP7_75t_L g4601 ( 
.A(n_4573),
.B(n_4301),
.Y(n_4601)
);

BUFx2_ASAP7_75t_L g4602 ( 
.A(n_4570),
.Y(n_4602)
);

AOI21xp5_ASAP7_75t_L g4603 ( 
.A1(n_4568),
.A2(n_4207),
.B(n_4258),
.Y(n_4603)
);

NAND4xp25_ASAP7_75t_L g4604 ( 
.A(n_4567),
.B(n_4277),
.C(n_4251),
.D(n_4276),
.Y(n_4604)
);

AOI22xp5_ASAP7_75t_L g4605 ( 
.A1(n_4588),
.A2(n_4237),
.B1(n_4284),
.B2(n_4240),
.Y(n_4605)
);

INVx1_ASAP7_75t_L g4606 ( 
.A(n_4582),
.Y(n_4606)
);

NAND3xp33_ASAP7_75t_SL g4607 ( 
.A(n_4577),
.B(n_4237),
.C(n_4240),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_4589),
.B(n_4284),
.Y(n_4608)
);

NAND4xp25_ASAP7_75t_SL g4609 ( 
.A(n_4575),
.B(n_4238),
.C(n_4283),
.D(n_4291),
.Y(n_4609)
);

AOI221xp5_ASAP7_75t_L g4610 ( 
.A1(n_4587),
.A2(n_4238),
.B1(n_4283),
.B2(n_4172),
.C(n_4291),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_SL g4611 ( 
.A(n_4580),
.B(n_4224),
.Y(n_4611)
);

NAND4xp25_ASAP7_75t_L g4612 ( 
.A(n_4581),
.B(n_4289),
.C(n_4164),
.D(n_4295),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_4566),
.Y(n_4613)
);

NOR2xp33_ASAP7_75t_L g4614 ( 
.A(n_4590),
.B(n_4289),
.Y(n_4614)
);

NOR3xp33_ASAP7_75t_L g4615 ( 
.A(n_4565),
.B(n_4275),
.C(n_4223),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_SL g4616 ( 
.A(n_4586),
.B(n_4224),
.Y(n_4616)
);

NOR3xp33_ASAP7_75t_SL g4617 ( 
.A(n_4578),
.B(n_4243),
.C(n_4244),
.Y(n_4617)
);

AOI22xp5_ASAP7_75t_L g4618 ( 
.A1(n_4607),
.A2(n_4300),
.B1(n_4280),
.B2(n_4297),
.Y(n_4618)
);

NAND2xp5_ASAP7_75t_L g4619 ( 
.A(n_4593),
.B(n_4300),
.Y(n_4619)
);

AOI321xp33_ASAP7_75t_L g4620 ( 
.A1(n_4595),
.A2(n_4597),
.A3(n_4594),
.B1(n_4601),
.B2(n_4616),
.C(n_4611),
.Y(n_4620)
);

OAI22xp5_ASAP7_75t_L g4621 ( 
.A1(n_4605),
.A2(n_4270),
.B1(n_4243),
.B2(n_4244),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4608),
.Y(n_4622)
);

AOI221xp5_ASAP7_75t_L g4623 ( 
.A1(n_4613),
.A2(n_4270),
.B1(n_4300),
.B2(n_4297),
.C(n_4295),
.Y(n_4623)
);

OAI221xp5_ASAP7_75t_L g4624 ( 
.A1(n_4596),
.A2(n_4614),
.B1(n_4617),
.B2(n_4602),
.C(n_4600),
.Y(n_4624)
);

NAND2xp33_ASAP7_75t_R g4625 ( 
.A(n_4606),
.B(n_459),
.Y(n_4625)
);

NAND2xp33_ASAP7_75t_SL g4626 ( 
.A(n_4609),
.B(n_4297),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_L g4627 ( 
.A(n_4598),
.B(n_4280),
.Y(n_4627)
);

NOR2xp33_ASAP7_75t_R g4628 ( 
.A(n_4615),
.B(n_462),
.Y(n_4628)
);

NAND2xp5_ASAP7_75t_SL g4629 ( 
.A(n_4603),
.B(n_4271),
.Y(n_4629)
);

AND2x2_ASAP7_75t_L g4630 ( 
.A(n_4610),
.B(n_4111),
.Y(n_4630)
);

NAND3xp33_ASAP7_75t_L g4631 ( 
.A(n_4599),
.B(n_4271),
.C(n_4106),
.Y(n_4631)
);

HB1xp67_ASAP7_75t_L g4632 ( 
.A(n_4604),
.Y(n_4632)
);

NOR2x1_ASAP7_75t_L g4633 ( 
.A(n_4612),
.B(n_4280),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_4594),
.Y(n_4634)
);

NOR2x1p5_ASAP7_75t_L g4635 ( 
.A(n_4607),
.B(n_4290),
.Y(n_4635)
);

NOR2x1_ASAP7_75t_L g4636 ( 
.A(n_4624),
.B(n_4263),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_L g4637 ( 
.A(n_4630),
.B(n_4290),
.Y(n_4637)
);

NOR2x1_ASAP7_75t_L g4638 ( 
.A(n_4634),
.B(n_4263),
.Y(n_4638)
);

AND2x4_ASAP7_75t_L g4639 ( 
.A(n_4622),
.B(n_4303),
.Y(n_4639)
);

OAI21xp5_ASAP7_75t_L g4640 ( 
.A1(n_4627),
.A2(n_4223),
.B(n_4290),
.Y(n_4640)
);

OR2x2_ASAP7_75t_L g4641 ( 
.A(n_4631),
.B(n_4263),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_4620),
.Y(n_4642)
);

AOI22xp5_ASAP7_75t_L g4643 ( 
.A1(n_4625),
.A2(n_4303),
.B1(n_4254),
.B2(n_4200),
.Y(n_4643)
);

OR2x2_ASAP7_75t_L g4644 ( 
.A(n_4619),
.B(n_4303),
.Y(n_4644)
);

INVx1_ASAP7_75t_L g4645 ( 
.A(n_4629),
.Y(n_4645)
);

NOR4xp75_ASAP7_75t_L g4646 ( 
.A(n_4628),
.B(n_4254),
.C(n_469),
.D(n_474),
.Y(n_4646)
);

NOR2x1p5_ASAP7_75t_L g4647 ( 
.A(n_4632),
.B(n_4254),
.Y(n_4647)
);

NOR2x1_ASAP7_75t_L g4648 ( 
.A(n_4635),
.B(n_468),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4626),
.Y(n_4649)
);

OA22x2_ASAP7_75t_L g4650 ( 
.A1(n_4621),
.A2(n_4200),
.B1(n_477),
.B2(n_483),
.Y(n_4650)
);

NOR2x1_ASAP7_75t_L g4651 ( 
.A(n_4633),
.B(n_475),
.Y(n_4651)
);

AOI211xp5_ASAP7_75t_L g4652 ( 
.A1(n_4642),
.A2(n_4623),
.B(n_4618),
.C(n_488),
.Y(n_4652)
);

OAI22xp5_ASAP7_75t_L g4653 ( 
.A1(n_4636),
.A2(n_4200),
.B1(n_1425),
.B2(n_1433),
.Y(n_4653)
);

NOR3xp33_ASAP7_75t_L g4654 ( 
.A(n_4645),
.B(n_484),
.C(n_485),
.Y(n_4654)
);

NAND4xp25_ASAP7_75t_L g4655 ( 
.A(n_4648),
.B(n_490),
.C(n_491),
.D(n_492),
.Y(n_4655)
);

OR2x2_ASAP7_75t_L g4656 ( 
.A(n_4641),
.B(n_494),
.Y(n_4656)
);

NAND4xp75_ASAP7_75t_L g4657 ( 
.A(n_4651),
.B(n_499),
.C(n_502),
.D(n_503),
.Y(n_4657)
);

NAND4xp25_ASAP7_75t_L g4658 ( 
.A(n_4649),
.B(n_509),
.C(n_510),
.D(n_513),
.Y(n_4658)
);

NOR5xp2_ASAP7_75t_L g4659 ( 
.A(n_4640),
.B(n_516),
.C(n_520),
.D(n_521),
.E(n_522),
.Y(n_4659)
);

INVx1_ASAP7_75t_L g4660 ( 
.A(n_4637),
.Y(n_4660)
);

NAND4xp25_ASAP7_75t_SL g4661 ( 
.A(n_4644),
.B(n_524),
.C(n_532),
.D(n_1936),
.Y(n_4661)
);

AOI221x1_ASAP7_75t_L g4662 ( 
.A1(n_4646),
.A2(n_1936),
.B1(n_1923),
.B2(n_1902),
.C(n_1892),
.Y(n_4662)
);

NAND4xp75_ASAP7_75t_L g4663 ( 
.A(n_4638),
.B(n_1936),
.C(n_1923),
.D(n_1902),
.Y(n_4663)
);

NOR2x1_ASAP7_75t_L g4664 ( 
.A(n_4647),
.B(n_1443),
.Y(n_4664)
);

NOR3xp33_ASAP7_75t_L g4665 ( 
.A(n_4643),
.B(n_1443),
.C(n_1440),
.Y(n_4665)
);

XNOR2x1_ASAP7_75t_L g4666 ( 
.A(n_4650),
.B(n_1443),
.Y(n_4666)
);

NOR3xp33_ASAP7_75t_L g4667 ( 
.A(n_4639),
.B(n_1443),
.C(n_1440),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4637),
.Y(n_4668)
);

NAND2xp5_ASAP7_75t_L g4669 ( 
.A(n_4642),
.B(n_1440),
.Y(n_4669)
);

HB1xp67_ASAP7_75t_L g4670 ( 
.A(n_4657),
.Y(n_4670)
);

AOI221xp5_ASAP7_75t_SL g4671 ( 
.A1(n_4652),
.A2(n_1936),
.B1(n_1923),
.B2(n_1902),
.C(n_1892),
.Y(n_4671)
);

NOR2xp33_ASAP7_75t_R g4672 ( 
.A(n_4661),
.B(n_4656),
.Y(n_4672)
);

CKINVDCx5p33_ASAP7_75t_R g4673 ( 
.A(n_4660),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_4666),
.Y(n_4674)
);

OR2x2_ASAP7_75t_L g4675 ( 
.A(n_4655),
.B(n_1433),
.Y(n_4675)
);

CKINVDCx5p33_ASAP7_75t_R g4676 ( 
.A(n_4668),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_4669),
.Y(n_4677)
);

NAND4xp75_ASAP7_75t_L g4678 ( 
.A(n_4662),
.B(n_1923),
.C(n_1902),
.D(n_1892),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_4664),
.Y(n_4679)
);

CKINVDCx16_ASAP7_75t_R g4680 ( 
.A(n_4658),
.Y(n_4680)
);

AOI221xp5_ASAP7_75t_L g4681 ( 
.A1(n_4665),
.A2(n_1892),
.B1(n_1881),
.B2(n_1860),
.C(n_1838),
.Y(n_4681)
);

INVx1_ASAP7_75t_SL g4682 ( 
.A(n_4663),
.Y(n_4682)
);

OAI22xp33_ASAP7_75t_L g4683 ( 
.A1(n_4680),
.A2(n_4653),
.B1(n_4659),
.B2(n_4654),
.Y(n_4683)
);

OAI221xp5_ASAP7_75t_L g4684 ( 
.A1(n_4671),
.A2(n_4667),
.B1(n_1892),
.B2(n_1881),
.C(n_1860),
.Y(n_4684)
);

AOI221xp5_ASAP7_75t_L g4685 ( 
.A1(n_4682),
.A2(n_1881),
.B1(n_1860),
.B2(n_1838),
.C(n_1832),
.Y(n_4685)
);

AOI22xp33_ASAP7_75t_SL g4686 ( 
.A1(n_4673),
.A2(n_1881),
.B1(n_1860),
.B2(n_1838),
.Y(n_4686)
);

INVx2_ASAP7_75t_L g4687 ( 
.A(n_4675),
.Y(n_4687)
);

AND2x2_ASAP7_75t_L g4688 ( 
.A(n_4670),
.B(n_1881),
.Y(n_4688)
);

INVx2_ASAP7_75t_L g4689 ( 
.A(n_4678),
.Y(n_4689)
);

AOI22xp5_ASAP7_75t_L g4690 ( 
.A1(n_4683),
.A2(n_4676),
.B1(n_4674),
.B2(n_4677),
.Y(n_4690)
);

AOI22xp5_ASAP7_75t_SL g4691 ( 
.A1(n_4688),
.A2(n_4689),
.B1(n_4679),
.B2(n_4687),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4686),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4684),
.Y(n_4693)
);

AOI22xp5_ASAP7_75t_L g4694 ( 
.A1(n_4685),
.A2(n_4681),
.B1(n_4672),
.B2(n_1860),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4688),
.Y(n_4695)
);

OAI22x1_ASAP7_75t_L g4696 ( 
.A1(n_4689),
.A2(n_1299),
.B1(n_1308),
.B2(n_1322),
.Y(n_4696)
);

INVx2_ASAP7_75t_SL g4697 ( 
.A(n_4691),
.Y(n_4697)
);

NAND4xp25_ASAP7_75t_L g4698 ( 
.A(n_4690),
.B(n_1838),
.C(n_1832),
.D(n_1830),
.Y(n_4698)
);

NAND3x1_ASAP7_75t_L g4699 ( 
.A(n_4695),
.B(n_1838),
.C(n_1832),
.Y(n_4699)
);

NOR4xp25_ASAP7_75t_L g4700 ( 
.A(n_4692),
.B(n_1832),
.C(n_1830),
.D(n_1827),
.Y(n_4700)
);

AOI22xp5_ASAP7_75t_L g4701 ( 
.A1(n_4693),
.A2(n_1832),
.B1(n_1830),
.B2(n_1827),
.Y(n_4701)
);

XNOR2xp5_ASAP7_75t_L g4702 ( 
.A(n_4694),
.B(n_1830),
.Y(n_4702)
);

AO22x2_ASAP7_75t_L g4703 ( 
.A1(n_4697),
.A2(n_4696),
.B1(n_1830),
.B2(n_1827),
.Y(n_4703)
);

OAI22xp33_ASAP7_75t_L g4704 ( 
.A1(n_4701),
.A2(n_1827),
.B1(n_1824),
.B2(n_1822),
.Y(n_4704)
);

HB1xp67_ASAP7_75t_L g4705 ( 
.A(n_4702),
.Y(n_4705)
);

AOI21x1_ASAP7_75t_L g4706 ( 
.A1(n_4699),
.A2(n_1827),
.B(n_1824),
.Y(n_4706)
);

AND3x1_ASAP7_75t_L g4707 ( 
.A(n_4700),
.B(n_1793),
.C(n_1822),
.Y(n_4707)
);

OAI321xp33_ASAP7_75t_L g4708 ( 
.A1(n_4704),
.A2(n_4698),
.A3(n_1824),
.B1(n_1822),
.B2(n_1821),
.C(n_1817),
.Y(n_4708)
);

HB1xp67_ASAP7_75t_L g4709 ( 
.A(n_4706),
.Y(n_4709)
);

BUFx2_ASAP7_75t_L g4710 ( 
.A(n_4707),
.Y(n_4710)
);

NAND3xp33_ASAP7_75t_L g4711 ( 
.A(n_4705),
.B(n_1824),
.C(n_1822),
.Y(n_4711)
);

AOI21xp5_ASAP7_75t_L g4712 ( 
.A1(n_4710),
.A2(n_4703),
.B(n_1824),
.Y(n_4712)
);

INVxp33_ASAP7_75t_L g4713 ( 
.A(n_4709),
.Y(n_4713)
);

OAI21xp5_ASAP7_75t_SL g4714 ( 
.A1(n_4711),
.A2(n_1822),
.B(n_1821),
.Y(n_4714)
);

NAND2xp5_ASAP7_75t_L g4715 ( 
.A(n_4708),
.B(n_1821),
.Y(n_4715)
);

AOI22xp5_ASAP7_75t_L g4716 ( 
.A1(n_4711),
.A2(n_1821),
.B1(n_1817),
.B2(n_1793),
.Y(n_4716)
);

OA21x2_ASAP7_75t_L g4717 ( 
.A1(n_4712),
.A2(n_1821),
.B(n_1817),
.Y(n_4717)
);

AOI22xp5_ASAP7_75t_L g4718 ( 
.A1(n_4713),
.A2(n_1817),
.B1(n_1793),
.B2(n_1784),
.Y(n_4718)
);

OAI21x1_ASAP7_75t_L g4719 ( 
.A1(n_4715),
.A2(n_1817),
.B(n_1793),
.Y(n_4719)
);

AOI22x1_ASAP7_75t_L g4720 ( 
.A1(n_4714),
.A2(n_1793),
.B1(n_1784),
.B2(n_1778),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_4716),
.Y(n_4721)
);

OR2x2_ASAP7_75t_L g4722 ( 
.A(n_4713),
.B(n_1784),
.Y(n_4722)
);

XOR2xp5_ASAP7_75t_L g4723 ( 
.A(n_4713),
.B(n_1784),
.Y(n_4723)
);

INVx1_ASAP7_75t_L g4724 ( 
.A(n_4715),
.Y(n_4724)
);

AOI21xp33_ASAP7_75t_SL g4725 ( 
.A1(n_4713),
.A2(n_1784),
.B(n_1778),
.Y(n_4725)
);

O2A1O1Ixp33_ASAP7_75t_L g4726 ( 
.A1(n_4713),
.A2(n_1767),
.B(n_1757),
.C(n_1778),
.Y(n_4726)
);

OAI22xp5_ASAP7_75t_L g4727 ( 
.A1(n_4723),
.A2(n_1778),
.B1(n_1767),
.B2(n_1757),
.Y(n_4727)
);

OAI22xp33_ASAP7_75t_L g4728 ( 
.A1(n_4718),
.A2(n_1778),
.B1(n_1767),
.B2(n_1757),
.Y(n_4728)
);

OAI22xp33_ASAP7_75t_L g4729 ( 
.A1(n_4722),
.A2(n_1767),
.B1(n_1308),
.B2(n_1322),
.Y(n_4729)
);

AOI22xp5_ASAP7_75t_L g4730 ( 
.A1(n_4724),
.A2(n_1299),
.B1(n_1308),
.B2(n_1322),
.Y(n_4730)
);

AOI22xp5_ASAP7_75t_L g4731 ( 
.A1(n_4721),
.A2(n_1299),
.B1(n_1308),
.B2(n_1322),
.Y(n_4731)
);

AOI22xp5_ASAP7_75t_L g4732 ( 
.A1(n_4717),
.A2(n_1299),
.B1(n_1346),
.B2(n_1376),
.Y(n_4732)
);

OAI22xp5_ASAP7_75t_L g4733 ( 
.A1(n_4720),
.A2(n_4725),
.B1(n_4726),
.B2(n_4719),
.Y(n_4733)
);

OAI22xp5_ASAP7_75t_L g4734 ( 
.A1(n_4723),
.A2(n_1346),
.B1(n_1376),
.B2(n_1394),
.Y(n_4734)
);

AOI22xp5_ASAP7_75t_L g4735 ( 
.A1(n_4723),
.A2(n_1346),
.B1(n_1376),
.B2(n_1394),
.Y(n_4735)
);

OAI22xp33_ASAP7_75t_L g4736 ( 
.A1(n_4718),
.A2(n_1346),
.B1(n_1376),
.B2(n_1394),
.Y(n_4736)
);

AOI21xp5_ASAP7_75t_L g4737 ( 
.A1(n_4733),
.A2(n_1394),
.B(n_1396),
.Y(n_4737)
);

AOI221xp5_ASAP7_75t_L g4738 ( 
.A1(n_4728),
.A2(n_1396),
.B1(n_1437),
.B2(n_1438),
.C(n_1501),
.Y(n_4738)
);

AND2x2_ASAP7_75t_L g4739 ( 
.A(n_4732),
.B(n_1396),
.Y(n_4739)
);

OR2x6_ASAP7_75t_L g4740 ( 
.A(n_4734),
.B(n_4727),
.Y(n_4740)
);

NAND2xp5_ASAP7_75t_SL g4741 ( 
.A(n_4729),
.B(n_1396),
.Y(n_4741)
);

NAND2xp5_ASAP7_75t_SL g4742 ( 
.A(n_4735),
.B(n_1437),
.Y(n_4742)
);

NAND2xp5_ASAP7_75t_L g4743 ( 
.A(n_4736),
.B(n_1437),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4739),
.Y(n_4744)
);

OAI22xp33_ASAP7_75t_L g4745 ( 
.A1(n_4740),
.A2(n_4731),
.B1(n_4730),
.B2(n_1437),
.Y(n_4745)
);

HB1xp67_ASAP7_75t_L g4746 ( 
.A(n_4740),
.Y(n_4746)
);

AOI221x1_ASAP7_75t_L g4747 ( 
.A1(n_4744),
.A2(n_4737),
.B1(n_4743),
.B2(n_4742),
.C(n_4738),
.Y(n_4747)
);

AOI21xp5_ASAP7_75t_L g4748 ( 
.A1(n_4747),
.A2(n_4746),
.B(n_4745),
.Y(n_4748)
);

AOI211xp5_ASAP7_75t_L g4749 ( 
.A1(n_4748),
.A2(n_4741),
.B(n_1438),
.C(n_1483),
.Y(n_4749)
);


endmodule