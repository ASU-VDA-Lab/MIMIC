module real_jpeg_23725_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_1),
.A2(n_40),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_49),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_1),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_1),
.A2(n_49),
.B1(n_62),
.B2(n_63),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_67),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_67),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_2),
.A2(n_67),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_3),
.A2(n_55),
.B1(n_56),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_3),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_171),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_171),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_3),
.A2(n_33),
.B1(n_50),
.B2(n_171),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_4),
.A2(n_32),
.B1(n_40),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_4),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_4),
.A2(n_62),
.B1(n_63),
.B2(n_151),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_4),
.A2(n_55),
.B1(n_56),
.B2(n_151),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_151),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_6),
.A2(n_55),
.B1(n_56),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_6),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_6),
.A2(n_62),
.B1(n_63),
.B2(n_180),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_180),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_6),
.A2(n_38),
.B1(n_180),
.B2(n_290),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_8),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_39),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_9),
.A2(n_39),
.B1(n_55),
.B2(n_56),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_9),
.A2(n_39),
.B1(n_62),
.B2(n_63),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_10),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_10),
.A2(n_35),
.B1(n_55),
.B2(n_56),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_10),
.A2(n_35),
.B1(n_62),
.B2(n_63),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_11),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_11),
.A2(n_58),
.B(n_63),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_11),
.B(n_88),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_11),
.A2(n_108),
.B1(n_112),
.B2(n_198),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_11),
.A2(n_26),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_11),
.B(n_47),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_15),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_15),
.Y(n_112)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_15),
.Y(n_146)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_15),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_129),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_89),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_19),
.B(n_89),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_83),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_44),
.B1(n_81),
.B2(n_82),
.Y(n_20)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_52),
.C(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_21),
.A2(n_81),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_30),
.B(n_36),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_22),
.B(n_43),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_22),
.A2(n_42),
.B1(n_150),
.B2(n_289),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_23),
.A2(n_24),
.B1(n_32),
.B2(n_40),
.Y(n_43)
);

OAI32xp33_ASAP7_75t_L g258 ( 
.A1(n_23),
.A2(n_27),
.A3(n_33),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_24),
.B(n_26),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_26),
.A2(n_27),
.B1(n_73),
.B2(n_74),
.Y(n_78)
);

OAI32xp33_ASAP7_75t_L g221 ( 
.A1(n_26),
.A2(n_56),
.A3(n_73),
.B1(n_213),
.B2(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_27),
.B(n_168),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g276 ( 
.A1(n_32),
.A2(n_168),
.B(n_259),
.Y(n_276)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_33),
.Y(n_124)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_41),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_37),
.B(n_47),
.Y(n_126)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_38),
.Y(n_290)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_41),
.A2(n_47),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_41),
.A2(n_47),
.B1(n_277),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_42),
.A2(n_122),
.B(n_126),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_42),
.A2(n_150),
.B(n_152),
.Y(n_149)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_51),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_47),
.B(n_123),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_68),
.B1(n_69),
.B2(n_80),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_52),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_80),
.B1(n_84),
.B2(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_65),
.B(n_66),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_53),
.B(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_53),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_53),
.A2(n_65),
.B1(n_170),
.B2(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_53),
.A2(n_65),
.B1(n_179),
.B2(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_53),
.A2(n_66),
.B(n_119),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_61),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_56),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_55),
.B(n_74),
.Y(n_222)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_SL g172 ( 
.A1(n_56),
.A2(n_60),
.B(n_168),
.C(n_173),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_61),
.B(n_100),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_61),
.A2(n_116),
.B1(n_117),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_61),
.A2(n_116),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_61),
.B(n_168),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_61),
.A2(n_98),
.B(n_148),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_62),
.B(n_202),
.Y(n_201)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_66),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_71),
.A2(n_77),
.B(n_273),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_72),
.A2(n_76),
.B(n_103),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_72),
.A2(n_211),
.B1(n_214),
.B2(n_215),
.Y(n_210)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_75),
.A2(n_87),
.B(n_214),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_85),
.B1(n_88),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_77),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_77),
.A2(n_88),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_77),
.A2(n_88),
.B1(n_238),
.B2(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.C(n_104),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_90),
.A2(n_94),
.B1(n_95),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_95),
.A2(n_96),
.B(n_101),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_101),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_97),
.A2(n_116),
.B(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_120),
.B(n_121),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_106),
.B1(n_133),
.B2(n_135),
.Y(n_132)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_115),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_120),
.B1(n_121),
.B2(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_107),
.A2(n_115),
.B1(n_120),
.B2(n_323),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_112),
.B(n_113),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_108),
.A2(n_144),
.B(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_108),
.A2(n_146),
.B1(n_188),
.B2(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_108),
.A2(n_113),
.B(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_108),
.A2(n_224),
.B(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_109),
.B(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_109),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_109),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.Y(n_261)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_112),
.B(n_168),
.Y(n_202)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_115),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_124),
.B(n_168),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_157),
.B(n_338),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_154),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_131),
.B(n_154),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.C(n_138),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_132),
.A2(n_136),
.B1(n_137),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_132),
.Y(n_327)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_138),
.B(n_326),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_149),
.C(n_153),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_139),
.A2(n_140),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_147),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_141),
.B(n_147),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_142),
.A2(n_191),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_143),
.B(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_149),
.B(n_153),
.Y(n_320)
);

AOI311xp33_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_316),
.A3(n_328),
.B(n_332),
.C(n_333),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_279),
.C(n_311),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_253),
.B(n_278),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_231),
.B(n_252),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_206),
.B(n_230),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_184),
.B(n_205),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_174),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_164),
.B(n_174),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_172),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_165),
.A2(n_166),
.B1(n_172),
.B2(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_172),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_182),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_181),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_181),
.C(n_182),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_178),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_183),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_194),
.B(n_204),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_186),
.B(n_192),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_191),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_199),
.B(n_203),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_196),
.B(n_197),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_207),
.B(n_208),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_220),
.B1(n_228),
.B2(n_229),
.Y(n_208)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_209)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_215),
.Y(n_237)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_216),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_219),
.C(n_228),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_223),
.Y(n_247)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_232),
.B(n_233),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_245),
.B2(n_246),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_248),
.C(n_250),
.Y(n_254)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_241),
.C(n_242),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_246)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_247),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_248),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_254),
.B(n_255),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_270),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_257),
.B(n_269),
.C(n_270),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_261),
.B1(n_265),
.B2(n_266),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_258),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_265),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_261),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_264),
.Y(n_294)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_275),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_274),
.C(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI21xp33_ASAP7_75t_L g334 ( 
.A1(n_280),
.A2(n_335),
.B(n_336),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_296),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_281),
.B(n_296),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_291),
.C(n_292),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_282),
.A2(n_283),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_286),
.C(n_287),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_291),
.B(n_292),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_295),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_296)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_306),
.B2(n_307),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_298),
.B(n_307),
.C(n_310),
.Y(n_330)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_302),
.B2(n_305),
.Y(n_299)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_300),
.Y(n_305)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_304),
.C(n_305),
.Y(n_324)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_308),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_313),
.Y(n_335)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

O2A1O1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_317),
.A2(n_329),
.B(n_334),
.C(n_337),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_325),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_325),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.C(n_324),
.Y(n_318)
);

FAx1_ASAP7_75t_SL g331 ( 
.A(n_319),
.B(n_322),
.CI(n_324),
.CON(n_331),
.SN(n_331)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_330),
.B(n_331),
.Y(n_337)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_331),
.Y(n_339)
);


endmodule