module real_jpeg_4367_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_1),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_2),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_2),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_2),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_2),
.B(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_2),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_2),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_2),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_3),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_3),
.B(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_4),
.B(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_4),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_4),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_4),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_4),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_4),
.B(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_5),
.A2(n_75),
.B(n_77),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_5),
.B(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_5),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_5),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_5),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_5),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_5),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_5),
.B(n_299),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_6),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_6),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_6),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_6),
.B(n_235),
.Y(n_234)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_8),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_8),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_8),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_8),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_8),
.B(n_288),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_8),
.B(n_323),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_9),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_9),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_9),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g299 ( 
.A(n_9),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_10),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_10),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_10),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_10),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_10),
.B(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_10),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_10),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_10),
.B(n_340),
.Y(n_339)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_12),
.Y(n_76)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_12),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_12),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_12),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_13),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_13),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_14),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_14),
.Y(n_288)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_14),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_15),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_15),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_15),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_15),
.B(n_140),
.Y(n_149)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_15),
.B(n_185),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_15),
.B(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_214),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_213),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_170),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_20),
.B(n_170),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_112),
.C(n_144),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_21),
.B(n_112),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_72),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_22),
.B(n_73),
.C(n_88),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_43),
.C(n_58),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_24),
.B(n_59),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_25),
.B(n_131),
.C(n_132),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_29),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_37),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_31),
.Y(n_132)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_35),
.Y(n_261)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_36),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_36),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_37),
.Y(n_131)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_41),
.Y(n_137)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_42),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_42),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_43),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_49),
.C(n_54),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_44),
.A2(n_45),
.B1(n_54),
.B2(n_55),
.Y(n_147)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_49),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g302 ( 
.A(n_53),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.C(n_68),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_60),
.A2(n_68),
.B1(n_178),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_60),
.Y(n_224)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_63),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_64),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_68),
.A2(n_174),
.B1(n_178),
.B2(n_179),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_68),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_88),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_81),
.C(n_85),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_74),
.B(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_74),
.A2(n_77),
.B(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_81),
.B(n_85),
.Y(n_169)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_83),
.B(n_227),
.Y(n_306)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_98),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_93),
.B1(n_96),
.B2(n_97),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_93),
.B(n_96),
.C(n_98),
.Y(n_200)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_95),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_105),
.C(n_110),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_99),
.A2(n_100),
.B1(n_110),
.B2(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_99),
.A2(n_100),
.B1(n_183),
.B2(n_184),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_100),
.B(n_184),
.Y(n_232)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_104),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_105),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_109),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_110),
.Y(n_167)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_129),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_114),
.B(n_130),
.C(n_133),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_121),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_116),
.B(n_123),
.C(n_126),
.Y(n_211)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_128),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_122),
.A2(n_123),
.B1(n_159),
.B2(n_160),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_159),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_124),
.Y(n_295)
);

INVx8_ASAP7_75t_L g317 ( 
.A(n_124),
.Y(n_317)
);

BUFx8_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g325 ( 
.A(n_125),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_126),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_126),
.A2(n_128),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_126),
.A2(n_128),
.B1(n_301),
.B2(n_303),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_126),
.B(n_303),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_139),
.C(n_141),
.Y(n_181)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_144),
.B(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_163),
.C(n_168),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_145),
.B(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_157),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_146),
.B(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_148),
.A2(n_157),
.B1(n_158),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_148),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.C(n_154),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_149),
.A2(n_154),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_149),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_150),
.B(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_154),
.Y(n_254)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_156),
.Y(n_209)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_163),
.B(n_168),
.Y(n_220)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_212),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_197),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_180),
.Y(n_172)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_175),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_187),
.B2(n_188),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_196),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_211),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_210),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_274),
.B(n_369),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_246),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_217),
.A2(n_371),
.B(n_372),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_244),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_218),
.B(n_244),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.C(n_242),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_219),
.B(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_221),
.B(n_242),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.C(n_230),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_225),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.C(n_236),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_231),
.A2(n_232),
.B1(n_357),
.B2(n_358),
.Y(n_356)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_357)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_272),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_247),
.B(n_272),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.C(n_269),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_248),
.B(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_250),
.B(n_269),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_255),
.C(n_267),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_251),
.B(n_360),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_255),
.A2(n_267),
.B1(n_268),
.B2(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_255),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.C(n_262),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_256),
.A2(n_257),
.B1(n_262),
.B2(n_263),
.Y(n_349)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_259),
.B(n_349),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_261),
.Y(n_310)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_364),
.B(n_368),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_351),
.B(n_363),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_335),
.B(n_350),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_311),
.B(n_334),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_304),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_279),
.B(n_304),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_291),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_280),
.B(n_292),
.C(n_300),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_286),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_281),
.B(n_287),
.C(n_289),
.Y(n_347)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_300),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_296),
.Y(n_305)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.C(n_307),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_331),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_306),
.Y(n_332)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_328),
.B(n_333),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_321),
.B(n_327),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_320),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_320),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_318),
.Y(n_329)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_326),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_337),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_346),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_338),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_338),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_347),
.C(n_348),
.Y(n_362)
);

FAx1_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_344),
.CI(n_345),
.CON(n_338),
.SN(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_362),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_362),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_359),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_356),
.C(n_359),
.Y(n_365)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_357),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_365),
.B(n_366),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);


endmodule