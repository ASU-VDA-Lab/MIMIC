module fake_jpeg_19473_n_130 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_4),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_21),
.Y(n_33)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_17),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

AOI21xp33_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_0),
.B(n_1),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_37),
.Y(n_45)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_14),
.Y(n_52)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_52),
.B(n_55),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_33),
.B(n_24),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_71),
.B(n_1),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_33),
.B1(n_26),
.B2(n_24),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_48),
.B1(n_17),
.B2(n_2),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_13),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_58),
.C(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_63),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_68),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_18),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_70),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_18),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_26),
.B(n_15),
.C(n_14),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_39),
.B(n_7),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_72),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_7),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_73),
.Y(n_83)
);

AND2x6_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_77),
.Y(n_91)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_85),
.B(n_73),
.Y(n_92)
);

CKINVDCx10_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_1),
.B1(n_2),
.B2(n_11),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_93),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_64),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_95),
.B(n_99),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_52),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_85),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_64),
.B1(n_55),
.B2(n_88),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_57),
.B1(n_68),
.B2(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_72),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_80),
.C(n_86),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_103),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_86),
.C(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_94),
.Y(n_113)
);

OAI322xp33_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_78),
.A3(n_83),
.B1(n_93),
.B2(n_63),
.C1(n_61),
.C2(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_100),
.B(n_70),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_92),
.B(n_96),
.C(n_81),
.D(n_98),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_111),
.B(n_112),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_89),
.B1(n_83),
.B2(n_51),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_115),
.B(n_119),
.Y(n_122)
);

AOI31xp33_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_111),
.A3(n_109),
.B(n_71),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_123),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_121),
.B(n_66),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_109),
.B(n_90),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_84),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_66),
.C(n_60),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_60),
.B(n_2),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_128),
.C(n_126),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_84),
.Y(n_130)
);


endmodule