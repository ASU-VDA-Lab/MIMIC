module fake_jpeg_5498_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_34),
.B(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_8),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_40),
.Y(n_55)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx2_ASAP7_75t_SL g60 ( 
.A(n_36),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_27),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_44),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_17),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_17),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_19),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_56),
.Y(n_94)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_54),
.A2(n_65),
.B1(n_66),
.B2(n_36),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_25),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_24),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_61),
.B(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_22),
.B1(n_18),
.B2(n_24),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_24),
.B1(n_37),
.B2(n_17),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_36),
.A2(n_22),
.B1(n_33),
.B2(n_18),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_36),
.A2(n_22),
.B1(n_33),
.B2(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_68),
.B(n_51),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_42),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_76),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_19),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_36),
.B1(n_40),
.B2(n_44),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_80),
.B(n_62),
.C(n_79),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_68),
.B(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_29),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_79),
.B(n_37),
.Y(n_110)
);

NAND2x1_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_36),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_37),
.B(n_34),
.C(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_81),
.B(n_87),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_74),
.B1(n_94),
.B2(n_72),
.Y(n_100)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_83),
.Y(n_123)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_84),
.A2(n_91),
.B1(n_95),
.B2(n_96),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_33),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_57),
.A2(n_43),
.B1(n_39),
.B2(n_26),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_58),
.B1(n_67),
.B2(n_54),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_112),
.B1(n_72),
.B2(n_75),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_100),
.A2(n_107),
.B1(n_98),
.B2(n_121),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_52),
.B1(n_50),
.B2(n_45),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_119),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_55),
.C(n_39),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_89),
.C(n_75),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_43),
.B1(n_44),
.B2(n_40),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_108),
.A2(n_124),
.B(n_90),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_R g109 ( 
.A(n_94),
.B(n_55),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_110),
.B(n_113),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_81),
.A2(n_43),
.B1(n_29),
.B2(n_20),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_80),
.A2(n_20),
.B1(n_29),
.B2(n_49),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_73),
.B(n_46),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_76),
.B(n_49),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_20),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_88),
.B(n_59),
.Y(n_146)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_39),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_43),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_43),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_145),
.B1(n_108),
.B2(n_113),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_75),
.B1(n_87),
.B2(n_96),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_137),
.B1(n_138),
.B2(n_149),
.Y(n_154)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_134),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_136),
.Y(n_176)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_86),
.B1(n_85),
.B2(n_87),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_85),
.B1(n_87),
.B2(n_71),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_142),
.C(n_150),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_95),
.B1(n_84),
.B2(n_83),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_105),
.B(n_106),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_123),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_108),
.A2(n_90),
.B1(n_88),
.B2(n_92),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_110),
.Y(n_159)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

OAI22x1_ASAP7_75t_L g149 ( 
.A1(n_109),
.A2(n_39),
.B1(n_59),
.B2(n_53),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_39),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_100),
.B(n_23),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_152),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_98),
.B(n_23),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_153),
.A2(n_157),
.B1(n_129),
.B2(n_135),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_156),
.A2(n_163),
.B(n_166),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_143),
.A2(n_111),
.B1(n_105),
.B2(n_99),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_162),
.B(n_167),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_118),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_115),
.A3(n_116),
.B1(n_124),
.B2(n_111),
.C1(n_117),
.C2(n_118),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_169),
.C(n_170),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_117),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_120),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_177),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_104),
.C(n_114),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_124),
.C(n_39),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_178),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_124),
.B(n_27),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_172),
.A2(n_173),
.B1(n_23),
.B2(n_32),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_27),
.B(n_39),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_147),
.A2(n_92),
.B(n_59),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_92),
.C(n_53),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_32),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_53),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_179),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_181),
.B(n_183),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_189),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_126),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_198),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_188),
.A2(n_163),
.B1(n_154),
.B2(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_176),
.A2(n_130),
.B1(n_151),
.B2(n_127),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_192),
.B1(n_193),
.B2(n_199),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_175),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_191),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_157),
.A2(n_127),
.B1(n_144),
.B2(n_136),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_148),
.B1(n_131),
.B2(n_128),
.Y(n_193)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_179),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_179),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_174),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_197),
.B(n_206),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_166),
.A2(n_32),
.B1(n_28),
.B2(n_26),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_128),
.B1(n_32),
.B2(n_28),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_200),
.A2(n_208),
.B1(n_167),
.B2(n_162),
.Y(n_225)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_154),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_172),
.B1(n_175),
.B2(n_156),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_209),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_187),
.Y(n_211)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_212),
.B(n_228),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_155),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_222),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_155),
.C(n_178),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_220),
.C(n_226),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_191),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_219),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_177),
.C(n_170),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_159),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_169),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_204),
.Y(n_251)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_225),
.A2(n_183),
.B1(n_198),
.B2(n_203),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_163),
.C(n_28),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_28),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_185),
.C(n_190),
.Y(n_242)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_231),
.B(n_188),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_184),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_186),
.B1(n_196),
.B2(n_181),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_236),
.A2(n_234),
.B1(n_216),
.B2(n_221),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_199),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_237),
.A2(n_250),
.B1(n_257),
.B2(n_224),
.Y(n_273)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_230),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_245),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_248),
.C(n_254),
.Y(n_266)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_223),
.B(n_182),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_251),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_189),
.C(n_186),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_212),
.B(n_23),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_257),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_195),
.C(n_26),
.Y(n_254)
);

INVxp33_ASAP7_75t_SL g255 ( 
.A(n_211),
.Y(n_255)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_26),
.C(n_16),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_214),
.C(n_232),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_214),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_257)
);

NOR3xp33_ASAP7_75t_SL g258 ( 
.A(n_237),
.B(n_252),
.C(n_255),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_262),
.Y(n_286)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

XNOR2x1_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_226),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_270),
.Y(n_287)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_269),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_267),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_243),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_227),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_274),
.C(n_16),
.Y(n_284)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_232),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_8),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_215),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_276),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_229),
.B1(n_225),
.B2(n_254),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_258),
.A2(n_240),
.B1(n_234),
.B2(n_224),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_278),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_280),
.A2(n_281),
.B1(n_292),
.B2(n_288),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_239),
.B1(n_256),
.B2(n_210),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_239),
.B1(n_249),
.B2(n_16),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_282),
.B(n_290),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_293),
.C(n_272),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_289),
.A2(n_10),
.B(n_14),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_8),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_271),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_0),
.C(n_1),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_274),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_297),
.C(n_300),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_268),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_296),
.B(n_299),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_291),
.B(n_267),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_307),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_286),
.B(n_266),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_259),
.C(n_263),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_301),
.B(n_302),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_281),
.B(n_259),
.Y(n_302)
);

INVxp33_ASAP7_75t_SL g304 ( 
.A(n_285),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_292),
.B(n_283),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_9),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_305),
.B(n_306),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_10),
.Y(n_306)
);

NAND3xp33_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_287),
.C(n_293),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_309),
.A2(n_310),
.B(n_311),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_279),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_15),
.C(n_13),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_300),
.C(n_13),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_15),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_3),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_1),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_317),
.A2(n_10),
.B(n_15),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_324),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_320),
.B(n_321),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_13),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_318),
.A2(n_308),
.B(n_312),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_322),
.A2(n_327),
.B(n_11),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_4),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_318),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_SL g326 ( 
.A1(n_313),
.A2(n_3),
.B(n_4),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_326),
.A2(n_12),
.B1(n_6),
.B2(n_7),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_11),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_325),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_SL g334 ( 
.A(n_328),
.B(n_326),
.Y(n_334)
);

NOR3xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_331),
.C(n_332),
.Y(n_335)
);

NOR4xp25_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_329),
.C(n_333),
.D(n_12),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_335),
.B(n_6),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_7),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_5),
.C(n_6),
.Y(n_339)
);


endmodule