module fake_jpeg_25845_n_379 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_379);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_379;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_50),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_28),
.B1(n_19),
.B2(n_26),
.Y(n_68)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_57),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_61),
.Y(n_102)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_13),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_30),
.B(n_13),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_21),
.Y(n_96)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_68),
.A2(n_87),
.B1(n_52),
.B2(n_51),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_73),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_43),
.B(n_30),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_72),
.B(n_96),
.Y(n_135)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_40),
.A2(n_28),
.B1(n_21),
.B2(n_23),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_75),
.A2(n_104),
.B1(n_106),
.B2(n_108),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_42),
.A2(n_28),
.B1(n_26),
.B2(n_23),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_76),
.Y(n_115)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_29),
.B1(n_32),
.B2(n_16),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

BUFx16f_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_39),
.Y(n_129)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_60),
.A2(n_37),
.B1(n_36),
.B2(n_33),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_65),
.A2(n_37),
.B1(n_36),
.B2(n_33),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_107),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_54),
.A2(n_25),
.B1(n_24),
.B2(n_29),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_84),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_111),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_49),
.B(n_53),
.C(n_46),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_112),
.A2(n_120),
.B1(n_132),
.B2(n_90),
.Y(n_162)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_114),
.B(n_137),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_84),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_138),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_109),
.A2(n_25),
.B1(n_29),
.B2(n_12),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_67),
.B1(n_16),
.B2(n_32),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_93),
.A2(n_25),
.B1(n_24),
.B2(n_32),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_122),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_16),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_123),
.B(n_125),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_124),
.A2(n_131),
.B1(n_127),
.B2(n_126),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_47),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_127),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_47),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_93),
.A2(n_47),
.B1(n_55),
.B2(n_45),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_83),
.A2(n_52),
.B1(n_51),
.B2(n_12),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_12),
.A3(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_148),
.B(n_7),
.C(n_9),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_L g134 ( 
.A1(n_83),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_140),
.B1(n_7),
.B2(n_9),
.Y(n_170)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_80),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_78),
.B(n_11),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_139),
.B(n_141),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_89),
.A2(n_0),
.B1(n_1),
.B2(n_6),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_80),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_94),
.A2(n_10),
.B1(n_7),
.B2(n_8),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_146),
.B1(n_150),
.B2(n_81),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_99),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_145),
.B(n_90),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_97),
.A2(n_10),
.B1(n_7),
.B2(n_8),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_6),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_149),
.Y(n_184)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_108),
.A2(n_105),
.A3(n_86),
.B1(n_88),
.B2(n_97),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_82),
.B(n_6),
.Y(n_149)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_159),
.Y(n_203)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_160),
.B(n_165),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_137),
.B(n_114),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_162),
.A2(n_167),
.B1(n_170),
.B2(n_178),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_70),
.C(n_101),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_181),
.C(n_156),
.Y(n_213)
);

AO22x1_ASAP7_75t_L g164 ( 
.A1(n_112),
.A2(n_81),
.B1(n_86),
.B2(n_105),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_166),
.A2(n_150),
.B1(n_136),
.B2(n_117),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_115),
.A2(n_95),
.B1(n_103),
.B2(n_92),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_135),
.B(n_10),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_173),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_135),
.B(n_10),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_172),
.B(n_179),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_113),
.B(n_98),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_177),
.A2(n_121),
.B1(n_117),
.B2(n_144),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_116),
.A2(n_103),
.B1(n_92),
.B2(n_79),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_149),
.B(n_147),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_125),
.A2(n_79),
.B1(n_107),
.B2(n_124),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_144),
.B1(n_162),
.B2(n_182),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_120),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_182),
.A2(n_138),
.B(n_145),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_133),
.B(n_122),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_183),
.B(n_132),
.Y(n_191)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_131),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_167),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_187),
.A2(n_208),
.B1(n_218),
.B2(n_207),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_190),
.A2(n_191),
.B(n_202),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_192),
.A2(n_195),
.B(n_215),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_176),
.B(n_111),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_193),
.B(n_194),
.Y(n_231)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

AOI32xp33_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_118),
.A3(n_141),
.B1(n_150),
.B2(n_110),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_110),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_196),
.B(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_185),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_198),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_117),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_205),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_130),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_200),
.B(n_212),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_201),
.Y(n_247)
);

OA21x2_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_121),
.B(n_130),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_185),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_204),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_220),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_153),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_184),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_211),
.A2(n_219),
.B1(n_206),
.B2(n_195),
.Y(n_243)
);

A2O1A1O1Ixp25_ASAP7_75t_L g212 ( 
.A1(n_183),
.A2(n_182),
.B(n_180),
.C(n_184),
.D(n_179),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_219),
.C(n_211),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_152),
.A2(n_159),
.B(n_153),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_L g217 ( 
.A1(n_177),
.A2(n_154),
.B1(n_164),
.B2(n_178),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_217),
.A2(n_223),
.B1(n_208),
.B2(n_187),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_206),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_170),
.A2(n_152),
.B1(n_163),
.B2(n_175),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_171),
.B(n_172),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_173),
.B(n_160),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_155),
.Y(n_233)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_164),
.A2(n_174),
.B1(n_169),
.B2(n_155),
.Y(n_223)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_227),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_212),
.B(n_169),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_229),
.B(n_237),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_233),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_190),
.A2(n_155),
.B(n_192),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_234),
.A2(n_235),
.B(n_236),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_191),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_213),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_239),
.Y(n_281)
);

INVx13_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_240),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_241),
.B(n_253),
.C(n_242),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_209),
.C(n_203),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_202),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_202),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_194),
.B(n_197),
.Y(n_244)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_244),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_255),
.B(n_202),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_188),
.B(n_216),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_246),
.B(n_188),
.Y(n_259)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

AOI322xp5_ASAP7_75t_L g253 ( 
.A1(n_187),
.A2(n_189),
.A3(n_221),
.B1(n_193),
.B2(n_216),
.C1(n_220),
.C2(n_204),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_198),
.B(n_189),
.Y(n_255)
);

OA22x2_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_243),
.B1(n_250),
.B2(n_245),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_230),
.Y(n_257)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_259),
.B(n_266),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_230),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_260),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_232),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_261),
.B(n_264),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_263),
.A2(n_270),
.B(n_255),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_232),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_268),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_210),
.Y(n_268)
);

OAI21xp33_ASAP7_75t_L g270 ( 
.A1(n_234),
.A2(n_210),
.B(n_236),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_224),
.B(n_241),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_258),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_233),
.Y(n_304)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_226),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_278),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_254),
.A2(n_245),
.B1(n_235),
.B2(n_256),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_282),
.B1(n_247),
.B2(n_248),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_225),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_272),
.C(n_229),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_254),
.A2(n_235),
.B1(n_247),
.B2(n_250),
.Y(n_282)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_292),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_290),
.A2(n_295),
.B1(n_266),
.B2(n_283),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_293),
.C(n_294),
.Y(n_309)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_224),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_277),
.A2(n_282),
.B1(n_274),
.B2(n_270),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_257),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_298),
.Y(n_318)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_268),
.B(n_246),
.C(n_239),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_305),
.C(n_279),
.Y(n_321)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_300),
.Y(n_325)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_301),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_302),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_269),
.B(n_255),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_303),
.Y(n_316)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_304),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_267),
.B(n_244),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_262),
.A2(n_252),
.B1(n_231),
.B2(n_228),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_306),
.Y(n_320)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_286),
.B(n_259),
.CI(n_228),
.CON(n_307),
.SN(n_307)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_307),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_311),
.A2(n_317),
.B1(n_324),
.B2(n_284),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_287),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_314),
.Y(n_326)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_285),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_315),
.A2(n_304),
.B(n_302),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_295),
.A2(n_271),
.B1(n_283),
.B2(n_281),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_291),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_280),
.C(n_281),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_323),
.C(n_286),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_288),
.B(n_280),
.C(n_265),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_290),
.A2(n_273),
.B1(n_275),
.B2(n_249),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_327),
.B(n_328),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_329),
.Y(n_350)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_320),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_330),
.B(n_331),
.Y(n_348)
);

NOR3xp33_ASAP7_75t_SL g331 ( 
.A(n_320),
.B(n_297),
.C(n_293),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_310),
.A2(n_315),
.B(n_312),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_332),
.A2(n_334),
.B(n_335),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_325),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_335),
.Y(n_342)
);

XNOR2x1_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_305),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_292),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_317),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_339),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_314),
.B(n_299),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_337),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_338),
.A2(n_312),
.B1(n_318),
.B2(n_308),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_309),
.B(n_294),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_342),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_326),
.B(n_319),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_343),
.A2(n_347),
.B(n_351),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_344),
.A2(n_324),
.B1(n_316),
.B2(n_325),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_332),
.A2(n_310),
.B(n_318),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_340),
.A2(n_308),
.B(n_313),
.Y(n_351)
);

A2O1A1Ixp33_ASAP7_75t_L g352 ( 
.A1(n_331),
.A2(n_316),
.B(n_323),
.C(n_311),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_352),
.A2(n_334),
.B(n_284),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_355),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_300),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_345),
.B(n_327),
.C(n_321),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_356),
.B(n_345),
.C(n_346),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_346),
.B(n_339),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_309),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_358),
.A2(n_352),
.B(n_347),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_348),
.A2(n_307),
.B1(n_251),
.B2(n_226),
.Y(n_360)
);

AOI322xp5_ASAP7_75t_L g366 ( 
.A1(n_360),
.A2(n_307),
.A3(n_350),
.B1(n_349),
.B2(n_344),
.C1(n_240),
.C2(n_328),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_238),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_361),
.B(n_362),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_351),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_365),
.Y(n_373)
);

INVxp33_ASAP7_75t_L g364 ( 
.A(n_353),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_364),
.B(n_369),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_366),
.A2(n_350),
.B1(n_359),
.B2(n_358),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_370),
.B(n_371),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_367),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_372),
.B(n_356),
.Y(n_375)
);

AOI31xp33_ASAP7_75t_L g376 ( 
.A1(n_375),
.A2(n_364),
.A3(n_357),
.B(n_373),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_376),
.A2(n_368),
.B(n_353),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_377),
.A2(n_374),
.B(n_238),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_378),
.Y(n_379)
);


endmodule