module fake_jpeg_9097_n_229 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_46),
.Y(n_67)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_45),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_34),
.B(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_60),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_32),
.B1(n_34),
.B2(n_17),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_70),
.B1(n_73),
.B2(n_17),
.Y(n_85)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_74),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_61),
.Y(n_79)
);

AO22x2_ASAP7_75t_L g66 ( 
.A1(n_37),
.A2(n_18),
.B1(n_30),
.B2(n_35),
.Y(n_66)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_66),
.A2(n_49),
.A3(n_27),
.B1(n_2),
.B2(n_3),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_68),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_29),
.B1(n_28),
.B2(n_26),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_32),
.B1(n_18),
.B2(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_76),
.Y(n_99)
);

CKINVDCx12_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_28),
.C(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_79),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_66),
.A2(n_47),
.B1(n_40),
.B2(n_20),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_80),
.A2(n_106),
.B1(n_87),
.B2(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_81),
.B(n_82),
.Y(n_125)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_95),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_93),
.B(n_84),
.C(n_88),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_40),
.B1(n_41),
.B2(n_36),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_86),
.A2(n_92),
.B1(n_107),
.B2(n_0),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_41),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_52),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_66),
.A2(n_20),
.B1(n_22),
.B2(n_24),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_57),
.A2(n_39),
.B1(n_38),
.B2(n_19),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_102),
.B1(n_0),
.B2(n_5),
.Y(n_126)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_19),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_63),
.B(n_38),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_49),
.C(n_59),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_24),
.B1(n_27),
.B2(n_2),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_104),
.Y(n_121)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_59),
.B(n_8),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_11),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_72),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_127),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_119),
.B1(n_105),
.B2(n_106),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_12),
.Y(n_154)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_114),
.B(n_115),
.Y(n_153)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_120),
.Y(n_132)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_123),
.B(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_59),
.Y(n_124)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_101),
.B1(n_6),
.B2(n_8),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_5),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_6),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_81),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_145),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_96),
.C(n_99),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_125),
.C(n_111),
.Y(n_165)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_142),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_141),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_143),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_86),
.B(n_95),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_148),
.B(n_152),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_5),
.B(n_104),
.Y(n_148)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_112),
.A2(n_101),
.B(n_14),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_154),
.B(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_158),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_166),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_117),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_162),
.B(n_145),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_119),
.Y(n_164)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_169),
.C(n_172),
.Y(n_182)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_168),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_114),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_150),
.B1(n_146),
.B2(n_142),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_131),
.C(n_115),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_113),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_165),
.C(n_169),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_147),
.B1(n_137),
.B2(n_140),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_178),
.A2(n_179),
.B1(n_156),
.B2(n_173),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_155),
.A2(n_145),
.B1(n_144),
.B2(n_140),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_168),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_186),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_154),
.B(n_136),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_183),
.A2(n_184),
.B(n_154),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_164),
.B(n_161),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_188),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

AOI322xp5_ASAP7_75t_SL g192 ( 
.A1(n_183),
.A2(n_172),
.A3(n_175),
.B1(n_180),
.B2(n_187),
.C1(n_136),
.C2(n_182),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_193),
.C(n_197),
.Y(n_206)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_157),
.Y(n_195)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_171),
.B1(n_162),
.B2(n_184),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_196),
.B(n_198),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_158),
.C(n_152),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_139),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_199),
.Y(n_208)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_200),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_198),
.B(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_201),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_179),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_203),
.B(n_190),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_208),
.A2(n_196),
.B(n_195),
.C(n_191),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_193),
.B1(n_197),
.B2(n_120),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_145),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_159),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_213),
.B(n_214),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_207),
.B(n_188),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_202),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_151),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_209),
.A3(n_204),
.B1(n_205),
.B2(n_206),
.C1(n_201),
.C2(n_202),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_14),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_218),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_15),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_215),
.C(n_118),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_222),
.A2(n_223),
.B(n_224),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_221),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_220),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_225),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_15),
.Y(n_229)
);


endmodule