module real_aes_7408_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_884;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_356;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_869;
wire n_613;
wire n_642;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_898;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_741;
wire n_314;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_0), .A2(n_243), .B1(n_369), .B2(n_374), .Y(n_769) );
XOR2x2_ASAP7_75t_L g502 ( .A(n_1), .B(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_2), .A2(n_172), .B1(n_351), .B2(n_355), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_3), .A2(n_54), .B1(n_337), .B2(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g611 ( .A(n_4), .Y(n_611) );
AOI222xp33_ASAP7_75t_L g522 ( .A1(n_5), .A2(n_25), .B1(n_233), .B2(n_523), .C1(n_524), .C2(n_526), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_6), .Y(n_748) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_7), .A2(n_170), .B1(n_381), .B2(n_385), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_8), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_9), .B(n_506), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_10), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_11), .A2(n_73), .B1(n_512), .B2(n_514), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_12), .A2(n_153), .B1(n_495), .B2(n_496), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_13), .A2(n_531), .B1(n_567), .B2(n_568), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_13), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_14), .A2(n_211), .B1(n_566), .B2(n_760), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_15), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g368 ( .A1(n_16), .A2(n_62), .B1(n_369), .B2(n_374), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g897 ( .A(n_17), .Y(n_897) );
XOR2x2_ASAP7_75t_L g423 ( .A(n_18), .B(n_424), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_19), .A2(n_205), .B1(n_350), .B2(n_354), .Y(n_349) );
INVx1_ASAP7_75t_L g417 ( .A(n_20), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_21), .A2(n_88), .B1(n_526), .B2(n_541), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_22), .A2(n_76), .B1(n_732), .B2(n_855), .Y(n_854) );
AO22x2_ASAP7_75t_L g311 ( .A1(n_23), .A2(n_82), .B1(n_312), .B2(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g833 ( .A(n_23), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g895 ( .A(n_24), .Y(n_895) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_26), .A2(n_287), .B(n_295), .C(n_835), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_27), .Y(n_630) );
AOI22xp33_ASAP7_75t_SL g719 ( .A1(n_28), .A2(n_196), .B1(n_520), .B2(n_564), .Y(n_719) );
INVx1_ASAP7_75t_L g812 ( .A(n_29), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_30), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_31), .A2(n_185), .B1(n_419), .B2(n_420), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_32), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_33), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_34), .A2(n_48), .B1(n_380), .B2(n_406), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_35), .A2(n_36), .B1(n_412), .B2(n_506), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_37), .A2(n_219), .B1(n_385), .B2(n_390), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_38), .A2(n_51), .B1(n_524), .B2(n_884), .Y(n_883) );
AO22x2_ASAP7_75t_L g315 ( .A1(n_39), .A2(n_85), .B1(n_312), .B2(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g834 ( .A(n_39), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_40), .A2(n_238), .B1(n_475), .B2(n_622), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_41), .A2(n_129), .B1(n_628), .B2(n_629), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g882 ( .A(n_42), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_43), .A2(n_210), .B1(n_406), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_SL g787 ( .A1(n_44), .A2(n_118), .B1(n_512), .B2(n_596), .Y(n_787) );
AOI22xp33_ASAP7_75t_SL g790 ( .A1(n_45), .A2(n_46), .B1(n_445), .B2(n_791), .Y(n_790) );
AOI22xp33_ASAP7_75t_SL g781 ( .A1(n_47), .A2(n_271), .B1(n_524), .B2(n_583), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_49), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_50), .B(n_412), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_52), .Y(n_664) );
AOI22xp5_ASAP7_75t_SL g400 ( .A1(n_53), .A2(n_267), .B1(n_401), .B2(n_403), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_55), .A2(n_242), .B1(n_456), .B2(n_457), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_56), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_57), .Y(n_464) );
AOI22xp33_ASAP7_75t_SL g788 ( .A1(n_58), .A2(n_245), .B1(n_374), .B2(n_598), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_59), .Y(n_665) );
XOR2x2_ASAP7_75t_L g776 ( .A(n_60), .B(n_777), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_61), .A2(n_262), .B1(n_524), .B2(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_63), .B(n_438), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_64), .A2(n_837), .B1(n_838), .B2(n_860), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_64), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_65), .A2(n_241), .B1(n_391), .B2(n_444), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_66), .A2(n_263), .B1(n_350), .B2(n_414), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_67), .A2(n_218), .B1(n_381), .B2(n_482), .Y(n_521) );
AOI22xp33_ASAP7_75t_SL g612 ( .A1(n_68), .A2(n_270), .B1(n_420), .B2(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_69), .B(n_617), .Y(n_616) );
CKINVDCx20_ASAP7_75t_R g888 ( .A(n_70), .Y(n_888) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_71), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_72), .B(n_337), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_74), .A2(n_186), .B1(n_408), .B2(n_732), .Y(n_731) );
AOI22xp33_ASAP7_75t_SL g683 ( .A1(n_75), .A2(n_148), .B1(n_354), .B2(n_430), .Y(n_683) );
AOI22xp33_ASAP7_75t_SL g707 ( .A1(n_77), .A2(n_123), .B1(n_496), .B2(n_708), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_78), .A2(n_154), .B1(n_553), .B2(n_603), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_79), .A2(n_95), .B1(n_564), .B2(n_566), .Y(n_563) );
AOI22xp33_ASAP7_75t_SL g359 ( .A1(n_80), .A2(n_113), .B1(n_360), .B2(n_365), .Y(n_359) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_81), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_83), .A2(n_142), .B1(n_375), .B2(n_482), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_84), .A2(n_171), .B1(n_355), .B2(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_86), .A2(n_222), .B1(n_370), .B2(n_518), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_87), .A2(n_217), .B1(n_391), .B2(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g293 ( .A(n_89), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_90), .B(n_435), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_91), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_92), .B(n_753), .Y(n_752) );
AOI22xp33_ASAP7_75t_SL g694 ( .A1(n_93), .A2(n_188), .B1(n_520), .B2(n_566), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_94), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g290 ( .A(n_96), .Y(n_290) );
INVx1_ASAP7_75t_L g421 ( .A(n_97), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_98), .A2(n_212), .B1(n_518), .B2(n_763), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_99), .A2(n_144), .B1(n_518), .B2(n_603), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_100), .A2(n_244), .B1(n_375), .B2(n_385), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_101), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_102), .A2(n_195), .B1(n_362), .B2(n_444), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_103), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g880 ( .A(n_104), .Y(n_880) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_105), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_106), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g842 ( .A(n_107), .Y(n_842) );
INVx1_ASAP7_75t_L g815 ( .A(n_108), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_109), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_110), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_111), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_112), .A2(n_206), .B1(n_561), .B2(n_562), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_114), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_115), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_116), .A2(n_128), .B1(n_475), .B2(n_596), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_117), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_119), .A2(n_163), .B1(n_420), .B2(n_508), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_120), .A2(n_125), .B1(n_495), .B2(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g808 ( .A(n_121), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_122), .A2(n_231), .B1(n_406), .B2(n_447), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_124), .A2(n_257), .B1(n_512), .B2(n_768), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_126), .A2(n_277), .B1(n_518), .B2(n_520), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_127), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_130), .A2(n_133), .B1(n_721), .B2(n_732), .Y(n_799) );
INVx1_ASAP7_75t_L g810 ( .A(n_131), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_132), .A2(n_204), .B1(n_375), .B2(n_482), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_134), .A2(n_174), .B1(n_457), .B2(n_598), .Y(n_733) );
AOI222xp33_ASAP7_75t_L g817 ( .A1(n_135), .A2(n_184), .B1(n_193), .B2(n_309), .C1(n_332), .C2(n_508), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_136), .A2(n_256), .B1(n_350), .B2(n_440), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_137), .A2(n_201), .B1(n_447), .B2(n_449), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_138), .A2(n_203), .B1(n_449), .B2(n_478), .Y(n_477) );
AOI22x1_ASAP7_75t_L g640 ( .A1(n_139), .A2(n_641), .B1(n_673), .B2(n_674), .Y(n_640) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_139), .Y(n_673) );
AOI222xp33_ASAP7_75t_L g742 ( .A1(n_140), .A2(n_175), .B1(n_221), .B2(n_309), .C1(n_548), .C2(n_613), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_141), .A2(n_279), .B1(n_710), .B2(n_711), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_143), .A2(n_261), .B1(n_449), .B2(n_721), .Y(n_720) );
AOI22xp33_ASAP7_75t_SL g387 ( .A1(n_145), .A2(n_187), .B1(n_388), .B2(n_391), .Y(n_387) );
INVx2_ASAP7_75t_L g294 ( .A(n_146), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_147), .A2(n_247), .B1(n_430), .B2(n_431), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g716 ( .A1(n_149), .A2(n_214), .B1(n_453), .B2(n_717), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_150), .Y(n_747) );
AOI222xp33_ASAP7_75t_L g497 ( .A1(n_151), .A2(n_165), .B1(n_225), .B2(n_309), .C1(n_419), .C2(n_498), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_152), .Y(n_549) );
AOI22xp33_ASAP7_75t_SL g597 ( .A1(n_155), .A2(n_168), .B1(n_598), .B2(n_599), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_156), .A2(n_230), .B1(n_452), .B2(n_453), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_157), .A2(n_250), .B1(n_354), .B2(n_541), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_158), .A2(n_278), .B1(n_401), .B2(n_599), .Y(n_892) );
AND2x6_ASAP7_75t_L g289 ( .A(n_159), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_159), .Y(n_827) );
AO22x2_ASAP7_75t_L g319 ( .A1(n_160), .A2(n_239), .B1(n_312), .B2(n_316), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_161), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_162), .A2(n_269), .B1(n_453), .B2(n_457), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_164), .Y(n_545) );
AOI22xp33_ASAP7_75t_SL g323 ( .A1(n_166), .A2(n_209), .B1(n_324), .B2(n_332), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_167), .A2(n_240), .B1(n_557), .B2(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g695 ( .A(n_169), .Y(n_695) );
AOI22xp33_ASAP7_75t_SL g379 ( .A1(n_173), .A2(n_282), .B1(n_380), .B2(n_383), .Y(n_379) );
XNOR2xp5_ASAP7_75t_L g696 ( .A(n_176), .B(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_SL g714 ( .A1(n_177), .A2(n_179), .B1(n_360), .B2(n_715), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_178), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_180), .A2(n_276), .B1(n_565), .B2(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g802 ( .A(n_181), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_182), .A2(n_572), .B1(n_573), .B2(n_604), .Y(n_571) );
CKINVDCx14_ASAP7_75t_R g604 ( .A(n_182), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_183), .A2(n_228), .B1(n_369), .B2(n_374), .Y(n_654) );
INVx1_ASAP7_75t_L g818 ( .A(n_189), .Y(n_818) );
AOI22xp33_ASAP7_75t_SL g691 ( .A1(n_190), .A2(n_234), .B1(n_512), .B2(n_624), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_191), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_192), .B(n_506), .Y(n_686) );
AO22x2_ASAP7_75t_L g321 ( .A1(n_194), .A2(n_249), .B1(n_312), .B2(n_313), .Y(n_321) );
AOI22xp33_ASAP7_75t_SL g621 ( .A1(n_197), .A2(n_254), .B1(n_565), .B2(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_198), .B(n_337), .Y(n_783) );
XOR2x2_ASAP7_75t_L g728 ( .A(n_199), .B(n_729), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g652 ( .A(n_200), .Y(n_652) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_202), .A2(n_208), .B1(n_482), .B2(n_624), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_207), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_213), .A2(n_258), .B1(n_496), .B2(n_541), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g849 ( .A(n_215), .Y(n_849) );
INVx1_ASAP7_75t_L g851 ( .A(n_216), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_220), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_223), .A2(n_744), .B1(n_770), .B2(n_771), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_223), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_224), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_226), .A2(n_280), .B1(n_351), .B2(n_613), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_227), .B(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_SL g792 ( .A1(n_229), .A2(n_273), .B1(n_765), .B2(n_793), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_232), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g899 ( .A(n_235), .Y(n_899) );
CKINVDCx20_ASAP7_75t_R g879 ( .A(n_236), .Y(n_879) );
XOR2x2_ASAP7_75t_L g302 ( .A(n_237), .B(n_303), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_239), .B(n_832), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_246), .A2(n_252), .B1(n_452), .B2(n_741), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_248), .Y(n_466) );
INVx1_ASAP7_75t_L g830 ( .A(n_249), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_251), .A2(n_281), .B1(n_337), .B2(n_710), .Y(n_735) );
INVx1_ASAP7_75t_L g322 ( .A(n_253), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_255), .Y(n_645) );
CKINVDCx16_ASAP7_75t_R g870 ( .A(n_259), .Y(n_870) );
OA22x2_ASAP7_75t_L g872 ( .A1(n_259), .A2(n_870), .B1(n_873), .B2(n_874), .Y(n_872) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_260), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_264), .A2(n_266), .B1(n_364), .B2(n_603), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_265), .Y(n_780) );
INVx1_ASAP7_75t_L g312 ( .A(n_268), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_268), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_272), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_274), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_275), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g844 ( .A(n_283), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_284), .B(n_436), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_285), .A2(n_461), .B1(n_499), .B2(n_500), .Y(n_460) );
CKINVDCx16_ASAP7_75t_R g499 ( .A(n_285), .Y(n_499) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_290), .Y(n_826) );
OAI21xp5_ASAP7_75t_L g868 ( .A1(n_291), .A2(n_825), .B(n_869), .Y(n_868) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_292), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_725), .B1(n_820), .B2(n_821), .C(n_822), .Y(n_295) );
INVx1_ASAP7_75t_L g820 ( .A(n_296), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B1(n_638), .B2(n_639), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_458), .B1(n_636), .B2(n_637), .Y(n_298) );
INVxp67_ASAP7_75t_SL g636 ( .A(n_299), .Y(n_636) );
XOR2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_394), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND3x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_358), .C(n_378), .Y(n_303) );
NOR2x1_ASAP7_75t_SL g304 ( .A(n_305), .B(n_335), .Y(n_304) );
OAI21xp5_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_322), .B(n_323), .Y(n_305) );
OAI222xp33_ASAP7_75t_L g543 ( .A1(n_306), .A2(n_544), .B1(n_545), .B2(n_546), .C1(n_547), .C2(n_549), .Y(n_543) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx2_ASAP7_75t_L g416 ( .A(n_308), .Y(n_416) );
INVx4_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_SL g427 ( .A(n_309), .Y(n_427) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_309), .Y(n_523) );
BUFx3_ASAP7_75t_L g610 ( .A(n_309), .Y(n_610) );
INVx2_ASAP7_75t_L g681 ( .A(n_309), .Y(n_681) );
AND2x6_ASAP7_75t_L g309 ( .A(n_310), .B(n_317), .Y(n_309) );
AND2x4_ASAP7_75t_L g355 ( .A(n_310), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g591 ( .A(n_310), .Y(n_591) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_315), .Y(n_310) );
AND2x2_ASAP7_75t_L g331 ( .A(n_311), .B(n_319), .Y(n_331) );
INVx2_ASAP7_75t_L g341 ( .A(n_311), .Y(n_341) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g316 ( .A(n_314), .Y(n_316) );
INVx2_ASAP7_75t_L g330 ( .A(n_315), .Y(n_330) );
AND2x2_ASAP7_75t_L g340 ( .A(n_315), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g348 ( .A(n_315), .B(n_341), .Y(n_348) );
INVx1_ASAP7_75t_L g353 ( .A(n_315), .Y(n_353) );
AND2x6_ASAP7_75t_L g364 ( .A(n_317), .B(n_347), .Y(n_364) );
AND2x2_ASAP7_75t_L g382 ( .A(n_317), .B(n_367), .Y(n_382) );
AND2x4_ASAP7_75t_L g390 ( .A(n_317), .B(n_340), .Y(n_390) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
AND2x2_ASAP7_75t_L g342 ( .A(n_318), .B(n_321), .Y(n_342) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g373 ( .A(n_319), .B(n_357), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_319), .B(n_321), .Y(n_377) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g329 ( .A(n_321), .Y(n_329) );
INVx1_ASAP7_75t_L g357 ( .A(n_321), .Y(n_357) );
INVx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx4_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g702 ( .A(n_326), .Y(n_702) );
BUFx2_ASAP7_75t_L g884 ( .A(n_326), .Y(n_884) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx2_ASAP7_75t_L g419 ( .A(n_327), .Y(n_419) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_327), .Y(n_440) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_327), .Y(n_508) );
BUFx4f_ASAP7_75t_SL g613 ( .A(n_327), .Y(n_613) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_331), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g334 ( .A(n_329), .Y(n_334) );
AND2x2_ASAP7_75t_L g367 ( .A(n_330), .B(n_341), .Y(n_367) );
INVx1_ASAP7_75t_L g588 ( .A(n_330), .Y(n_588) );
AND2x4_ASAP7_75t_L g333 ( .A(n_331), .B(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g351 ( .A(n_331), .B(n_352), .Y(n_351) );
NAND2x1p5_ASAP7_75t_L g587 ( .A(n_331), .B(n_588), .Y(n_587) );
BUFx4f_ASAP7_75t_L g753 ( .A(n_332), .Y(n_753) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx12f_ASAP7_75t_L g420 ( .A(n_333), .Y(n_420) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_333), .Y(n_430) );
INVx1_ASAP7_75t_L g704 ( .A(n_333), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_343), .C(n_349), .Y(n_335) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g711 ( .A(n_338), .Y(n_711) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
BUFx2_ASAP7_75t_L g438 ( .A(n_339), .Y(n_438) );
BUFx4f_ASAP7_75t_L g506 ( .A(n_339), .Y(n_506) );
AND2x6_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
AND2x2_ASAP7_75t_L g372 ( .A(n_340), .B(n_373), .Y(n_372) );
NAND2x1p5_ASAP7_75t_L g492 ( .A(n_340), .B(n_342), .Y(n_492) );
AND2x4_ASAP7_75t_L g346 ( .A(n_342), .B(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g366 ( .A(n_342), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g487 ( .A(n_342), .Y(n_487) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g412 ( .A(n_345), .Y(n_412) );
INVx5_ASAP7_75t_L g436 ( .A(n_345), .Y(n_436) );
INVx2_ASAP7_75t_L g617 ( .A(n_345), .Y(n_617) );
INVx4_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g486 ( .A(n_348), .B(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx3_ASAP7_75t_L g495 ( .A(n_351), .Y(n_495) );
INVx1_ASAP7_75t_L g542 ( .A(n_351), .Y(n_542) );
BUFx2_ASAP7_75t_L g708 ( .A(n_351), .Y(n_708) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x6_ASAP7_75t_L g376 ( .A(n_353), .B(n_377), .Y(n_376) );
BUFx2_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_355), .Y(n_414) );
BUFx3_ASAP7_75t_L g496 ( .A(n_355), .Y(n_496) );
BUFx2_ASAP7_75t_SL g526 ( .A(n_355), .Y(n_526) );
INVx1_ASAP7_75t_L g592 ( .A(n_356), .Y(n_592) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_368), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g406 ( .A(n_363), .Y(n_406) );
INVx5_ASAP7_75t_SL g480 ( .A(n_363), .Y(n_480) );
INVx4_ASAP7_75t_L g553 ( .A(n_363), .Y(n_553) );
INVx1_ASAP7_75t_L g741 ( .A(n_363), .Y(n_741) );
INVx11_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx11_ASAP7_75t_L g519 ( .A(n_364), .Y(n_519) );
INVx4_ASAP7_75t_L g409 ( .A(n_365), .Y(n_409) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx3_ASAP7_75t_L g456 ( .A(n_366), .Y(n_456) );
BUFx3_ASAP7_75t_L g475 ( .A(n_366), .Y(n_475) );
INVx2_ASAP7_75t_L g513 ( .A(n_366), .Y(n_513) );
BUFx3_ASAP7_75t_L g629 ( .A(n_366), .Y(n_629) );
AND2x2_ASAP7_75t_L g386 ( .A(n_367), .B(n_373), .Y(n_386) );
AND2x4_ASAP7_75t_L g392 ( .A(n_367), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_367), .B(n_373), .Y(n_469) );
BUFx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_370), .Y(n_598) );
INVx5_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx4_ASAP7_75t_L g402 ( .A(n_371), .Y(n_402) );
BUFx3_ASAP7_75t_L g454 ( .A(n_371), .Y(n_454) );
INVx2_ASAP7_75t_L g482 ( .A(n_371), .Y(n_482) );
INVx3_ASAP7_75t_L g557 ( .A(n_371), .Y(n_557) );
INVx8_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g403 ( .A(n_375), .Y(n_403) );
BUFx2_ASAP7_75t_L g457 ( .A(n_375), .Y(n_457) );
BUFx2_ASAP7_75t_L g599 ( .A(n_375), .Y(n_599) );
INVx6_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g558 ( .A(n_376), .Y(n_558) );
INVx1_ASAP7_75t_SL g717 ( .A(n_376), .Y(n_717) );
INVx1_ASAP7_75t_L g393 ( .A(n_377), .Y(n_393) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_387), .Y(n_378) );
INVx1_ASAP7_75t_SL g472 ( .A(n_380), .Y(n_472) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx3_ASAP7_75t_L g561 ( .A(n_381), .Y(n_561) );
INVx3_ASAP7_75t_L g644 ( .A(n_381), .Y(n_644) );
BUFx3_ASAP7_75t_L g768 ( .A(n_381), .Y(n_768) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g448 ( .A(n_382), .Y(n_448) );
BUFx2_ASAP7_75t_SL g596 ( .A(n_382), .Y(n_596) );
BUFx2_ASAP7_75t_SL g732 ( .A(n_382), .Y(n_732) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx3_ASAP7_75t_L g445 ( .A(n_386), .Y(n_445) );
BUFx3_ASAP7_75t_L g565 ( .A(n_386), .Y(n_565) );
BUFx3_ASAP7_75t_L g855 ( .A(n_386), .Y(n_855) );
INVx2_ASAP7_75t_L g465 ( .A(n_388), .Y(n_465) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g452 ( .A(n_389), .Y(n_452) );
INVx2_ASAP7_75t_L g562 ( .A(n_389), .Y(n_562) );
INVx3_ASAP7_75t_L g603 ( .A(n_389), .Y(n_603) );
INVx6_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx3_ASAP7_75t_L g520 ( .A(n_390), .Y(n_520) );
BUFx3_ASAP7_75t_L g765 ( .A(n_390), .Y(n_765) );
BUFx2_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
BUFx3_ASAP7_75t_L g449 ( .A(n_392), .Y(n_449) );
INVx1_ASAP7_75t_L g515 ( .A(n_392), .Y(n_515) );
BUFx3_ASAP7_75t_L g566 ( .A(n_392), .Y(n_566) );
BUFx2_ASAP7_75t_L g622 ( .A(n_392), .Y(n_622) );
BUFx3_ASAP7_75t_L g739 ( .A(n_392), .Y(n_739) );
BUFx2_ASAP7_75t_SL g791 ( .A(n_392), .Y(n_791) );
AND2x2_ASAP7_75t_L g624 ( .A(n_393), .B(n_588), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_422), .B2(n_423), .Y(n_394) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
XOR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_421), .Y(n_396) );
NOR4xp75_ASAP7_75t_L g397 ( .A(n_398), .B(n_404), .C(n_410), .D(n_415), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_399), .B(n_400), .Y(n_398) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2x1_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
INVx4_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI221xp5_ASAP7_75t_SL g551 ( .A1(n_409), .A2(n_552), .B1(n_554), .B2(n_555), .C(n_556), .Y(n_551) );
INVx3_ASAP7_75t_L g721 ( .A(n_409), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_411), .B(n_413), .Y(n_410) );
INVx1_ASAP7_75t_SL g432 ( .A(n_414), .Y(n_432) );
OAI21xp5_ASAP7_75t_SL g415 ( .A1(n_416), .A2(n_417), .B(n_418), .Y(n_415) );
OAI21xp5_ASAP7_75t_SL g580 ( .A1(n_416), .A2(n_581), .B(n_582), .Y(n_580) );
INVx2_ASAP7_75t_L g525 ( .A(n_420), .Y(n_525) );
BUFx4f_ASAP7_75t_SL g548 ( .A(n_420), .Y(n_548) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_425), .B(n_441), .Y(n_424) );
NOR2xp33_ASAP7_75t_SL g425 ( .A(n_426), .B(n_433), .Y(n_425) );
OAI21xp5_ASAP7_75t_SL g426 ( .A1(n_427), .A2(n_428), .B(n_429), .Y(n_426) );
BUFx2_ASAP7_75t_L g498 ( .A(n_430), .Y(n_498) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_437), .C(n_439), .Y(n_433) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_436), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_440), .Y(n_544) );
NOR2x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_450), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_446), .Y(n_442) );
BUFx4f_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g628 ( .A(n_448), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_455), .Y(n_450) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_456), .Y(n_647) );
INVx1_ASAP7_75t_L g898 ( .A(n_456), .Y(n_898) );
INVx1_ASAP7_75t_SL g637 ( .A(n_458), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_529), .B1(n_634), .B2(n_635), .Y(n_458) );
INVx1_ASAP7_75t_L g635 ( .A(n_459), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_501), .B1(n_527), .B2(n_528), .Y(n_459) );
INVx1_ASAP7_75t_L g527 ( .A(n_460), .Y(n_527) );
INVx2_ASAP7_75t_SL g500 ( .A(n_461), .Y(n_500) );
AND4x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_476), .C(n_483), .D(n_497), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_470), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_466), .B2(n_467), .Y(n_463) );
OAI221xp5_ASAP7_75t_SL g651 ( .A1(n_465), .A2(n_467), .B1(n_652), .B2(n_653), .C(n_654), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_465), .A2(n_467), .B1(n_894), .B2(n_895), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_467), .A2(n_808), .B1(n_809), .B2(n_810), .Y(n_807) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B1(n_473), .B2(n_474), .Y(n_470) );
INVxp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_481), .Y(n_476) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OAI221xp5_ASAP7_75t_SL g484 ( .A1(n_485), .A2(n_488), .B1(n_489), .B2(n_493), .C(n_494), .Y(n_484) );
INVx1_ASAP7_75t_L g878 ( .A(n_485), .Y(n_878) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g535 ( .A(n_486), .Y(n_535) );
BUFx3_ASAP7_75t_L g843 ( .A(n_486), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_489), .A2(n_534), .B1(n_747), .B2(n_748), .Y(n_746) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx3_ASAP7_75t_L g579 ( .A(n_491), .Y(n_579) );
BUFx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g538 ( .A(n_492), .Y(n_538) );
INVxp67_ASAP7_75t_L g528 ( .A(n_501), .Y(n_528) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND4xp75_ASAP7_75t_L g503 ( .A(n_504), .B(n_509), .C(n_516), .D(n_522), .Y(n_503) );
AND2x2_ASAP7_75t_SL g504 ( .A(n_505), .B(n_507), .Y(n_504) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_508), .Y(n_583) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_515), .A2(n_897), .B1(n_898), .B2(n_899), .Y(n_896) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_521), .Y(n_516) );
INVx4_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_SL g793 ( .A(n_519), .Y(n_793) );
INVx3_ASAP7_75t_L g814 ( .A(n_519), .Y(n_814) );
INVx2_ASAP7_75t_L g663 ( .A(n_523), .Y(n_663) );
INVx2_ASAP7_75t_SL g700 ( .A(n_523), .Y(n_700) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g634 ( .A(n_529), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_569), .B1(n_570), .B2(n_633), .Y(n_529) );
INVx1_ASAP7_75t_SL g633 ( .A(n_530), .Y(n_633) );
INVx1_ASAP7_75t_L g568 ( .A(n_531), .Y(n_568) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_550), .Y(n_531) );
NOR2xp33_ASAP7_75t_SL g532 ( .A(n_533), .B(n_543), .Y(n_532) );
OAI221xp5_ASAP7_75t_SL g533 ( .A1(n_534), .A2(n_536), .B1(n_537), .B2(n_539), .C(n_540), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_534), .A2(n_657), .B1(n_658), .B2(n_659), .Y(n_656) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g577 ( .A(n_535), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_537), .A2(n_842), .B1(n_843), .B2(n_844), .Y(n_841) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g659 ( .A(n_538), .Y(n_659) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OAI222xp33_ASAP7_75t_L g660 ( .A1(n_547), .A2(n_661), .B1(n_662), .B2(n_663), .C1(n_664), .C2(n_665), .Y(n_660) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_559), .Y(n_550) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
NAND2xp33_ASAP7_75t_SL g559 ( .A(n_560), .B(n_563), .Y(n_559) );
BUFx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g761 ( .A(n_565), .Y(n_761) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_566), .Y(n_650) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
AO22x1_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_605), .B1(n_631), .B2(n_632), .Y(n_570) );
INVx1_ASAP7_75t_L g632 ( .A(n_571), .Y(n_632) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_593), .Y(n_573) );
NOR3xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_580), .C(n_584), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B1(n_578), .B2(n_579), .Y(n_575) );
OA211x2_ASAP7_75t_L g801 ( .A1(n_579), .A2(n_802), .B(n_803), .C(n_805), .Y(n_801) );
OAI22xp5_ASAP7_75t_SL g876 ( .A1(n_579), .A2(n_877), .B1(n_879), .B2(n_880), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_586), .B1(n_589), .B2(n_590), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_586), .A2(n_671), .B1(n_755), .B2(n_756), .Y(n_754) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx4_ASAP7_75t_L g669 ( .A(n_587), .Y(n_669) );
BUFx3_ASAP7_75t_L g850 ( .A(n_587), .Y(n_850) );
OAI22xp33_ASAP7_75t_SL g885 ( .A1(n_587), .A2(n_886), .B1(n_887), .B2(n_888), .Y(n_885) );
CKINVDCx16_ASAP7_75t_R g672 ( .A(n_590), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_590), .A2(n_849), .B1(n_850), .B2(n_851), .Y(n_848) );
OR2x6_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_600), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g816 ( .A(n_603), .Y(n_816) );
INVx3_ASAP7_75t_SL g631 ( .A(n_605), .Y(n_631) );
XOR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_630), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_607), .B(n_619), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_614), .Y(n_607) );
OAI21xp5_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_611), .B(n_612), .Y(n_608) );
OAI21xp33_ASAP7_75t_L g845 ( .A1(n_609), .A2(n_846), .B(n_847), .Y(n_845) );
OAI21xp33_ASAP7_75t_SL g881 ( .A1(n_609), .A2(n_882), .B(n_883), .Y(n_881) );
INVx3_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g661 ( .A(n_613), .Y(n_661) );
NAND3xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .C(n_618), .Y(n_614) );
BUFx2_ASAP7_75t_L g804 ( .A(n_617), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_625), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_675), .B1(n_723), .B2(n_724), .Y(n_639) );
INVx1_ASAP7_75t_L g723 ( .A(n_640), .Y(n_723) );
INVx1_ASAP7_75t_L g674 ( .A(n_641), .Y(n_674) );
AND2x2_ASAP7_75t_SL g641 ( .A(n_642), .B(n_655), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_651), .Y(n_642) );
OAI221xp5_ASAP7_75t_SL g643 ( .A1(n_644), .A2(n_645), .B1(n_646), .B2(n_648), .C(n_649), .Y(n_643) );
INVx2_ASAP7_75t_L g715 ( .A(n_644), .Y(n_715) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NOR3xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_660), .C(n_666), .Y(n_655) );
OAI221xp5_ASAP7_75t_L g749 ( .A1(n_661), .A2(n_700), .B1(n_750), .B2(n_751), .C(n_752), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_670), .B2(n_671), .Y(n_666) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g887 ( .A(n_672), .Y(n_887) );
INVx2_ASAP7_75t_L g724 ( .A(n_675), .Y(n_724) );
OA22x2_ASAP7_75t_SL g675 ( .A1(n_676), .A2(n_677), .B1(n_696), .B2(n_722), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
XOR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_695), .Y(n_677) );
NAND2x1_ASAP7_75t_L g678 ( .A(n_679), .B(n_688), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_684), .Y(n_679) );
OAI21xp5_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_682), .B(n_683), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .C(n_687), .Y(n_684) );
NOR2x1_ASAP7_75t_L g688 ( .A(n_689), .B(n_692), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g722 ( .A(n_696), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_712), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_706), .Y(n_698) );
OAI222xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_702), .B2(n_703), .C1(n_704), .C2(n_705), .Y(n_699) );
OAI21xp5_ASAP7_75t_SL g779 ( .A1(n_700), .A2(n_780), .B(n_781), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_718), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
INVx1_ASAP7_75t_L g821 ( .A(n_725), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B1(n_774), .B2(n_775), .Y(n_725) );
INVx3_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OA22x2_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_743), .B1(n_772), .B2(n_773), .Y(n_727) );
INVx1_ASAP7_75t_L g773 ( .A(n_728), .Y(n_773) );
NAND4xp75_ASAP7_75t_L g729 ( .A(n_730), .B(n_734), .C(n_737), .D(n_742), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .Y(n_730) );
AND2x2_ASAP7_75t_SL g734 ( .A(n_735), .B(n_736), .Y(n_734) );
AND2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_740), .Y(n_737) );
INVxp67_ASAP7_75t_L g809 ( .A(n_739), .Y(n_809) );
INVx1_ASAP7_75t_L g772 ( .A(n_743), .Y(n_772) );
INVx2_ASAP7_75t_L g771 ( .A(n_744), .Y(n_771) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_757), .Y(n_744) );
NOR3xp33_ASAP7_75t_L g745 ( .A(n_746), .B(n_749), .C(n_754), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_766), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_762), .Y(n_758) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx3_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_769), .Y(n_766) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
OAI22xp5_ASAP7_75t_SL g775 ( .A1(n_776), .A2(n_794), .B1(n_795), .B2(n_819), .Y(n_775) );
INVx1_ASAP7_75t_L g819 ( .A(n_776), .Y(n_819) );
NAND3xp33_ASAP7_75t_L g777 ( .A(n_778), .B(n_786), .C(n_789), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_782), .Y(n_778) );
NAND3xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .C(n_785), .Y(n_782) );
AND2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
AND2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_792), .Y(n_789) );
INVx1_ASAP7_75t_SL g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
XOR2x2_ASAP7_75t_L g796 ( .A(n_797), .B(n_818), .Y(n_796) );
NAND4xp75_ASAP7_75t_L g797 ( .A(n_798), .B(n_801), .C(n_806), .D(n_817), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_811), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_813), .B1(n_815), .B2(n_816), .Y(n_811) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_SL g822 ( .A(n_823), .Y(n_822) );
NOR2x1_ASAP7_75t_L g823 ( .A(n_824), .B(n_828), .Y(n_823) );
OR2x2_ASAP7_75t_SL g902 ( .A(n_824), .B(n_829), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_825), .B(n_827), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_825), .Y(n_862) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_826), .B(n_866), .Y(n_869) );
CKINVDCx16_ASAP7_75t_R g866 ( .A(n_827), .Y(n_866) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_829), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
OAI322xp33_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_861), .A3(n_863), .B1(n_867), .B2(n_870), .C1(n_871), .C2(n_900), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_838), .Y(n_837) );
HB1xp67_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_840), .B(n_852), .Y(n_839) );
NOR3xp33_ASAP7_75t_L g840 ( .A(n_841), .B(n_845), .C(n_848), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_853), .B(n_857), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_854), .B(n_856), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_858), .B(n_859), .Y(n_857) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
HB1xp67_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_868), .Y(n_867) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_889), .Y(n_874) );
NOR3xp33_ASAP7_75t_L g875 ( .A(n_876), .B(n_881), .C(n_885), .Y(n_875) );
INVx2_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
NOR3xp33_ASAP7_75t_L g889 ( .A(n_890), .B(n_893), .C(n_896), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_891), .B(n_892), .Y(n_890) );
CKINVDCx20_ASAP7_75t_R g900 ( .A(n_901), .Y(n_900) );
CKINVDCx20_ASAP7_75t_R g901 ( .A(n_902), .Y(n_901) );
endmodule