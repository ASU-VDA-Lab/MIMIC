module fake_aes_2891_n_24 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_24);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_24;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
wire n_21;
INVx3_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
BUFx3_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_11), .Y(n_17) );
O2A1O1Ixp33_ASAP7_75t_SL g18 ( .A1(n_15), .A2(n_0), .B(n_2), .C(n_3), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
AOI21xp33_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_12), .B(n_14), .Y(n_21) );
NAND2xp5_ASAP7_75t_SL g22 ( .A(n_21), .B(n_16), .Y(n_22) );
AO21x2_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_18), .B(n_13), .Y(n_23) );
AOI21xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_8), .B(n_9), .Y(n_24) );
endmodule