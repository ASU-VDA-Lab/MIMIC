module fake_netlist_1_7275_n_707 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_707);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_707;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g81 ( .A(n_41), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_23), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_54), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_61), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_58), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_22), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_14), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_28), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_8), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_62), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_34), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_49), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_78), .Y(n_93) );
INVx1_ASAP7_75t_SL g94 ( .A(n_2), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_6), .Y(n_95) );
CKINVDCx14_ASAP7_75t_R g96 ( .A(n_56), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_4), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_52), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_75), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_39), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_20), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_1), .Y(n_102) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_71), .Y(n_103) );
NOR2xp67_ASAP7_75t_L g104 ( .A(n_50), .B(n_48), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_17), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_10), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_64), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_26), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_46), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_31), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_18), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_36), .Y(n_112) );
INVxp33_ASAP7_75t_SL g113 ( .A(n_4), .Y(n_113) );
NOR2xp67_ASAP7_75t_L g114 ( .A(n_63), .B(n_1), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_79), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_76), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_59), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_27), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_19), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_67), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_29), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_35), .Y(n_122) );
NOR2xp67_ASAP7_75t_L g123 ( .A(n_15), .B(n_17), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_42), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_53), .Y(n_125) );
INVxp67_ASAP7_75t_L g126 ( .A(n_33), .Y(n_126) );
INVx1_ASAP7_75t_SL g127 ( .A(n_8), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_25), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_70), .Y(n_129) );
INVx1_ASAP7_75t_SL g130 ( .A(n_82), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_82), .Y(n_131) );
NAND2x1p5_ASAP7_75t_L g132 ( .A(n_111), .B(n_32), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_103), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_92), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_91), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_92), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_105), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_103), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_87), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_91), .Y(n_140) );
NOR2xp67_ASAP7_75t_L g141 ( .A(n_124), .B(n_0), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_105), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_107), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_107), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_93), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_96), .B(n_0), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_83), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_117), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_117), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_89), .B(n_2), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_81), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_111), .B(n_3), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_103), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_95), .B(n_3), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_101), .B(n_5), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_106), .B(n_5), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_81), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_103), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_103), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_84), .B(n_6), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_93), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_85), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_86), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_98), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_88), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_98), .Y(n_166) );
OAI21x1_ASAP7_75t_L g167 ( .A1(n_90), .A2(n_40), .B(n_77), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_99), .B(n_7), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_100), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_113), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_108), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_109), .Y(n_172) );
AND2x6_ASAP7_75t_L g173 ( .A(n_110), .B(n_38), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_115), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_119), .B(n_7), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_162), .Y(n_176) );
AND3x4_ASAP7_75t_L g177 ( .A(n_141), .B(n_123), .C(n_114), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_162), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_162), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_162), .Y(n_180) );
INVx1_ASAP7_75t_SL g181 ( .A(n_130), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_162), .Y(n_182) );
OAI22xp33_ASAP7_75t_L g183 ( .A1(n_170), .A2(n_113), .B1(n_97), .B2(n_102), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_162), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_146), .B(n_94), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_171), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_143), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_152), .A2(n_127), .B1(n_120), .B2(n_129), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_171), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_146), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_147), .B(n_128), .Y(n_191) );
AND2x6_ASAP7_75t_L g192 ( .A(n_152), .B(n_118), .Y(n_192) );
INVx2_ASAP7_75t_SL g193 ( .A(n_163), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_147), .B(n_126), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_151), .A2(n_87), .B1(n_97), .B2(n_102), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_157), .B(n_125), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_171), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_135), .B(n_112), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_144), .B(n_122), .Y(n_199) );
AND2x6_ASAP7_75t_L g200 ( .A(n_135), .B(n_116), .Y(n_200) );
NOR2x1p5_ASAP7_75t_L g201 ( .A(n_131), .B(n_9), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_140), .B(n_121), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_169), .B(n_104), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_171), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_171), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_148), .B(n_43), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_140), .B(n_9), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_169), .B(n_10), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_171), .Y(n_209) );
INVx1_ASAP7_75t_SL g210 ( .A(n_149), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_133), .Y(n_211) );
BUFx2_ASAP7_75t_L g212 ( .A(n_164), .Y(n_212) );
INVx3_ASAP7_75t_L g213 ( .A(n_145), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_134), .Y(n_214) );
BUFx3_ASAP7_75t_L g215 ( .A(n_173), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_136), .Y(n_216) );
INVx6_ASAP7_75t_L g217 ( .A(n_173), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_166), .B(n_45), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_133), .Y(n_219) );
INVx4_ASAP7_75t_SL g220 ( .A(n_173), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_133), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_161), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_159), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_161), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_161), .Y(n_225) );
INVx5_ASAP7_75t_L g226 ( .A(n_173), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_138), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_145), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_159), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_172), .B(n_44), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_172), .B(n_11), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_138), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_145), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_159), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_138), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_145), .Y(n_236) );
NOR3xp33_ASAP7_75t_SL g237 ( .A(n_183), .B(n_175), .C(n_150), .Y(n_237) );
AND2x2_ASAP7_75t_SL g238 ( .A(n_207), .B(n_208), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_222), .Y(n_239) );
NAND2xp33_ASAP7_75t_SL g240 ( .A(n_207), .B(n_174), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_207), .A2(n_173), .B1(n_174), .B2(n_165), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_213), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_215), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_208), .Y(n_244) );
INVx4_ASAP7_75t_L g245 ( .A(n_226), .Y(n_245) );
NOR3xp33_ASAP7_75t_SL g246 ( .A(n_214), .B(n_154), .C(n_156), .Y(n_246) );
BUFx3_ASAP7_75t_L g247 ( .A(n_215), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_176), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_226), .Y(n_249) );
NOR3xp33_ASAP7_75t_SL g250 ( .A(n_214), .B(n_155), .C(n_160), .Y(n_250) );
CKINVDCx8_ASAP7_75t_R g251 ( .A(n_216), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_222), .Y(n_252) );
INVx2_ASAP7_75t_SL g253 ( .A(n_192), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_224), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_193), .A2(n_167), .B(n_173), .Y(n_255) );
BUFx3_ASAP7_75t_L g256 ( .A(n_217), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_176), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_202), .B(n_165), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_182), .Y(n_259) );
BUFx10_ASAP7_75t_L g260 ( .A(n_192), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_208), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_182), .Y(n_262) );
NAND2x1_ASAP7_75t_L g263 ( .A(n_200), .B(n_173), .Y(n_263) );
NAND3xp33_ASAP7_75t_SL g264 ( .A(n_181), .B(n_139), .C(n_132), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_213), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_202), .B(n_165), .Y(n_266) );
CKINVDCx11_ASAP7_75t_R g267 ( .A(n_210), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_186), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_192), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_192), .A2(n_173), .B1(n_163), .B2(n_165), .Y(n_270) );
INVx3_ASAP7_75t_L g271 ( .A(n_213), .Y(n_271) );
NOR3xp33_ASAP7_75t_SL g272 ( .A(n_216), .B(n_168), .C(n_142), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_186), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_198), .B(n_191), .Y(n_274) );
NAND3xp33_ASAP7_75t_SL g275 ( .A(n_187), .B(n_132), .C(n_142), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_198), .B(n_163), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_193), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_190), .B(n_163), .Y(n_278) );
INVx3_ASAP7_75t_L g279 ( .A(n_224), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_197), .Y(n_280) );
INVx1_ASAP7_75t_SL g281 ( .A(n_212), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_192), .A2(n_141), .B1(n_132), .B2(n_137), .Y(n_282) );
NOR2xp33_ASAP7_75t_R g283 ( .A(n_187), .B(n_137), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_217), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_226), .Y(n_285) );
OR2x6_ASAP7_75t_L g286 ( .A(n_201), .B(n_167), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_197), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_228), .Y(n_288) );
OAI22xp33_ASAP7_75t_L g289 ( .A1(n_195), .A2(n_137), .B1(n_158), .B2(n_153), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_212), .B(n_137), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_204), .Y(n_291) );
NAND3xp33_ASAP7_75t_SL g292 ( .A(n_177), .B(n_153), .C(n_158), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_226), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_228), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_226), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_233), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_233), .Y(n_297) );
NOR3xp33_ASAP7_75t_SL g298 ( .A(n_199), .B(n_11), .C(n_12), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_236), .Y(n_299) );
NAND2xp33_ASAP7_75t_SL g300 ( .A(n_201), .B(n_159), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_185), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_236), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_196), .B(n_55), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_185), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_253), .B(n_276), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_279), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_253), .B(n_190), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_276), .B(n_192), .Y(n_308) );
OAI22xp5_ASAP7_75t_SL g309 ( .A1(n_281), .A2(n_177), .B1(n_188), .B2(n_194), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_279), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_279), .Y(n_311) );
NOR2x1_ASAP7_75t_L g312 ( .A(n_264), .B(n_177), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_238), .B(n_192), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_238), .Y(n_314) );
NOR2xp67_ASAP7_75t_L g315 ( .A(n_275), .B(n_203), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_274), .B(n_200), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_258), .B(n_200), .Y(n_317) );
BUFx10_ASAP7_75t_L g318 ( .A(n_304), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_266), .B(n_200), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_239), .Y(n_320) );
NOR2xp67_ASAP7_75t_L g321 ( .A(n_292), .B(n_206), .Y(n_321) );
CKINVDCx16_ASAP7_75t_R g322 ( .A(n_283), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_304), .Y(n_323) );
BUFx4_ASAP7_75t_SL g324 ( .A(n_290), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_239), .Y(n_325) );
INVx3_ASAP7_75t_SL g326 ( .A(n_290), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_240), .A2(n_200), .B1(n_217), .B2(n_231), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_278), .B(n_200), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_247), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_260), .Y(n_330) );
BUFx12f_ASAP7_75t_L g331 ( .A(n_267), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_278), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_269), .B(n_220), .Y(n_333) );
INVx6_ASAP7_75t_SL g334 ( .A(n_260), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_244), .B(n_200), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_252), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_261), .B(n_218), .Y(n_337) );
NOR2xp33_ASAP7_75t_R g338 ( .A(n_267), .B(n_217), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_252), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_240), .A2(n_225), .B1(n_226), .B2(n_220), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_251), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_254), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_301), .B(n_225), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_255), .A2(n_230), .B(n_178), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_254), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_241), .A2(n_209), .B(n_178), .Y(n_346) );
INVx8_ASAP7_75t_L g347 ( .A(n_286), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_269), .A2(n_220), .B1(n_179), .B2(n_180), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_251), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_260), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_246), .B(n_220), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_282), .B(n_179), .Y(n_352) );
NAND2x1p5_ASAP7_75t_L g353 ( .A(n_263), .B(n_179), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_288), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_237), .A2(n_209), .B1(n_180), .B2(n_184), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_294), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_296), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_247), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_263), .A2(n_184), .B(n_189), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_297), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_299), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_329), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_309), .A2(n_289), .B1(n_300), .B2(n_286), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_332), .A2(n_250), .B1(n_272), .B2(n_300), .C(n_298), .Y(n_364) );
AO21x1_ASAP7_75t_L g365 ( .A1(n_342), .A2(n_189), .B(n_205), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_320), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_323), .A2(n_286), .B1(n_242), .B2(n_265), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_320), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_342), .A2(n_286), .B1(n_270), .B2(n_303), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_324), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_325), .B(n_302), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_325), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_329), .Y(n_373) );
OAI221xp5_ASAP7_75t_L g374 ( .A1(n_312), .A2(n_326), .B1(n_315), .B2(n_355), .C(n_354), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_336), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_336), .Y(n_376) );
A2O1A1Ixp33_ASAP7_75t_L g377 ( .A1(n_357), .A2(n_277), .B(n_242), .C(n_265), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_326), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_345), .B(n_271), .Y(n_379) );
INVx3_ASAP7_75t_L g380 ( .A(n_329), .Y(n_380) );
INVx3_ASAP7_75t_L g381 ( .A(n_329), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g382 ( .A1(n_347), .A2(n_265), .B1(n_242), .B2(n_271), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_345), .B(n_271), .Y(n_383) );
INVx4_ASAP7_75t_L g384 ( .A(n_347), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_357), .B(n_243), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_339), .A2(n_153), .B1(n_158), .B2(n_243), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_343), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_343), .B(n_256), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_308), .B(n_256), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_361), .B(n_243), .Y(n_390) );
BUFx12f_ASAP7_75t_L g391 ( .A(n_331), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_314), .A2(n_284), .B1(n_243), .B2(n_245), .Y(n_392) );
BUFx4f_ASAP7_75t_L g393 ( .A(n_347), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_308), .B(n_284), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_331), .Y(n_395) );
OAI22xp33_ASAP7_75t_L g396 ( .A1(n_314), .A2(n_243), .B1(n_205), .B2(n_159), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_310), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_384), .B(n_361), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_387), .B(n_314), .Y(n_399) );
AOI221xp5_ASAP7_75t_SL g400 ( .A1(n_363), .A2(n_360), .B1(n_356), .B2(n_352), .C(n_313), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_372), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_374), .A2(n_314), .B1(n_318), .B2(n_308), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_378), .Y(n_403) );
AND2x4_ASAP7_75t_L g404 ( .A(n_384), .B(n_314), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_387), .B(n_356), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_369), .A2(n_344), .B(n_346), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_364), .A2(n_349), .B1(n_341), .B2(n_305), .C(n_307), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_372), .Y(n_408) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_366), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_376), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_363), .A2(n_347), .B1(n_360), .B2(n_327), .Y(n_411) );
BUFx3_ASAP7_75t_L g412 ( .A(n_393), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_374), .A2(n_318), .B1(n_307), .B2(n_305), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_376), .A2(n_316), .B1(n_310), .B2(n_321), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_366), .B(n_305), .Y(n_415) );
OAI211xp5_ASAP7_75t_SL g416 ( .A1(n_364), .A2(n_337), .B(n_318), .C(n_328), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_366), .B(n_307), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_368), .B(n_311), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_378), .Y(n_419) );
AOI22xp33_ASAP7_75t_SL g420 ( .A1(n_370), .A2(n_322), .B1(n_338), .B2(n_341), .Y(n_420) );
AOI22xp33_ASAP7_75t_SL g421 ( .A1(n_370), .A2(n_351), .B1(n_358), .B2(n_311), .Y(n_421) );
AOI22xp33_ASAP7_75t_SL g422 ( .A1(n_393), .A2(n_351), .B1(n_358), .B2(n_306), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_368), .B(n_351), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_368), .Y(n_424) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_367), .A2(n_319), .B1(n_317), .B2(n_335), .C(n_340), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_369), .A2(n_329), .B1(n_353), .B2(n_333), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_388), .A2(n_333), .B1(n_353), .B2(n_334), .Y(n_427) );
BUFx10_ASAP7_75t_L g428 ( .A(n_398), .Y(n_428) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_407), .A2(n_382), .B1(n_377), .B2(n_393), .C(n_395), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_416), .A2(n_388), .B1(n_393), .B2(n_384), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_405), .B(n_375), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_401), .B(n_375), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_413), .A2(n_371), .B1(n_375), .B2(n_382), .Y(n_433) );
OR2x2_ASAP7_75t_SL g434 ( .A(n_403), .B(n_391), .Y(n_434) );
CKINVDCx16_ASAP7_75t_R g435 ( .A(n_412), .Y(n_435) );
AOI222xp33_ASAP7_75t_L g436 ( .A1(n_402), .A2(n_391), .B1(n_388), .B2(n_371), .C1(n_384), .C2(n_383), .Y(n_436) );
A2O1A1Ixp33_ASAP7_75t_L g437 ( .A1(n_412), .A2(n_379), .B(n_383), .C(n_390), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_419), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_424), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g440 ( .A1(n_412), .A2(n_391), .B1(n_362), .B2(n_381), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g441 ( .A1(n_398), .A2(n_380), .B1(n_362), .B2(n_381), .Y(n_441) );
OAI222xp33_ASAP7_75t_L g442 ( .A1(n_426), .A2(n_379), .B1(n_396), .B2(n_385), .C1(n_390), .C2(n_397), .Y(n_442) );
AOI221xp5_ASAP7_75t_SL g443 ( .A1(n_411), .A2(n_386), .B1(n_396), .B2(n_385), .C(n_397), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_401), .B(n_397), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_426), .A2(n_381), .B1(n_373), .B2(n_380), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_409), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_408), .B(n_362), .Y(n_447) );
OAI221xp5_ASAP7_75t_L g448 ( .A1(n_420), .A2(n_386), .B1(n_392), .B2(n_353), .C(n_381), .Y(n_448) );
OAI22xp33_ASAP7_75t_L g449 ( .A1(n_405), .A2(n_362), .B1(n_380), .B2(n_373), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_424), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_409), .Y(n_451) );
AOI33xp33_ASAP7_75t_L g452 ( .A1(n_421), .A2(n_204), .A3(n_235), .B1(n_232), .B2(n_221), .B3(n_219), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_408), .B(n_394), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_398), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_398), .A2(n_380), .B1(n_373), .B2(n_389), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_404), .B(n_373), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_410), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_399), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_409), .Y(n_459) );
BUFx3_ASAP7_75t_L g460 ( .A(n_404), .Y(n_460) );
NAND4xp25_ASAP7_75t_SL g461 ( .A(n_422), .B(n_365), .C(n_13), .D(n_14), .Y(n_461) );
OAI22xp33_ASAP7_75t_L g462 ( .A1(n_411), .A2(n_334), .B1(n_389), .B2(n_394), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_458), .B(n_431), .Y(n_463) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_436), .B(n_400), .C(n_410), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_438), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_434), .A2(n_427), .B1(n_404), .B2(n_399), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_432), .B(n_409), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_432), .B(n_409), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_457), .B(n_415), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_434), .B(n_404), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_457), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_439), .Y(n_472) );
OAI221xp5_ASAP7_75t_L g473 ( .A1(n_429), .A2(n_400), .B1(n_414), .B2(n_425), .C(n_406), .Y(n_473) );
AOI31xp33_ASAP7_75t_L g474 ( .A1(n_440), .A2(n_423), .A3(n_414), .B(n_415), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_439), .B(n_409), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_450), .B(n_418), .Y(n_476) );
OAI21x1_ASAP7_75t_L g477 ( .A1(n_445), .A2(n_365), .B(n_359), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_431), .B(n_418), .Y(n_478) );
AOI221x1_ASAP7_75t_L g479 ( .A1(n_437), .A2(n_423), .B1(n_159), .B2(n_417), .C(n_389), .Y(n_479) );
NAND4xp25_ASAP7_75t_SL g480 ( .A(n_430), .B(n_417), .C(n_13), .D(n_15), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_450), .B(n_12), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_454), .B(n_16), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g483 ( .A(n_452), .B(n_229), .C(n_223), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_444), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_444), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g486 ( .A1(n_461), .A2(n_394), .B1(n_389), .B2(n_211), .C(n_219), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_447), .B(n_16), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_447), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_460), .B(n_359), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_446), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_462), .A2(n_394), .B1(n_333), .B2(n_334), .Y(n_491) );
INVx4_ASAP7_75t_L g492 ( .A(n_428), .Y(n_492) );
INVx2_ASAP7_75t_SL g493 ( .A(n_428), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_460), .B(n_18), .Y(n_494) );
BUFx2_ASAP7_75t_L g495 ( .A(n_446), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_459), .Y(n_496) );
NAND4xp25_ASAP7_75t_L g497 ( .A(n_443), .B(n_19), .C(n_20), .D(n_227), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_451), .Y(n_498) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_435), .Y(n_499) );
NOR2x1_ASAP7_75t_L g500 ( .A(n_442), .B(n_350), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_459), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_451), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_453), .B(n_235), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_449), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_456), .B(n_21), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_428), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_456), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_456), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_455), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_435), .B(n_232), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_433), .A2(n_350), .B1(n_330), .B2(n_348), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_471), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_465), .B(n_448), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_463), .B(n_441), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_471), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_485), .B(n_443), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_499), .B(n_24), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_492), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_507), .B(n_30), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_472), .Y(n_520) );
NAND3xp33_ASAP7_75t_L g521 ( .A(n_497), .B(n_229), .C(n_223), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_467), .B(n_37), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_510), .Y(n_523) );
OR2x6_ASAP7_75t_L g524 ( .A(n_492), .B(n_350), .Y(n_524) );
OAI31xp33_ASAP7_75t_L g525 ( .A1(n_480), .A2(n_330), .A3(n_227), .B(n_221), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_472), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_467), .B(n_47), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_496), .Y(n_528) );
OAI21xp5_ASAP7_75t_SL g529 ( .A1(n_474), .A2(n_470), .B(n_497), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_476), .B(n_211), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_463), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_510), .Y(n_532) );
NOR2xp33_ASAP7_75t_R g533 ( .A(n_492), .B(n_51), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_488), .B(n_57), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_488), .B(n_60), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_484), .B(n_65), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_468), .B(n_66), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_496), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_468), .B(n_475), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_494), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_501), .Y(n_541) );
INVxp67_ASAP7_75t_SL g542 ( .A(n_495), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_475), .B(n_68), .Y(n_543) );
INVxp67_ASAP7_75t_L g544 ( .A(n_494), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_507), .B(n_69), .Y(n_545) );
NAND2x1p5_ASAP7_75t_L g546 ( .A(n_492), .B(n_330), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_476), .B(n_72), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_507), .B(n_73), .Y(n_548) );
BUFx2_ASAP7_75t_L g549 ( .A(n_495), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_508), .B(n_74), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_493), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_484), .B(n_80), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_501), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_490), .Y(n_554) );
BUFx3_ASAP7_75t_L g555 ( .A(n_493), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_490), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_498), .B(n_223), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_506), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_498), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_508), .B(n_223), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_487), .B(n_223), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_487), .B(n_481), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_502), .B(n_229), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_502), .Y(n_564) );
NAND3xp33_ASAP7_75t_L g565 ( .A(n_464), .B(n_229), .C(n_234), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_504), .B(n_229), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_504), .B(n_234), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_489), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_489), .B(n_234), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_478), .B(n_234), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_521), .A2(n_483), .B(n_479), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_526), .Y(n_572) );
AOI222xp33_ASAP7_75t_L g573 ( .A1(n_529), .A2(n_464), .B1(n_481), .B2(n_473), .C1(n_509), .C2(n_466), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g574 ( .A1(n_513), .A2(n_469), .B1(n_509), .B2(n_506), .C(n_482), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_526), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_531), .B(n_509), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_518), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_512), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_523), .B(n_482), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_532), .B(n_489), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_518), .Y(n_581) );
OAI31xp33_ASAP7_75t_L g582 ( .A1(n_525), .A2(n_483), .A3(n_505), .B(n_491), .Y(n_582) );
OAI21xp33_ASAP7_75t_L g583 ( .A1(n_533), .A2(n_500), .B(n_505), .Y(n_583) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_562), .A2(n_479), .B1(n_500), .B2(n_489), .Y(n_584) );
OAI21xp5_ASAP7_75t_L g585 ( .A1(n_565), .A2(n_486), .B(n_511), .Y(n_585) );
OAI221xp5_ASAP7_75t_L g586 ( .A1(n_517), .A2(n_503), .B1(n_234), .B2(n_248), .C(n_273), .Y(n_586) );
AOI222xp33_ASAP7_75t_L g587 ( .A1(n_544), .A2(n_477), .B1(n_248), .B2(n_280), .C1(n_257), .C2(n_259), .Y(n_587) );
AOI211xp5_ASAP7_75t_L g588 ( .A1(n_540), .A2(n_477), .B(n_280), .C(n_257), .Y(n_588) );
INVxp67_ASAP7_75t_SL g589 ( .A(n_557), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_512), .Y(n_590) );
AOI221x1_ASAP7_75t_L g591 ( .A1(n_547), .A2(n_273), .B1(n_291), .B2(n_259), .C(n_262), .Y(n_591) );
OAI32xp33_ASAP7_75t_L g592 ( .A1(n_551), .A2(n_245), .A3(n_291), .B1(n_262), .B2(n_268), .Y(n_592) );
AOI221x1_ASAP7_75t_L g593 ( .A1(n_561), .A2(n_268), .B1(n_287), .B2(n_245), .C(n_285), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_539), .B(n_287), .Y(n_594) );
NOR2xp67_ASAP7_75t_L g595 ( .A(n_558), .B(n_249), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_514), .A2(n_249), .B1(n_285), .B2(n_293), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_539), .B(n_249), .Y(n_597) );
AOI21xp33_ASAP7_75t_L g598 ( .A1(n_558), .A2(n_249), .B(n_285), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_515), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_514), .A2(n_249), .B1(n_285), .B2(n_293), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_556), .B(n_285), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_556), .B(n_293), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_564), .B(n_515), .Y(n_603) );
INVxp67_ASAP7_75t_SL g604 ( .A(n_557), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_520), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_536), .A2(n_293), .B1(n_295), .B2(n_535), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_549), .B(n_293), .Y(n_607) );
AOI221x1_ASAP7_75t_L g608 ( .A1(n_516), .A2(n_295), .B1(n_564), .B2(n_550), .C(n_519), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_520), .B(n_295), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_568), .B(n_295), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_554), .B(n_295), .Y(n_611) );
NOR2xp67_ASAP7_75t_SL g612 ( .A(n_536), .B(n_535), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_554), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_555), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_568), .B(n_559), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_559), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_555), .B(n_542), .Y(n_617) );
OAI211xp5_ASAP7_75t_L g618 ( .A1(n_549), .A2(n_522), .B(n_537), .C(n_527), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_534), .A2(n_546), .B1(n_524), .B2(n_522), .Y(n_619) );
AOI222xp33_ASAP7_75t_L g620 ( .A1(n_552), .A2(n_530), .B1(n_537), .B2(n_527), .C1(n_543), .C2(n_567), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_543), .Y(n_621) );
INVxp67_ASAP7_75t_SL g622 ( .A(n_563), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_528), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_572), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_615), .B(n_541), .Y(n_625) );
INVxp67_ASAP7_75t_SL g626 ( .A(n_589), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_574), .A2(n_552), .B1(n_553), .B2(n_566), .C(n_567), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_603), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g629 ( .A(n_583), .B(n_534), .Y(n_629) );
NOR2x1_ASAP7_75t_L g630 ( .A(n_577), .B(n_524), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_572), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_575), .Y(n_632) );
NOR4xp25_ASAP7_75t_SL g633 ( .A(n_586), .B(n_546), .C(n_524), .D(n_519), .Y(n_633) );
NOR2xp33_ASAP7_75t_R g634 ( .A(n_581), .B(n_570), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_575), .Y(n_635) );
OAI21xp33_ASAP7_75t_L g636 ( .A1(n_573), .A2(n_569), .B(n_566), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_578), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_623), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_589), .B(n_541), .Y(n_639) );
INVx3_ASAP7_75t_L g640 ( .A(n_623), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_615), .B(n_528), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_590), .Y(n_642) );
OAI21xp5_ASAP7_75t_SL g643 ( .A1(n_618), .A2(n_546), .B(n_550), .Y(n_643) );
NOR2xp67_ASAP7_75t_L g644 ( .A(n_571), .B(n_519), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_599), .Y(n_645) );
NOR3xp33_ASAP7_75t_SL g646 ( .A(n_582), .B(n_524), .C(n_570), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_604), .B(n_538), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_605), .Y(n_648) );
HAxp5_ASAP7_75t_SL g649 ( .A(n_596), .B(n_550), .CON(n_649), .SN(n_649) );
AOI21xp33_ASAP7_75t_L g650 ( .A1(n_579), .A2(n_563), .B(n_569), .Y(n_650) );
NAND2xp33_ASAP7_75t_SL g651 ( .A(n_612), .B(n_550), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_613), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_616), .Y(n_653) );
OAI221xp5_ASAP7_75t_L g654 ( .A1(n_585), .A2(n_538), .B1(n_545), .B2(n_548), .C(n_560), .Y(n_654) );
NAND2xp33_ASAP7_75t_SL g655 ( .A(n_619), .B(n_519), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_580), .B(n_560), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_622), .B(n_545), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_614), .B(n_548), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_576), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_630), .B(n_584), .Y(n_660) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_646), .A2(n_584), .B(n_595), .Y(n_661) );
AOI322xp5_ASAP7_75t_L g662 ( .A1(n_655), .A2(n_636), .A3(n_626), .B1(n_651), .B2(n_629), .C1(n_659), .C2(n_627), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_628), .B(n_617), .Y(n_663) );
NOR2xp33_ASAP7_75t_SL g664 ( .A(n_643), .B(n_621), .Y(n_664) );
XNOR2xp5_ASAP7_75t_L g665 ( .A(n_656), .B(n_594), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_656), .B(n_620), .Y(n_666) );
AND2x4_ASAP7_75t_L g667 ( .A(n_644), .B(n_608), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g668 ( .A(n_649), .B(n_588), .C(n_587), .Y(n_668) );
XOR2x2_ASAP7_75t_L g669 ( .A(n_658), .B(n_606), .Y(n_669) );
O2A1O1Ixp5_ASAP7_75t_L g670 ( .A1(n_655), .A2(n_592), .B(n_598), .C(n_607), .Y(n_670) );
NOR2x1p5_ASAP7_75t_L g671 ( .A(n_649), .B(n_597), .Y(n_671) );
OAI322xp33_ASAP7_75t_L g672 ( .A1(n_639), .A2(n_600), .A3(n_602), .B1(n_601), .B2(n_609), .C1(n_611), .C2(n_610), .Y(n_672) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_640), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_637), .B(n_610), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_625), .B(n_593), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g676 ( .A1(n_651), .A2(n_591), .B1(n_654), .B2(n_650), .C(n_647), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_633), .A2(n_657), .B1(n_640), .B2(n_634), .Y(n_677) );
INVx1_ASAP7_75t_SL g678 ( .A(n_641), .Y(n_678) );
NAND3xp33_ASAP7_75t_SL g679 ( .A(n_662), .B(n_653), .C(n_652), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_660), .A2(n_640), .B(n_652), .Y(n_680) );
INVx1_ASAP7_75t_SL g681 ( .A(n_665), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_666), .B(n_645), .Y(n_682) );
O2A1O1Ixp5_ASAP7_75t_L g683 ( .A1(n_660), .A2(n_642), .B(n_648), .C(n_638), .Y(n_683) );
XNOR2xp5_ASAP7_75t_L g684 ( .A(n_671), .B(n_641), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_674), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_668), .A2(n_624), .B1(n_631), .B2(n_632), .Y(n_686) );
NAND4xp25_ASAP7_75t_L g687 ( .A(n_661), .B(n_632), .C(n_638), .D(n_635), .Y(n_687) );
OAI22xp5_ASAP7_75t_SL g688 ( .A1(n_676), .A2(n_635), .B1(n_677), .B2(n_667), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_663), .B(n_669), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_664), .A2(n_670), .B1(n_673), .B2(n_678), .C(n_675), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_673), .A2(n_671), .B1(n_664), .B2(n_668), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_672), .A2(n_671), .B1(n_643), .B2(n_660), .Y(n_692) );
INVxp67_ASAP7_75t_SL g693 ( .A(n_673), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g694 ( .A(n_662), .B(n_660), .C(n_676), .Y(n_694) );
NOR3xp33_ASAP7_75t_L g695 ( .A(n_694), .B(n_688), .C(n_692), .Y(n_695) );
CKINVDCx5p33_ASAP7_75t_R g696 ( .A(n_681), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_683), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_682), .B(n_689), .Y(n_698) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_690), .A2(n_686), .B1(n_693), .B2(n_685), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_695), .A2(n_679), .B(n_691), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_696), .Y(n_701) );
OR2x2_ASAP7_75t_L g702 ( .A(n_698), .B(n_687), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_701), .Y(n_703) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_702), .Y(n_704) );
INVx1_ASAP7_75t_SL g705 ( .A(n_703), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_705), .A2(n_700), .B1(n_704), .B2(n_697), .Y(n_706) );
AOI211xp5_ASAP7_75t_L g707 ( .A1(n_706), .A2(n_684), .B(n_680), .C(n_699), .Y(n_707) );
endmodule