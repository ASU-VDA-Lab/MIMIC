module fake_netlist_5_916_n_5557 (n_137, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_619, n_408, n_61, n_664, n_376, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_667, n_515, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_649, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_629, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_668, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_650, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_636, n_600, n_660, n_223, n_392, n_158, n_655, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_662, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_661, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_614, n_663, n_50, n_337, n_430, n_313, n_631, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_613, n_241, n_637, n_357, n_598, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_638, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_648, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_159, n_334, n_599, n_541, n_391, n_434, n_645, n_539, n_175, n_538, n_666, n_262, n_238, n_639, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_5557);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_619;
input n_408;
input n_61;
input n_664;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_667;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_649;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_629;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_668;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_650;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_661;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_638;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_666;
input n_262;
input n_238;
input n_639;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_5557;

wire n_924;
wire n_2253;
wire n_2417;
wire n_977;
wire n_2756;
wire n_4706;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_5287;
wire n_2327;
wire n_1488;
wire n_2899;
wire n_790;
wire n_5484;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_2395;
wire n_5161;
wire n_5512;
wire n_5207;
wire n_2347;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_2391;
wire n_5035;
wire n_5282;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_2059;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_671;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_1462;
wire n_4211;
wire n_3448;
wire n_3019;
wire n_2096;
wire n_877;
wire n_3776;
wire n_2530;
wire n_4517;
wire n_1696;
wire n_2483;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1285;
wire n_1860;
wire n_4615;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_5480;
wire n_2147;
wire n_3010;
wire n_2770;
wire n_4131;
wire n_5402;
wire n_2584;
wire n_3188;
wire n_5509;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_1242;
wire n_3283;
wire n_5469;
wire n_2323;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_5453;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_731;
wire n_5202;
wire n_1314;
wire n_1512;
wire n_1490;
wire n_3214;
wire n_2091;
wire n_1517;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_1449;
wire n_4678;
wire n_2032;
wire n_1566;
wire n_2587;
wire n_5406;
wire n_3947;
wire n_3490;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_5241;
wire n_882;
wire n_2384;
wire n_3156;
wire n_696;
wire n_3376;
wire n_5037;
wire n_4468;
wire n_3653;
wire n_3702;
wire n_1040;
wire n_4976;
wire n_2202;
wire n_2648;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_5398;
wire n_2276;
wire n_2089;
wire n_3420;
wire n_1561;
wire n_1165;
wire n_5144;
wire n_1034;
wire n_3361;
wire n_4758;
wire n_1600;
wire n_845;
wire n_4255;
wire n_1796;
wire n_901;
wire n_4484;
wire n_3668;
wire n_4237;
wire n_2934;
wire n_1672;
wire n_1880;
wire n_3550;
wire n_1626;
wire n_2079;
wire n_2238;
wire n_1151;
wire n_1405;
wire n_1706;
wire n_3418;
wire n_4901;
wire n_2859;
wire n_1075;
wire n_3395;
wire n_4917;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_2968;
wire n_1585;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_1599;
wire n_4421;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_4469;
wire n_4414;
wire n_5184;
wire n_4532;
wire n_3339;
wire n_3349;
wire n_3735;
wire n_2248;
wire n_3007;
wire n_1000;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_5463;
wire n_2100;
wire n_5236;
wire n_3310;
wire n_3487;
wire n_2258;
wire n_748;
wire n_1667;
wire n_1058;
wire n_838;
wire n_3983;
wire n_1053;
wire n_1224;
wire n_4405;
wire n_5433;
wire n_1926;
wire n_1331;
wire n_4195;
wire n_1014;
wire n_4969;
wire n_1241;
wire n_4504;
wire n_1385;
wire n_793;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_2987;
wire n_1527;
wire n_4567;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_2175;
wire n_5055;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_5397;
wire n_4471;
wire n_5031;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_3208;
wire n_3331;
wire n_2379;
wire n_4983;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_3649;
wire n_4302;
wire n_2514;
wire n_5189;
wire n_5381;
wire n_4786;
wire n_3257;
wire n_1027;
wire n_4160;
wire n_2293;
wire n_5516;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_1276;
wire n_1412;
wire n_3981;
wire n_1199;
wire n_1038;
wire n_1841;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_1711;
wire n_870;
wire n_1891;
wire n_5254;
wire n_3526;
wire n_2546;
wire n_965;
wire n_3790;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_4613;
wire n_4649;
wire n_1888;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_4028;
wire n_5479;
wire n_1690;
wire n_3819;
wire n_2449;
wire n_5083;
wire n_1194;
wire n_2297;
wire n_4186;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_2227;
wire n_4618;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_2876;
wire n_4099;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_2479;
wire n_1464;
wire n_4295;
wire n_5303;
wire n_1444;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_4697;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_4810;
wire n_3317;
wire n_1121;
wire n_4391;
wire n_949;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_1001;
wire n_1503;
wire n_4638;
wire n_1468;
wire n_3455;
wire n_5047;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_5346;
wire n_1994;
wire n_5517;
wire n_1195;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_5109;
wire n_2796;
wire n_757;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_3095;
wire n_2805;
wire n_1145;
wire n_4918;
wire n_1153;
wire n_3856;
wire n_741;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_1207;
wire n_5010;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_2857;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_940;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1596;
wire n_2947;
wire n_978;
wire n_4299;
wire n_4801;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_3515;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_1208;
wire n_3287;
wire n_3378;
wire n_5435;
wire n_1431;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_5373;
wire n_4294;
wire n_1732;
wire n_5279;
wire n_4125;
wire n_4232;
wire n_4949;
wire n_2941;
wire n_2457;
wire n_5493;
wire n_4790;
wire n_962;
wire n_723;
wire n_2536;
wire n_1336;
wire n_1758;
wire n_2952;
wire n_4847;
wire n_5321;
wire n_3058;
wire n_5096;
wire n_4365;
wire n_1878;
wire n_3505;
wire n_4610;
wire n_3730;
wire n_4489;
wire n_974;
wire n_727;
wire n_5210;
wire n_4967;
wire n_957;
wire n_4992;
wire n_3001;
wire n_3945;
wire n_4542;
wire n_2261;
wire n_2729;
wire n_3597;
wire n_1612;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_4534;
wire n_4500;
wire n_5014;
wire n_3185;
wire n_1300;
wire n_1127;
wire n_3523;
wire n_1785;
wire n_2829;
wire n_4597;
wire n_4329;
wire n_1006;
wire n_4087;
wire n_3811;
wire n_1270;
wire n_3200;
wire n_1664;
wire n_2231;
wire n_2017;
wire n_2604;
wire n_4257;
wire n_3453;
wire n_2390;
wire n_3213;
wire n_1041;
wire n_3077;
wire n_1562;
wire n_3474;
wire n_3984;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_1913;
wire n_1823;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_4189;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_3707;
wire n_1846;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_860;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_4687;
wire n_948;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_4037;
wire n_2922;
wire n_3499;
wire n_3275;
wire n_2645;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_1552;
wire n_3618;
wire n_2593;
wire n_5262;
wire n_3683;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_824;
wire n_1327;
wire n_4763;
wire n_1684;
wire n_3590;
wire n_5310;
wire n_815;
wire n_4594;
wire n_3424;
wire n_1381;
wire n_1037;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_5146;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_3171;
wire n_1437;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_5441;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_1123;
wire n_1467;
wire n_2163;
wire n_2254;
wire n_1382;
wire n_925;
wire n_3546;
wire n_2647;
wire n_1311;
wire n_1519;
wire n_950;
wire n_4443;
wire n_5461;
wire n_4507;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_3244;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_912;
wire n_968;
wire n_4452;
wire n_4348;
wire n_5430;
wire n_5362;
wire n_4355;
wire n_3494;
wire n_5050;
wire n_885;
wire n_5063;
wire n_5229;
wire n_2125;
wire n_3771;
wire n_5199;
wire n_683;
wire n_3110;
wire n_1057;
wire n_1051;
wire n_721;
wire n_1157;
wire n_3073;
wire n_4572;
wire n_5527;
wire n_802;
wire n_5416;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_1608;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_1305;
wire n_5266;
wire n_3178;
wire n_873;
wire n_5355;
wire n_2334;
wire n_690;
wire n_4521;
wire n_4488;
wire n_2289;
wire n_3051;
wire n_1343;
wire n_2783;
wire n_2263;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_1288;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_4519;
wire n_5551;
wire n_3715;
wire n_972;
wire n_3040;
wire n_1938;
wire n_1200;
wire n_2499;
wire n_3568;
wire n_5475;
wire n_3737;
wire n_1185;
wire n_991;
wire n_1967;
wire n_1329;
wire n_3255;
wire n_4856;
wire n_2997;
wire n_4400;
wire n_5168;
wire n_943;
wire n_3326;
wire n_3734;
wire n_4778;
wire n_2429;
wire n_883;
wire n_5322;
wire n_856;
wire n_1793;
wire n_4352;
wire n_4441;
wire n_918;
wire n_4761;
wire n_942;
wire n_1804;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_2364;
wire n_2533;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_5371;
wire n_2291;
wire n_4043;
wire n_1636;
wire n_3601;
wire n_5418;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_2094;
wire n_1096;
wire n_1575;
wire n_2393;
wire n_1697;
wire n_5316;
wire n_3831;
wire n_3801;
wire n_2043;
wire n_2751;
wire n_4893;
wire n_5032;
wire n_1549;
wire n_1934;
wire n_4948;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_1446;
wire n_4406;
wire n_2758;
wire n_1458;
wire n_1807;
wire n_2618;
wire n_5112;
wire n_5386;
wire n_2559;
wire n_763;
wire n_4748;
wire n_2295;
wire n_3931;
wire n_1219;
wire n_4010;
wire n_2840;
wire n_5017;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_2795;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_3380;
wire n_2098;
wire n_1296;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_5424;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_4728;
wire n_789;
wire n_4247;
wire n_4933;
wire n_4018;
wire n_3900;
wire n_1105;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_3872;
wire n_4336;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_836;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_3877;
wire n_2995;
wire n_5496;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_1102;
wire n_4052;
wire n_3459;
wire n_1499;
wire n_4398;
wire n_3155;
wire n_2633;
wire n_4954;
wire n_2435;
wire n_1392;
wire n_1164;
wire n_2097;
wire n_5460;
wire n_4304;
wire n_3911;
wire n_5333;
wire n_1303;
wire n_4431;
wire n_4192;
wire n_3736;
wire n_4805;
wire n_4885;
wire n_1661;
wire n_3565;
wire n_4701;
wire n_2575;
wire n_5040;
wire n_861;
wire n_1658;
wire n_1904;
wire n_1345;
wire n_1899;
wire n_1003;
wire n_2067;
wire n_2219;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_4631;
wire n_1726;
wire n_3035;
wire n_5194;
wire n_5464;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_3639;
wire n_708;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_1915;
wire n_1109;
wire n_5239;
wire n_1310;
wire n_2605;
wire n_4747;
wire n_5197;
wire n_1399;
wire n_1979;
wire n_2924;
wire n_4111;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_5305;
wire n_4538;
wire n_766;
wire n_1117;
wire n_2754;
wire n_687;
wire n_1742;
wire n_5376;
wire n_2489;
wire n_5204;
wire n_2012;
wire n_1291;
wire n_4094;
wire n_3503;
wire n_2866;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_4150;
wire n_827;
wire n_4878;
wire n_1703;
wire n_1650;
wire n_1137;
wire n_3934;
wire n_4985;
wire n_3922;
wire n_3846;
wire n_2103;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_850;
wire n_3074;
wire n_1999;
wire n_2372;
wire n_3673;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_2430;
wire n_2433;
wire n_3293;
wire n_5508;
wire n_4022;
wire n_1531;
wire n_840;
wire n_1334;
wire n_4852;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_2817;
wire n_3139;
wire n_5292;
wire n_2598;
wire n_4601;
wire n_2687;
wire n_1120;
wire n_1890;
wire n_714;
wire n_4220;
wire n_1944;
wire n_909;
wire n_1497;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_4515;
wire n_4351;
wire n_5264;
wire n_3126;
wire n_4403;
wire n_1981;
wire n_1663;
wire n_1718;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_5504;
wire n_1518;
wire n_4223;
wire n_1281;
wire n_1889;
wire n_1489;
wire n_5025;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_1569;
wire n_2188;
wire n_756;
wire n_1429;
wire n_4644;
wire n_4456;
wire n_5060;
wire n_5334;
wire n_2448;
wire n_4346;
wire n_3170;
wire n_2748;
wire n_3311;
wire n_3272;
wire n_2898;
wire n_2717;
wire n_1861;
wire n_760;
wire n_3628;
wire n_3691;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_2573;
wire n_4435;
wire n_2939;
wire n_3807;
wire n_2447;
wire n_4764;
wire n_886;
wire n_1221;
wire n_5394;
wire n_2774;
wire n_1707;
wire n_853;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_751;
wire n_4827;
wire n_2488;
wire n_3477;
wire n_5421;
wire n_2476;
wire n_704;
wire n_4399;
wire n_2781;
wire n_5309;
wire n_2778;
wire n_771;
wire n_4782;
wire n_1520;
wire n_4363;
wire n_2887;
wire n_1287;
wire n_4864;
wire n_1262;
wire n_2691;
wire n_1411;
wire n_3054;
wire n_4335;
wire n_2526;
wire n_2703;
wire n_2167;
wire n_5428;
wire n_3391;
wire n_4259;
wire n_5541;
wire n_2709;
wire n_5543;
wire n_816;
wire n_1536;
wire n_4865;
wire n_4056;
wire n_1344;
wire n_4564;
wire n_1246;
wire n_3840;
wire n_1339;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_2173;
wire n_1842;
wire n_871;
wire n_3738;
wire n_685;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_1555;
wire n_3245;
wire n_4417;
wire n_4899;
wire n_796;
wire n_2119;
wire n_1502;
wire n_2552;
wire n_2157;
wire n_1012;
wire n_5411;
wire n_2453;
wire n_4798;
wire n_1525;
wire n_740;
wire n_3509;
wire n_3352;
wire n_3076;
wire n_3535;
wire n_2182;
wire n_1061;
wire n_3251;
wire n_2931;
wire n_5185;
wire n_1193;
wire n_3118;
wire n_3511;
wire n_1226;
wire n_3443;
wire n_2146;
wire n_1487;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_781;
wire n_3521;
wire n_5379;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_1515;
wire n_2918;
wire n_3232;
wire n_1673;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_3114;
wire n_3125;
wire n_4981;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_4430;
wire n_4081;
wire n_1103;
wire n_3132;
wire n_4407;
wire n_3951;
wire n_4894;
wire n_3238;
wire n_3210;
wire n_2036;
wire n_3267;
wire n_4995;
wire n_695;
wire n_5524;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_3884;
wire n_3726;
wire n_805;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_3577;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1741;
wire n_1160;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_3347;
wire n_1074;
wire n_3216;
wire n_1621;
wire n_3809;
wire n_2113;
wire n_1448;
wire n_4288;
wire n_3567;
wire n_5066;
wire n_1634;
wire n_3939;
wire n_5401;
wire n_4241;
wire n_3321;
wire n_3212;
wire n_1433;
wire n_2256;
wire n_3152;
wire n_5106;
wire n_5468;
wire n_2920;
wire n_4265;
wire n_1186;
wire n_5319;
wire n_1018;
wire n_2247;
wire n_713;
wire n_1622;
wire n_1180;
wire n_3705;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_5455;
wire n_2268;
wire n_3778;
wire n_5337;
wire n_3304;
wire n_1378;
wire n_3912;
wire n_1729;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_5223;
wire n_3795;
wire n_5020;
wire n_4419;
wire n_4477;
wire n_3179;
wire n_3256;
wire n_2386;
wire n_1501;
wire n_3086;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_1099;
wire n_2568;
wire n_5364;
wire n_1738;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_1021;
wire n_4639;
wire n_3713;
wire n_3663;
wire n_5046;
wire n_5166;
wire n_3246;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_819;
wire n_5088;
wire n_2302;
wire n_5457;
wire n_951;
wire n_5532;
wire n_1494;
wire n_2069;
wire n_3434;
wire n_1806;
wire n_933;
wire n_1563;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_755;
wire n_4243;
wire n_4982;
wire n_3695;
wire n_4330;
wire n_2482;
wire n_2677;
wire n_5544;
wire n_3832;
wire n_3987;
wire n_902;
wire n_5352;
wire n_4991;
wire n_5538;
wire n_1698;
wire n_2329;
wire n_1098;
wire n_2142;
wire n_5410;
wire n_3332;
wire n_1135;
wire n_3048;
wire n_3937;
wire n_2203;
wire n_4525;
wire n_1243;
wire n_3782;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_3786;
wire n_2888;
wire n_3638;
wire n_5503;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_2306;
wire n_3022;
wire n_4264;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_5129;
wire n_2149;
wire n_1078;
wire n_5500;
wire n_3060;
wire n_4276;
wire n_5219;
wire n_3013;
wire n_1984;
wire n_5170;
wire n_2408;
wire n_5320;
wire n_1877;
wire n_3049;
wire n_1723;
wire n_5107;
wire n_4485;
wire n_4626;
wire n_1036;
wire n_1097;
wire n_798;
wire n_2659;
wire n_1414;
wire n_4975;
wire n_1852;
wire n_3089;
wire n_2470;
wire n_5405;
wire n_3985;
wire n_5253;
wire n_1391;
wire n_670;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_2551;
wire n_1587;
wire n_2682;
wire n_813;
wire n_1284;
wire n_3440;
wire n_1748;
wire n_4569;
wire n_2699;
wire n_4897;
wire n_888;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_5491;
wire n_2615;
wire n_3940;
wire n_1064;
wire n_858;
wire n_2985;
wire n_691;
wire n_5065;
wire n_2753;
wire n_1582;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_5492;
wire n_3141;
wire n_5084;
wire n_3164;
wire n_3570;
wire n_5260;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_5328;
wire n_3936;
wire n_4503;
wire n_3507;
wire n_3821;
wire n_2700;
wire n_1211;
wire n_3367;
wire n_4464;
wire n_907;
wire n_3096;
wire n_3496;
wire n_4114;
wire n_989;
wire n_2544;
wire n_2356;
wire n_892;
wire n_4556;
wire n_5454;
wire n_2620;
wire n_1581;
wire n_4089;
wire n_2919;
wire n_4327;
wire n_953;
wire n_4218;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_2757;
wire n_963;
wire n_1052;
wire n_954;
wire n_4353;
wire n_2042;
wire n_884;
wire n_1754;
wire n_1623;
wire n_2921;
wire n_2720;
wire n_1854;
wire n_4990;
wire n_5529;
wire n_1856;
wire n_4959;
wire n_4161;
wire n_832;
wire n_1319;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_1387;
wire n_4466;
wire n_2262;
wire n_2462;
wire n_1532;
wire n_3625;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_686;
wire n_2837;
wire n_847;
wire n_4844;
wire n_2979;
wire n_5257;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_702;
wire n_2548;
wire n_822;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_4388;
wire n_4206;
wire n_1538;
wire n_1779;
wire n_4738;
wire n_1369;
wire n_3909;
wire n_3207;
wire n_3944;
wire n_809;
wire n_4434;
wire n_4837;
wire n_3042;
wire n_1942;
wire n_2510;
wire n_4219;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_5012;
wire n_1293;
wire n_1876;
wire n_4620;
wire n_1810;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_2222;
wire n_3510;
wire n_3218;
wire n_2667;
wire n_3150;
wire n_747;
wire n_4325;
wire n_1733;
wire n_2413;
wire n_851;
wire n_843;
wire n_705;
wire n_3775;
wire n_4133;
wire n_678;
wire n_4184;
wire n_5203;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_4379;
wire n_2181;
wire n_1829;
wire n_4030;
wire n_4490;
wire n_3138;
wire n_4397;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_1734;
wire n_4820;
wire n_3770;
wire n_1308;
wire n_5094;
wire n_4938;
wire n_4179;
wire n_3469;
wire n_5336;
wire n_677;
wire n_2723;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_5548;
wire n_3855;
wire n_1008;
wire n_2054;
wire n_5339;
wire n_1559;
wire n_4931;
wire n_1765;
wire n_3158;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_3113;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_2856;
wire n_1832;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_3828;
wire n_3288;
wire n_5514;
wire n_4404;
wire n_5091;
wire n_1509;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_878;
wire n_5486;
wire n_1306;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_906;
wire n_919;
wire n_4356;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_1740;
wire n_1586;
wire n_4291;
wire n_5403;
wire n_4386;
wire n_4149;
wire n_1492;
wire n_1692;
wire n_2982;
wire n_2481;
wire n_3545;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_1095;
wire n_1614;
wire n_2339;
wire n_4637;
wire n_4935;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_3741;
wire n_3410;
wire n_2029;
wire n_995;
wire n_1609;
wire n_5298;
wire n_1887;
wire n_4413;
wire n_1073;
wire n_2346;
wire n_3990;
wire n_4493;
wire n_3475;
wire n_1215;
wire n_1592;
wire n_2882;
wire n_1721;
wire n_2338;
wire n_3672;
wire n_5290;
wire n_3197;
wire n_3109;
wire n_2721;
wire n_1043;
wire n_5095;
wire n_3002;
wire n_5324;
wire n_3897;
wire n_1159;
wire n_3845;
wire n_2081;
wire n_4570;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_2418;
wire n_2179;
wire n_1416;
wire n_1724;
wire n_2521;
wire n_3458;
wire n_1420;
wire n_3330;
wire n_1132;
wire n_4606;
wire n_4774;
wire n_2477;
wire n_3887;
wire n_4093;
wire n_1486;
wire n_4672;
wire n_3519;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_4766;
wire n_2896;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_1927;
wire n_1349;
wire n_4460;
wire n_1031;
wire n_3645;
wire n_3223;
wire n_3929;
wire n_834;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1965;
wire n_1902;
wire n_1941;
wire n_5501;
wire n_3938;
wire n_5377;
wire n_2878;
wire n_874;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_3189;
wire n_2066;
wire n_993;
wire n_3154;
wire n_1551;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4349;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_1084;
wire n_970;
wire n_1935;
wire n_3366;
wire n_1534;
wire n_1351;
wire n_2696;
wire n_4863;
wire n_1205;
wire n_3242;
wire n_3525;
wire n_3486;
wire n_2405;
wire n_3995;
wire n_2088;
wire n_2953;
wire n_4036;
wire n_921;
wire n_5100;
wire n_1795;
wire n_2578;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_5367;
wire n_2656;
wire n_1080;
wire n_1274;
wire n_3524;
wire n_5034;
wire n_1708;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2092;
wire n_2075;
wire n_3658;
wire n_1776;
wire n_4807;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_1757;
wire n_890;
wire n_1919;
wire n_960;
wire n_4230;
wire n_3419;
wire n_1290;
wire n_1047;
wire n_2053;
wire n_1958;
wire n_1252;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_1808;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_5003;
wire n_5252;
wire n_967;
wire n_2731;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_1357;
wire n_3979;
wire n_4582;
wire n_2998;
wire n_4684;
wire n_4840;
wire n_3162;
wire n_983;
wire n_2760;
wire n_3377;
wire n_3749;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_762;
wire n_1283;
wire n_5325;
wire n_2637;
wire n_5375;
wire n_4384;
wire n_4423;
wire n_4096;
wire n_2881;
wire n_1203;
wire n_3282;
wire n_821;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_4996;
wire n_2475;
wire n_4598;
wire n_5064;
wire n_4478;
wire n_2646;
wire n_5536;
wire n_1605;
wire n_5173;
wire n_1228;
wire n_3920;
wire n_4890;
wire n_5027;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_828;
wire n_779;
wire n_4106;
wire n_3717;
wire n_2743;
wire n_2675;
wire n_1439;
wire n_3052;
wire n_5215;
wire n_945;
wire n_3743;
wire n_1932;
wire n_4721;
wire n_984;
wire n_694;
wire n_1983;
wire n_4029;
wire n_1594;
wire n_900;
wire n_3870;
wire n_4496;
wire n_3529;
wire n_1977;
wire n_1147;
wire n_2153;
wire n_4338;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_1470;
wire n_1735;
wire n_2318;
wire n_833;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_3442;
wire n_1201;
wire n_1114;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_669;
wire n_1176;
wire n_1149;
wire n_1020;
wire n_5121;
wire n_1824;
wire n_1917;
wire n_3386;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_5555;
wire n_2446;
wire n_3488;
wire n_1035;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_4668;
wire n_4953;
wire n_5466;
wire n_3898;
wire n_849;
wire n_1786;
wire n_5284;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_2627;
wire n_4759;
wire n_1413;
wire n_801;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_3552;
wire n_875;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_2361;
wire n_1173;
wire n_1603;
wire n_1401;
wire n_969;
wire n_4113;
wire n_1019;
wire n_1998;
wire n_4686;
wire n_5530;
wire n_3759;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_3933;
wire n_3206;
wire n_5506;
wire n_3966;
wire n_5243;
wire n_5449;
wire n_1702;
wire n_5221;
wire n_4183;
wire n_778;
wire n_1122;
wire n_4068;
wire n_4872;
wire n_4233;
wire n_3192;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_2649;
wire n_1187;
wire n_1929;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_3324;
wire n_1174;
wire n_3914;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_3742;
wire n_2252;
wire n_4819;
wire n_1685;
wire n_917;
wire n_1714;
wire n_1541;
wire n_2576;
wire n_4900;
wire n_3390;
wire n_1573;
wire n_3746;
wire n_2373;
wire n_1713;
wire n_3817;
wire n_2745;
wire n_1253;
wire n_1737;
wire n_774;
wire n_2493;
wire n_4930;
wire n_5276;
wire n_1059;
wire n_1133;
wire n_5078;
wire n_4537;
wire n_2885;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_4282;
wire n_3485;
wire n_4180;
wire n_3839;
wire n_1440;
wire n_5205;
wire n_3333;
wire n_2845;
wire n_4143;
wire n_4659;
wire n_2602;
wire n_4579;
wire n_4616;
wire n_1496;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_2401;
wire n_3135;
wire n_5476;
wire n_2003;
wire n_1457;
wire n_5446;
wire n_4895;
wire n_3573;
wire n_3148;
wire n_2264;
wire n_3534;
wire n_1482;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3438;
wire n_4098;
wire n_872;
wire n_1297;
wire n_4789;
wire n_1972;
wire n_2806;
wire n_1184;
wire n_2184;
wire n_5312;
wire n_985;
wire n_3217;
wire n_3425;
wire n_3404;
wire n_5111;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_676;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_1602;
wire n_1178;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_2065;
wire n_4017;
wire n_3397;
wire n_3740;
wire n_1081;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_703;
wire n_1318;
wire n_780;
wire n_2977;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_3600;
wire n_4134;
wire n_1388;
wire n_2836;
wire n_672;
wire n_1625;
wire n_2130;
wire n_5167;
wire n_898;
wire n_3239;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_1452;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_1326;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_4740;
wire n_5301;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_1192;
wire n_2221;
wire n_3576;
wire n_1024;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_4049;
wire n_941;
wire n_3862;
wire n_5214;
wire n_5487;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_5497;
wire n_4724;
wire n_1238;
wire n_1772;
wire n_752;
wire n_1476;
wire n_1108;
wire n_5526;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_4546;
wire n_862;
wire n_3584;
wire n_3756;
wire n_2889;
wire n_5021;
wire n_2772;
wire n_5444;
wire n_1675;
wire n_1924;
wire n_4382;
wire n_1554;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_5211;
wire n_5230;
wire n_2260;
wire n_5389;
wire n_1813;
wire n_4833;
wire n_3056;
wire n_2345;
wire n_1172;
wire n_5110;
wire n_1341;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_5425;
wire n_3289;
wire n_1973;
wire n_786;
wire n_1142;
wire n_2579;
wire n_1770;
wire n_4228;
wire n_4401;
wire n_1756;
wire n_1716;
wire n_2788;
wire n_2984;
wire n_3364;
wire n_1873;
wire n_3201;
wire n_1087;
wire n_3472;
wire n_2874;
wire n_5179;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_4968;
wire n_1272;
wire n_5030;
wire n_3949;
wire n_3543;
wire n_1247;
wire n_3050;
wire n_1478;
wire n_3903;
wire n_4834;
wire n_1210;
wire n_1364;
wire n_5272;
wire n_2742;
wire n_2183;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_5361;
wire n_4171;
wire n_4045;
wire n_1367;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_1460;
wire n_2834;
wire n_2531;
wire n_5015;
wire n_2702;
wire n_2030;
wire n_903;
wire n_3115;
wire n_4749;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_1404;
wire n_1794;
wire n_2234;
wire n_4804;
wire n_5545;
wire n_2209;
wire n_4270;
wire n_2797;
wire n_1255;
wire n_5152;
wire n_2321;
wire n_722;
wire n_3680;
wire n_844;
wire n_3497;
wire n_1601;
wire n_5409;
wire n_2940;
wire n_2612;
wire n_1495;
wire n_5128;
wire n_4566;
wire n_979;
wire n_2841;
wire n_3322;
wire n_4576;
wire n_846;
wire n_2427;
wire n_2505;
wire n_4061;
wire n_2070;
wire n_3250;
wire n_2594;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_5307;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_3112;
wire n_2349;
wire n_1379;
wire n_3874;
wire n_5415;
wire n_4676;
wire n_4544;
wire n_2170;
wire n_1091;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_4591;
wire n_3266;
wire n_4646;
wire n_1130;
wire n_4563;
wire n_4725;
wire n_2210;
wire n_4169;
wire n_5331;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_2426;
wire n_4320;
wire n_5341;
wire n_4881;
wire n_5271;
wire n_5089;
wire n_5263;
wire n_3613;
wire n_3444;
wire n_1181;
wire n_1505;
wire n_4012;
wire n_5518;
wire n_4636;
wire n_4584;
wire n_807;
wire n_3910;
wire n_4711;
wire n_835;
wire n_3319;
wire n_5240;
wire n_3335;
wire n_3413;
wire n_5495;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_1138;
wire n_5546;
wire n_927;
wire n_2689;
wire n_3259;
wire n_5482;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_3688;
wire n_3016;
wire n_1693;
wire n_5393;
wire n_2599;
wire n_904;
wire n_3338;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_4209;
wire n_1271;
wire n_1542;
wire n_5041;
wire n_1423;
wire n_1166;
wire n_1751;
wire n_5431;
wire n_1508;
wire n_785;
wire n_2200;
wire n_3261;
wire n_5026;
wire n_1161;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_1150;
wire n_5059;
wire n_5505;
wire n_3127;
wire n_1780;
wire n_3732;
wire n_4250;
wire n_5329;
wire n_1055;
wire n_3596;
wire n_4699;
wire n_3906;
wire n_4127;
wire n_880;
wire n_3297;
wire n_2683;
wire n_1370;
wire n_1360;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_4202;
wire n_5212;
wire n_5000;
wire n_2853;
wire n_1323;
wire n_688;
wire n_3766;
wire n_1353;
wire n_800;
wire n_2880;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_915;
wire n_864;
wire n_5420;
wire n_1264;
wire n_4412;
wire n_3599;
wire n_3407;
wire n_3621;
wire n_1580;
wire n_5234;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1607;
wire n_2538;
wire n_2105;
wire n_5259;
wire n_3163;
wire n_5440;
wire n_1118;
wire n_1686;
wire n_947;
wire n_3710;
wire n_4155;
wire n_1359;
wire n_2031;
wire n_3891;
wire n_1230;
wire n_4144;
wire n_2165;
wire n_929;
wire n_3379;
wire n_4374;
wire n_3532;
wire n_1124;
wire n_5131;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1257;
wire n_1182;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_4548;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_1016;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_1845;
wire n_2193;
wire n_2478;
wire n_5140;
wire n_4816;
wire n_1483;
wire n_2983;
wire n_3810;
wire n_1289;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_5306;
wire n_4483;
wire n_5342;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_2651;
wire n_4358;
wire n_5147;
wire n_3656;
wire n_2071;
wire n_2561;
wire n_2643;
wire n_1374;
wire n_4793;
wire n_4168;
wire n_3446;
wire n_955;
wire n_5511;
wire n_3028;
wire n_4806;
wire n_1146;
wire n_4350;
wire n_5533;
wire n_897;
wire n_5280;
wire n_1428;
wire n_1216;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1931;
wire n_4187;
wire n_1070;
wire n_4166;
wire n_5206;
wire n_1030;
wire n_3222;
wire n_1071;
wire n_1267;
wire n_1801;
wire n_5419;
wire n_1513;
wire n_2970;
wire n_2235;
wire n_673;
wire n_837;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_680;
wire n_1473;
wire n_3755;
wire n_4258;
wire n_4498;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_2506;
wire n_675;
wire n_4064;
wire n_4936;
wire n_5387;
wire n_1556;
wire n_1863;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_2944;
wire n_881;
wire n_2407;
wire n_4907;
wire n_5058;
wire n_3262;
wire n_1450;
wire n_5018;
wire n_4006;
wire n_4861;
wire n_1322;
wire n_3690;
wire n_889;
wire n_2358;
wire n_973;
wire n_5192;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_2370;
wire n_5159;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_736;
wire n_5097;
wire n_2750;
wire n_3899;
wire n_1278;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_4069;
wire n_2784;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_2557;
wire n_5300;
wire n_1248;
wire n_4850;
wire n_3781;
wire n_4813;
wire n_4912;
wire n_2590;
wire n_2330;
wire n_2942;
wire n_5525;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_944;
wire n_3889;
wire n_4256;
wire n_4224;
wire n_3508;
wire n_4024;
wire n_2218;
wire n_2267;
wire n_857;
wire n_2636;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_5400;
wire n_2759;
wire n_4415;
wire n_5552;
wire n_4702;
wire n_4252;
wire n_4457;
wire n_971;
wire n_5139;
wire n_1393;
wire n_2319;
wire n_3481;
wire n_5481;
wire n_2808;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_4491;
wire n_2930;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_2611;
wire n_4261;
wire n_1660;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_2698;
wire n_5043;
wire n_1662;
wire n_1481;
wire n_4001;
wire n_3047;
wire n_868;
wire n_2454;
wire n_4371;
wire n_914;
wire n_5281;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_5048;
wire n_5521;
wire n_5028;
wire n_1479;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_4194;
wire n_759;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1766;
wire n_1571;
wire n_3119;
wire n_4142;
wire n_1189;
wire n_4082;
wire n_3479;
wire n_4085;
wire n_4260;
wire n_4073;
wire n_1649;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_3279;
wire n_2621;
wire n_5073;
wire n_5024;
wire n_1537;
wire n_4262;
wire n_2671;
wire n_1798;
wire n_1790;
wire n_4720;
wire n_1647;
wire n_4685;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_1674;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_5515;
wire n_4014;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_2913;
wire n_2336;
wire n_1233;
wire n_1615;
wire n_4175;
wire n_2005;
wire n_1916;
wire n_4648;
wire n_1333;
wire n_5006;
wire n_1443;
wire n_946;
wire n_1539;
wire n_4892;
wire n_3823;
wire n_1866;
wire n_4173;
wire n_689;
wire n_738;
wire n_1624;
wire n_4970;
wire n_3816;
wire n_1279;
wire n_5404;
wire n_4108;
wire n_4486;
wire n_2960;
wire n_1090;
wire n_5438;
wire n_4627;
wire n_758;
wire n_2290;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_1049;
wire n_2145;
wire n_1639;
wire n_3030;
wire n_1068;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_5163;
wire n_2039;
wire n_4961;
wire n_3753;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_1362;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_3396;
wire n_1445;
wire n_4023;
wire n_4420;
wire n_1923;
wire n_5138;
wire n_1017;
wire n_5374;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1828;
wire n_2320;
wire n_1045;
wire n_5349;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_4640;
wire n_2583;
wire n_1033;
wire n_4396;
wire n_5127;
wire n_4367;
wire n_2087;
wire n_5485;
wire n_5216;
wire n_1009;
wire n_1989;
wire n_3818;
wire n_2523;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_1578;
wire n_3719;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_2725;
wire n_5175;
wire n_3883;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_773;
wire n_743;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_3466;
wire n_4962;
wire n_1237;
wire n_2595;
wire n_761;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_5171;
wire n_3586;
wire n_1390;
wire n_5554;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_5427;
wire n_3065;
wire n_4361;
wire n_1093;
wire n_5417;
wire n_4614;
wire n_1265;
wire n_2681;
wire n_3103;
wire n_765;
wire n_4945;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_1015;
wire n_1651;
wire n_2775;
wire n_4693;
wire n_5488;
wire n_1101;
wire n_1106;
wire n_4326;
wire n_3557;
wire n_2230;
wire n_5447;
wire n_5383;
wire n_4744;
wire n_2851;
wire n_4305;
wire n_1455;
wire n_767;
wire n_2490;
wire n_1407;
wire n_4213;
wire n_2849;
wire n_3692;
wire n_2204;
wire n_4929;
wire n_729;
wire n_1961;
wire n_4964;
wire n_911;
wire n_1430;
wire n_4802;
wire n_1354;
wire n_4139;
wire n_1044;
wire n_3029;
wire n_2508;
wire n_4031;
wire n_2416;
wire n_5437;
wire n_3881;
wire n_2461;
wire n_2243;
wire n_4583;
wire n_4210;
wire n_5245;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_1611;
wire n_2368;
wire n_2890;
wire n_2554;
wire n_3698;
wire n_3927;
wire n_1082;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_716;
wire n_1630;
wire n_4891;
wire n_701;
wire n_1023;
wire n_803;
wire n_1092;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_3993;
wire n_4940;
wire n_5208;
wire n_1056;
wire n_3588;
wire n_2308;
wire n_4590;
wire n_4830;
wire n_5231;
wire n_5237;
wire n_4664;
wire n_3860;
wire n_1029;
wire n_1206;
wire n_5456;
wire n_3160;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_3847;
wire n_4946;
wire n_1346;
wire n_4906;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_5390;
wire n_1060;
wire n_5347;
wire n_2824;
wire n_3033;
wire n_3298;
wire n_2440;
wire n_4883;
wire n_1386;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_2333;
wire n_2916;
wire n_4297;
wire n_1632;
wire n_1085;
wire n_1066;
wire n_3800;
wire n_2403;
wire n_5407;
wire n_4608;
wire n_5232;
wire n_2792;
wire n_2870;
wire n_3991;
wire n_1112;
wire n_3134;
wire n_4172;
wire n_4791;
wire n_4536;
wire n_5149;
wire n_2463;
wire n_5151;
wire n_4773;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_2472;
wire n_4611;
wire n_4755;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_1719;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2309;
wire n_2948;
wire n_1560;
wire n_5494;
wire n_4362;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_4422;
wire n_2589;
wire n_1363;
wire n_1301;
wire n_3482;
wire n_2233;
wire n_1312;
wire n_804;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_5228;
wire n_1504;
wire n_3956;
wire n_5323;
wire n_3572;
wire n_992;
wire n_4215;
wire n_4280;
wire n_3375;
wire n_4047;
wire n_5471;
wire n_842;
wire n_5434;
wire n_2082;
wire n_1643;
wire n_3167;
wire n_5350;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_5338;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3854;
wire n_2468;
wire n_1610;
wire n_1422;
wire n_1077;
wire n_3078;
wire n_894;
wire n_3253;
wire n_4027;
wire n_831;
wire n_2280;
wire n_4599;
wire n_3363;
wire n_4812;
wire n_1511;
wire n_3689;
wire n_2020;
wire n_4628;
wire n_1881;
wire n_988;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_3950;
wire n_4458;
wire n_4121;
wire n_1616;
wire n_5090;
wire n_4476;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_2303;
wire n_2810;
wire n_2747;
wire n_1848;
wire n_2126;
wire n_4573;
wire n_5289;
wire n_4118;
wire n_5513;
wire n_4803;
wire n_4079;
wire n_4091;
wire n_681;
wire n_1638;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_5132;
wire n_830;
wire n_5191;
wire n_3085;
wire n_1655;
wire n_749;
wire n_5359;
wire n_2574;
wire n_1134;
wire n_5293;
wire n_1358;
wire n_717;
wire n_4316;
wire n_939;
wire n_3697;
wire n_1232;
wire n_734;
wire n_2638;
wire n_4044;
wire n_4062;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_1338;
wire n_5510;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_2711;
wire n_5363;
wire n_5200;
wire n_1653;
wire n_1506;
wire n_2867;
wire n_990;
wire n_1894;
wire n_975;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_4253;
wire n_5356;
wire n_5369;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_770;
wire n_5255;
wire n_2852;
wire n_2392;
wire n_711;
wire n_3517;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_1834;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_1516;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_2409;
wire n_3402;
wire n_5295;
wire n_4679;
wire n_4115;
wire n_726;
wire n_4998;
wire n_2988;
wire n_1731;
wire n_818;
wire n_1970;
wire n_2766;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_2205;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_3401;
wire n_3226;
wire n_1410;
wire n_707;
wire n_3902;
wire n_4730;
wire n_937;
wire n_2779;
wire n_1584;
wire n_3654;
wire n_2164;
wire n_2115;
wire n_2232;
wire n_5327;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_5137;
wire n_2811;
wire n_3348;
wire n_895;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_5098;
wire n_1543;
wire n_1991;
wire n_2224;
wire n_732;
wire n_4743;
wire n_3805;
wire n_1067;
wire n_3825;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_2692;
wire n_2008;
wire n_4654;
wire n_5423;
wire n_799;
wire n_1213;
wire n_4733;
wire n_3792;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_1689;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_869;
wire n_3312;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_5069;
wire n_3285;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_684;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_2480;
wire n_2363;
wire n_4072;
wire n_916;
wire n_1115;
wire n_4781;
wire n_3606;
wire n_5004;
wire n_2550;
wire n_4424;
wire n_823;
wire n_725;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_3878;
wire n_4450;
wire n_3553;
wire n_719;
wire n_4746;
wire n_1683;
wire n_1530;
wire n_997;
wire n_932;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_1409;
wire n_3850;
wire n_788;
wire n_4459;
wire n_1268;
wire n_2996;
wire n_1320;
wire n_4050;
wire n_986;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_2102;
wire n_1063;
wire n_4853;
wire n_981;
wire n_867;
wire n_2422;
wire n_2239;
wire n_5256;
wire n_2950;
wire n_5220;
wire n_3852;
wire n_5178;
wire n_812;
wire n_4520;
wire n_2057;
wire n_4008;
wire n_5507;
wire n_905;
wire n_5077;
wire n_782;
wire n_3858;
wire n_1901;
wire n_4502;
wire n_3032;
wire n_4851;
wire n_1330;
wire n_3072;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_1745;
wire n_3924;
wire n_769;
wire n_4571;
wire n_2006;
wire n_934;
wire n_5314;
wire n_1618;
wire n_826;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_2535;
wire n_4205;
wire n_2726;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_1083;
wire n_4739;
wire n_2376;
wire n_5483;
wire n_3017;
wire n_787;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_4879;
wire n_5051;
wire n_930;
wire n_3926;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2854;
wire n_1701;
wire n_4181;
wire n_1550;
wire n_2764;
wire n_1498;
wire n_4225;
wire n_682;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_922;
wire n_1648;
wire n_4153;
wire n_5156;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_1769;
wire n_4783;
wire n_839;
wire n_2964;
wire n_3769;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_2442;
wire n_928;
wire n_1943;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_1396;
wire n_1348;
wire n_2883;
wire n_1752;
wire n_4182;
wire n_2912;
wire n_1315;
wire n_4825;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_5120;
wire n_5470;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_4839;
wire n_5222;
wire n_1028;
wire n_4016;
wire n_3435;
wire n_3575;
wire n_1546;
wire n_4231;
wire n_3165;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_4083;
wire n_1937;
wire n_4461;
wire n_3234;
wire n_5392;
wire n_745;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3024;
wire n_5443;
wire n_3512;
wire n_4939;
wire n_5169;
wire n_4389;
wire n_3930;
wire n_4448;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_2503;
wire n_1540;
wire n_1936;
wire n_5502;
wire n_2027;
wire n_2642;
wire n_720;
wire n_2500;
wire n_1918;
wire n_863;
wire n_4831;
wire n_2513;
wire n_2695;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_2414;
wire n_1402;
wire n_3662;
wire n_4319;
wire n_5474;
wire n_2229;
wire n_1397;
wire n_4596;
wire n_5413;
wire n_2004;
wire n_5412;
wire n_3694;
wire n_2586;
wire n_4726;
wire n_1398;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_1196;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_811;
wire n_4119;
wire n_3799;
wire n_4298;
wire n_5201;
wire n_4474;
wire n_1089;
wire n_5217;
wire n_1004;
wire n_2511;
wire n_1681;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_5490;
wire n_5029;
wire n_2704;
wire n_4214;
wire n_5158;
wire n_4884;
wire n_4366;
wire n_1251;
wire n_4009;
wire n_4580;
wire n_1263;
wire n_1126;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_1859;
wire n_1677;
wire n_5472;
wire n_2955;
wire n_4112;
wire n_4337;
wire n_4138;
wire n_5396;
wire n_1528;
wire n_5335;
wire n_1292;
wire n_2520;
wire n_1198;
wire n_956;
wire n_2134;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_1347;
wire n_5143;
wire n_4238;
wire n_1451;
wire n_1022;
wire n_2374;
wire n_1545;
wire n_859;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_2396;
wire n_1799;
wire n_854;
wire n_4734;
wire n_674;
wire n_1939;
wire n_2486;
wire n_4635;
wire n_1152;
wire n_3501;
wire n_1869;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_4242;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_1896;
wire n_3180;
wire n_5283;
wire n_5268;
wire n_1705;
wire n_4561;
wire n_2639;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_1261;
wire n_938;
wire n_3186;
wire n_4955;
wire n_1154;
wire n_5556;
wire n_5462;
wire n_4501;
wire n_3696;
wire n_1280;
wire n_3650;
wire n_2761;
wire n_3157;
wire n_709;
wire n_2537;
wire n_2144;
wire n_920;
wire n_2515;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_1949;
wire n_976;
wire n_1946;
wire n_2936;
wire n_775;
wire n_1484;
wire n_1328;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_4369;
wire n_5378;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_5542;
wire n_1831;
wire n_1598;
wire n_4394;
wire n_1850;
wire n_5519;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_5278;
wire n_2663;
wire n_1394;
wire n_2693;
wire n_3798;
wire n_4065;
wire n_5187;
wire n_4944;
wire n_2249;
wire n_2180;
wire n_926;
wire n_4135;
wire n_1218;
wire n_2632;
wire n_1547;
wire n_777;
wire n_1755;
wire n_958;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_4716;
wire n_4942;
wire n_2432;
wire n_1521;
wire n_3405;
wire n_4745;
wire n_2337;
wire n_1167;
wire n_1384;
wire n_3907;
wire n_5344;
wire n_923;
wire n_4629;
wire n_2932;
wire n_2980;
wire n_5225;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_4752;
wire n_5265;
wire n_1750;
wire n_1459;
wire n_3986;
wire n_4376;
wire n_4753;
wire n_4552;
wire n_3885;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_1197;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_5126;
wire n_1039;
wire n_2214;
wire n_3427;
wire n_2055;
wire n_4067;
wire n_1403;
wire n_5553;
wire n_4042;
wire n_4176;
wire n_4385;
wire n_3320;
wire n_5009;
wire n_2688;
wire n_5368;
wire n_1202;
wire n_1463;
wire n_3651;
wire n_4333;
wire n_3359;
wire n_2865;
wire n_2706;
wire n_5499;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_4815;
wire n_4246;
wire n_3580;
wire n_2139;
wire n_4609;
wire n_5291;
wire n_5114;
wire n_2674;
wire n_1565;
wire n_4088;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_4472;
wire n_4462;
wire n_3433;
wire n_1072;
wire n_5288;
wire n_2305;
wire n_5540;
wire n_2450;
wire n_3447;
wire n_3305;
wire n_4148;
wire n_4151;
wire n_1712;
wire n_3528;
wire n_4373;
wire n_4934;
wire n_5218;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_4630;
wire n_5408;
wire n_4643;
wire n_4331;
wire n_3989;
wire n_4475;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_1775;
wire n_3296;
wire n_1368;
wire n_2762;
wire n_4683;
wire n_5366;
wire n_728;
wire n_1162;
wire n_1847;
wire n_2767;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_5477;
wire n_5451;
wire n_3923;
wire n_931;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_1544;
wire n_5086;
wire n_1629;
wire n_2801;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_1997;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_5053;
wire n_1259;
wire n_4553;
wire n_706;
wire n_746;
wire n_784;
wire n_3978;
wire n_4809;
wire n_5226;
wire n_1244;
wire n_1925;
wire n_3660;
wire n_1815;
wire n_1788;
wire n_2491;
wire n_5079;
wire n_913;
wire n_3833;
wire n_865;
wire n_697;
wire n_1222;
wire n_1679;
wire n_4841;
wire n_776;
wire n_2022;
wire n_3814;
wire n_1415;
wire n_2592;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_3513;
wire n_3133;
wire n_4645;
wire n_1191;
wire n_2992;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_2517;
wire n_3128;
wire n_5426;
wire n_744;
wire n_2631;
wire n_2178;
wire n_1767;
wire n_1529;
wire n_2469;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_5531;
wire n_3000;
wire n_5429;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_1837;
wire n_1839;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_2875;
wire n_936;
wire n_1500;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_5448;
wire n_3471;
wire n_5432;
wire n_999;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_1656;
wire n_3564;
wire n_1158;
wire n_3988;
wire n_3457;
wire n_1678;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_5445;
wire n_3630;
wire n_3271;
wire n_4771;
wire n_908;
wire n_4086;
wire n_2412;
wire n_4814;
wire n_724;
wire n_2084;
wire n_1781;
wire n_3648;
wire n_3075;
wire n_3173;
wire n_5332;
wire n_5108;
wire n_4692;
wire n_959;
wire n_3031;
wire n_3701;
wire n_3243;
wire n_1773;
wire n_1169;
wire n_2666;
wire n_3385;
wire n_2171;
wire n_4708;
wire n_2768;
wire n_2314;
wire n_4826;
wire n_3343;
wire n_2420;
wire n_1079;
wire n_5489;
wire n_1593;
wire n_3767;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_4589;
wire n_5057;
wire n_4578;
wire n_1640;
wire n_2162;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_3221;
wire n_742;
wire n_750;
wire n_5436;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_2359;
wire n_3674;
wire n_5286;
wire n_3502;
wire n_3098;
wire n_1383;
wire n_5013;
wire n_2312;
wire n_3015;
wire n_1171;
wire n_1920;
wire n_1065;
wire n_5439;
wire n_4147;
wire n_2048;
wire n_3607;
wire n_4925;
wire n_1921;
wire n_1309;
wire n_4974;
wire n_1800;
wire n_1548;
wire n_4932;
wire n_1421;
wire n_4510;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_3276;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_1119;
wire n_1240;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_4285;
wire n_4651;
wire n_700;
wire n_4818;
wire n_4514;
wire n_1366;
wire n_4800;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_1568;
wire n_2110;
wire n_1332;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_1591;
wire n_2033;
wire n_4341;
wire n_1682;
wire n_4312;
wire n_2628;
wire n_3399;
wire n_1249;
wire n_1111;
wire n_2132;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_4140;
wire n_3675;
wire n_5092;
wire n_1140;
wire n_891;
wire n_3387;
wire n_5186;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_2831;
wire n_1456;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_4832;
wire n_4207;
wire n_987;
wire n_4545;
wire n_3037;
wire n_4868;
wire n_1885;
wire n_2452;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_5238;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_1849;
wire n_1131;
wire n_5054;
wire n_2467;
wire n_1094;
wire n_2288;
wire n_4063;
wire n_5399;
wire n_1209;
wire n_3592;
wire n_4650;
wire n_4888;
wire n_5326;
wire n_1435;
wire n_879;
wire n_3394;
wire n_4874;
wire n_3793;
wire n_4669;
wire n_4339;
wire n_1645;
wire n_4041;
wire n_5459;
wire n_2858;
wire n_4060;
wire n_996;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_2128;
wire n_5528;
wire n_3097;
wire n_5391;
wire n_4541;
wire n_3824;
wire n_5422;
wire n_3388;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_5523;
wire n_3465;
wire n_1316;
wire n_4796;
wire n_1438;
wire n_3589;
wire n_952;
wire n_2534;
wire n_1229;
wire n_4799;
wire n_5153;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_2789;
wire n_4775;
wire n_2216;
wire n_5044;
wire n_1897;
wire n_764;
wire n_1424;
wire n_5365;
wire n_2933;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_5354;
wire n_4455;
wire n_2328;
wire n_4248;
wire n_5452;
wire n_4754;
wire n_4554;
wire n_4845;
wire n_3053;
wire n_1299;
wire n_3893;
wire n_1141;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_1699;
wire n_3334;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_5535;
wire n_1432;
wire n_3875;
wire n_5370;
wire n_4003;
wire n_5372;
wire n_5299;
wire n_2402;
wire n_4301;
wire n_841;
wire n_1050;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_1844;
wire n_3777;
wire n_4784;
wire n_2999;
wire n_1644;
wire n_5550;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_5209;
wire n_3080;
wire n_4199;
wire n_2701;
wire n_3362;
wire n_1631;
wire n_3105;
wire n_5478;
wire n_1179;
wire n_753;
wire n_1048;
wire n_4286;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_692;
wire n_820;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_3417;
wire n_1143;
wire n_1579;
wire n_4034;
wire n_1688;
wire n_3327;
wire n_5275;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_2755;
wire n_3237;
wire n_1992;
wire n_4402;
wire n_4239;
wire n_3400;
wire n_4550;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_3382;
wire n_3574;
wire n_5227;
wire n_2169;
wire n_1557;
wire n_4201;
wire n_896;
wire n_3316;
wire n_5242;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1730;
wire n_3603;
wire n_4123;
wire n_2192;
wire n_5520;
wire n_964;
wire n_3633;
wire n_4479;
wire n_1373;
wire n_2670;
wire n_1646;
wire n_1307;
wire n_4416;
wire n_3372;
wire n_4539;
wire n_814;
wire n_2707;
wire n_2471;
wire n_1472;
wire n_1671;
wire n_3230;
wire n_3342;
wire n_1062;
wire n_4682;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_1204;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_5458;
wire n_3861;
wire n_4736;
wire n_3780;
wire n_783;
wire n_1928;
wire n_5244;
wire n_5382;
wire n_1188;
wire n_3957;
wire n_5274;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_5384;
wire n_3608;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_2352;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_2619;
wire n_2444;
wire n_1110;
wire n_3123;
wire n_5056;
wire n_1088;
wire n_5249;
wire n_3393;
wire n_866;
wire n_5198;
wire n_5360;
wire n_5233;
wire n_4887;
wire n_4617;
wire n_5269;
wire n_3520;
wire n_2492;
wire n_4005;
wire n_1687;
wire n_1637;
wire n_4904;
wire n_1419;
wire n_693;
wire n_4792;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_1389;
wire n_1256;
wire n_4980;
wire n_1465;
wire n_4290;
wire n_5247;
wire n_1375;
wire n_3727;
wire n_5317;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_1597;
wire n_1659;
wire n_2431;
wire n_1371;
wire n_4956;
wire n_5380;
wire n_2206;
wire n_3182;
wire n_2564;
wire n_4947;
wire n_876;
wire n_4656;
wire n_1190;
wire n_3896;
wire n_3958;
wire n_3450;
wire n_966;
wire n_4729;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_1116;
wire n_2000;
wire n_1212;
wire n_2074;
wire n_3174;
wire n_982;
wire n_1453;
wire n_2217;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_3408;
wire n_899;
wire n_2722;
wire n_5388;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_1628;
wire n_3432;
wire n_1514;
wire n_1771;
wire n_1005;
wire n_679;
wire n_710;
wire n_3090;
wire n_2437;
wire n_3762;
wire n_1168;
wire n_2445;
wire n_1427;
wire n_1835;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_4529;
wire n_910;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_3972;
wire n_5539;
wire n_3308;
wire n_791;
wire n_1533;
wire n_5036;
wire n_5547;
wire n_4772;
wire n_3467;
wire n_4322;
wire n_1720;
wire n_2830;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_5273;
wire n_4677;
wire n_3901;
wire n_715;
wire n_1480;
wire n_5261;
wire n_3757;
wire n_3381;
wire n_5193;
wire n_1782;
wire n_2245;
wire n_4909;
wire n_1524;
wire n_1485;
wire n_810;
wire n_2965;
wire n_3635;
wire n_5022;
wire n_5005;
wire n_1144;
wire n_2814;
wire n_1570;
wire n_3882;
wire n_3046;
wire n_2213;
wire n_1170;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_855;
wire n_5534;
wire n_1461;
wire n_3204;
wire n_2136;
wire n_5174;
wire n_1273;
wire n_1822;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_1235;
wire n_4380;
wire n_980;
wire n_698;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1783;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_998;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_4880;
wire n_1907;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_1417;
wire n_1295;
wire n_5061;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_1762;
wire n_1013;
wire n_718;
wire n_3023;
wire n_4193;
wire n_4075;
wire n_3104;
wire n_4737;
wire n_3647;
wire n_825;
wire n_2819;
wire n_737;
wire n_5195;
wire n_3609;
wire n_4136;
wire n_1715;
wire n_1952;
wire n_4393;
wire n_3720;
wire n_4535;
wire n_733;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_4794;
wire n_3959;
wire n_792;
wire n_3140;
wire n_5246;
wire n_3724;
wire n_2104;
wire n_3011;
wire n_5164;
wire n_4196;
wire n_1425;
wire n_4592;
wire n_4675;
wire n_5340;
wire n_3069;
wire n_5498;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_5183;
wire n_3084;
wire n_1727;
wire n_2735;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_5549;
wire n_2411;
wire n_1046;
wire n_3761;
wire n_4889;
wire n_2014;
wire n_2986;
wire n_5442;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_4828;
wire n_5385;
wire n_4558;
wire n_2172;
wire n_4722;
wire n_1129;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_961;
wire n_2250;
wire n_1225;
wire n_4092;
wire n_3908;
wire n_2423;
wire n_3671;
wire n_994;
wire n_3344;
wire n_2194;
wire n_848;
wire n_4465;
wire n_3302;
wire n_5537;
wire n_5304;
wire n_1223;
wire n_2680;
wire n_5130;
wire n_1567;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_3842;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_1797;
wire n_2957;
wire n_2357;
wire n_1250;
wire n_3309;
wire n_772;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_1589;
wire n_4116;
wire n_2570;
wire n_1086;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_5473;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_2744;
wire n_4287;
wire n_2397;
wire n_2208;
wire n_3063;
wire n_5177;
wire n_3617;
wire n_1298;
wire n_1652;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_1676;
wire n_1113;
wire n_1277;
wire n_2591;
wire n_3384;
wire n_852;
wire n_4602;
wire n_5172;
wire n_4449;
wire n_1864;
wire n_5070;
wire n_1337;
wire n_4445;
wire n_699;
wire n_5414;
wire n_1627;
wire n_1245;
wire n_4870;
wire n_2438;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_3181;
wire n_2278;
wire n_4915;
wire n_5296;
wire n_2135;
wire n_5450;
wire n_3493;
wire n_5313;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_2823;
wire n_1076;
wire n_1408;
wire n_1761;
wire n_730;
wire n_5270;
wire n_795;
wire n_4345;
wire n_5188;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_1526;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_5465;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_712;
wire n_1583;
wire n_2826;
wire n_3539;
wire n_1042;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_4124;
wire n_5467;
wire n_5522;
wire n_4492;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_2225;
wire n_1507;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3853;
wire n_4216;
wire n_2019;
wire n_1340;
wire n_1558;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_1704;
wire n_3721;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1234;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_2614;
wire n_1032;
wire n_2991;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_3473;
wire n_4560;
wire n_5318;
wire n_2839;
wire n_1588;
wire n_5395;
wire n_2237;
wire n_3463;
wire n_3699;
wire n_5067;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_2728;
wire n_3857;

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_643),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_280),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_144),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_158),
.Y(n_672)
);

BUFx5_ASAP7_75t_L g673 ( 
.A(n_298),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_84),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_631),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_146),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_277),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_455),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_357),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_88),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_362),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_613),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_207),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_334),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_408),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_558),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_410),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_494),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_618),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_311),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_96),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_308),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_356),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_635),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_555),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_492),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_80),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_403),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_39),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_580),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_252),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_49),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_662),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_644),
.Y(n_704)
);

CKINVDCx14_ASAP7_75t_R g705 ( 
.A(n_525),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_30),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_188),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_391),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_137),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_211),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_256),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_578),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_474),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_338),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_42),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_467),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_475),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_205),
.Y(n_718)
);

CKINVDCx14_ASAP7_75t_R g719 ( 
.A(n_85),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_456),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_94),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_14),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_653),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_301),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_294),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_649),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_238),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_180),
.Y(n_728)
);

BUFx10_ASAP7_75t_L g729 ( 
.A(n_647),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_636),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_357),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_294),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_117),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_186),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_373),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_491),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_352),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_346),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_246),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_602),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_512),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_623),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_254),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_407),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_118),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_381),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_557),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_454),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_198),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_69),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_199),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_529),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_188),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_554),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_233),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_288),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_542),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_304),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_388),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_370),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_389),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_29),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_563),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_74),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_565),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_272),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_362),
.Y(n_767)
);

BUFx2_ASAP7_75t_SL g768 ( 
.A(n_113),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_639),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_358),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_84),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_615),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_646),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_147),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_526),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_458),
.Y(n_776)
);

INVxp33_ASAP7_75t_R g777 ( 
.A(n_19),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_638),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_201),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_240),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_338),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_521),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_637),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_172),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_667),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_376),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_291),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_626),
.Y(n_788)
);

BUFx10_ASAP7_75t_L g789 ( 
.A(n_622),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_534),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_311),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_211),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_290),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_659),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_264),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_184),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_39),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_661),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_432),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_405),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_243),
.Y(n_801)
);

BUFx5_ASAP7_75t_L g802 ( 
.A(n_304),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_547),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_581),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_341),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_24),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_645),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_276),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_634),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_535),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_185),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_651),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_197),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_251),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_26),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_245),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_451),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_663),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_450),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_161),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_231),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_640),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_648),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_206),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_11),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_329),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_65),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_605),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_593),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_465),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_628),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_599),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_13),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_81),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_108),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_488),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_665),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_206),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_390),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_232),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_274),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_594),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_560),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_587),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_589),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_478),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_90),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_228),
.Y(n_848)
);

BUFx10_ASAP7_75t_L g849 ( 
.A(n_20),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_668),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_276),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_498),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_505),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_264),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_420),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_482),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_534),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_12),
.Y(n_858)
);

CKINVDCx16_ASAP7_75t_R g859 ( 
.A(n_325),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_303),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_22),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_642),
.Y(n_862)
);

BUFx5_ASAP7_75t_L g863 ( 
.A(n_666),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_457),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_202),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_600),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_253),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_63),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_584),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_347),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_80),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_407),
.Y(n_872)
);

INVx1_ASAP7_75t_SL g873 ( 
.A(n_52),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_498),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_327),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_650),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_441),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_454),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_168),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_332),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_616),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_579),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_451),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_330),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_191),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_516),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_284),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_562),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_246),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_465),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_385),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_197),
.Y(n_892)
);

BUFx10_ASAP7_75t_L g893 ( 
.A(n_199),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_442),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_514),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_524),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_384),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_450),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_320),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_214),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_252),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_262),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_113),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_111),
.Y(n_904)
);

CKINVDCx16_ASAP7_75t_R g905 ( 
.A(n_162),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_633),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_654),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_545),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_161),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_395),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_434),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_467),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_358),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_25),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_58),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_25),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_522),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_224),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_553),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_256),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_171),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_177),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_341),
.Y(n_923)
);

BUFx10_ASAP7_75t_L g924 ( 
.A(n_540),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_255),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_99),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_514),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_166),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_583),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_31),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_70),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_477),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_475),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_528),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_481),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_244),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_102),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_356),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_46),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_510),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_160),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_462),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_310),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_272),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_397),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_446),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_487),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_588),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_114),
.Y(n_949)
);

BUFx10_ASAP7_75t_L g950 ( 
.A(n_74),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_115),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_408),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_470),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_170),
.Y(n_954)
);

BUFx5_ASAP7_75t_L g955 ( 
.A(n_469),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_333),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_656),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_585),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_76),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_156),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_184),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_12),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_402),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_133),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_95),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_496),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_141),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_81),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_484),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_391),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_106),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_632),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_493),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_367),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_424),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_45),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_484),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_283),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_97),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_320),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_388),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_426),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_93),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_529),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_590),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_462),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_507),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_131),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_417),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_344),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_627),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_82),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_457),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_261),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_260),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_319),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_137),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_564),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_122),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_210),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_598),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_250),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_293),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_541),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_69),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_346),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_177),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_156),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_360),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_46),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_22),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_23),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_520),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_364),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_148),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_0),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_354),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_556),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_378),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_518),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_351),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_455),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_310),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_533),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_510),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_11),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_66),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_415),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_287),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_508),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_507),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_511),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_239),
.Y(n_1033)
);

BUFx3_ASAP7_75t_L g1034 ( 
.A(n_3),
.Y(n_1034)
);

INVx1_ASAP7_75t_SL g1035 ( 
.A(n_571),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_657),
.Y(n_1036)
);

CKINVDCx16_ASAP7_75t_R g1037 ( 
.A(n_152),
.Y(n_1037)
);

INVx1_ASAP7_75t_SL g1038 ( 
.A(n_229),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_176),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_91),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_315),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_302),
.Y(n_1042)
);

CKINVDCx16_ASAP7_75t_R g1043 ( 
.A(n_7),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_533),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_652),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_447),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_610),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_270),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_54),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_463),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_351),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_606),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_285),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_352),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_171),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_179),
.Y(n_1056)
);

CKINVDCx16_ASAP7_75t_R g1057 ( 
.A(n_278),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_23),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_349),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_293),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_664),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_398),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_316),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_401),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_428),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_496),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_174),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_185),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_396),
.Y(n_1069)
);

CKINVDCx14_ASAP7_75t_R g1070 ( 
.A(n_528),
.Y(n_1070)
);

INVxp33_ASAP7_75t_L g1071 ( 
.A(n_51),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_314),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_322),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_512),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_160),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_103),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_504),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_82),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_641),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_497),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_108),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_487),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_655),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_503),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_577),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_329),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_617),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_79),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_434),
.Y(n_1089)
);

CKINVDCx14_ASAP7_75t_R g1090 ( 
.A(n_658),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_398),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_435),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_350),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_245),
.Y(n_1094)
);

CKINVDCx20_ASAP7_75t_R g1095 ( 
.A(n_331),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_370),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_502),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_121),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_130),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_515),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_630),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_552),
.Y(n_1102)
);

CKINVDCx11_ASAP7_75t_R g1103 ( 
.A(n_390),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_493),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_361),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_260),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_235),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_461),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_319),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_315),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_114),
.Y(n_1111)
);

BUFx8_ASAP7_75t_SL g1112 ( 
.A(n_289),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_386),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_53),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_24),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_515),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_500),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_326),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_331),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_263),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_403),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_187),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_472),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_472),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_535),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_420),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_122),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_314),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_28),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_221),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_344),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_100),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_660),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_485),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_225),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_222),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_141),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_253),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_470),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_259),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_611),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_448),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_404),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_569),
.Y(n_1144)
);

BUFx10_ASAP7_75t_L g1145 ( 
.A(n_32),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_222),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_136),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_174),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_77),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_612),
.Y(n_1150)
);

INVx1_ASAP7_75t_SL g1151 ( 
.A(n_324),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_603),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_476),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_297),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_405),
.Y(n_1155)
);

CKINVDCx16_ASAP7_75t_R g1156 ( 
.A(n_332),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_270),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_244),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_540),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_328),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_300),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_271),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_440),
.Y(n_1163)
);

BUFx10_ASAP7_75t_L g1164 ( 
.A(n_198),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_65),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_364),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_162),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_500),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_257),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_266),
.Y(n_1170)
);

INVxp67_ASAP7_75t_SL g1171 ( 
.A(n_807),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_673),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1112),
.Y(n_1173)
);

INVxp67_ASAP7_75t_SL g1174 ( 
.A(n_807),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_673),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_673),
.Y(n_1176)
);

INVxp67_ASAP7_75t_SL g1177 ( 
.A(n_823),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1103),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_673),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_673),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_673),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_673),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_673),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_673),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_802),
.Y(n_1185)
);

INVxp33_ASAP7_75t_L g1186 ( 
.A(n_1129),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_790),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_802),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_802),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_802),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_802),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_802),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_790),
.Y(n_1193)
);

CKINVDCx11_ASAP7_75t_R g1194 ( 
.A(n_849),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_802),
.Y(n_1195)
);

INVxp67_ASAP7_75t_SL g1196 ( 
.A(n_823),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_802),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_802),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_955),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_955),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_955),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_955),
.Y(n_1202)
);

INVxp33_ASAP7_75t_SL g1203 ( 
.A(n_824),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_705),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_719),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_955),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_955),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_955),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_955),
.Y(n_1209)
);

INVxp67_ASAP7_75t_SL g1210 ( 
.A(n_866),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_955),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_682),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_720),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_682),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_730),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_720),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_700),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_700),
.Y(n_1218)
);

INVxp33_ASAP7_75t_L g1219 ( 
.A(n_824),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_703),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_703),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_726),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_726),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_672),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_742),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_720),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_713),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_720),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_742),
.Y(n_1229)
);

INVxp67_ASAP7_75t_SL g1230 ( 
.A(n_866),
.Y(n_1230)
);

CKINVDCx16_ASAP7_75t_R g1231 ( 
.A(n_859),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_761),
.Y(n_1232)
);

INVxp33_ASAP7_75t_L g1233 ( 
.A(n_938),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_765),
.Y(n_1234)
);

INVxp67_ASAP7_75t_L g1235 ( 
.A(n_938),
.Y(n_1235)
);

INVxp33_ASAP7_75t_SL g1236 ( 
.A(n_1015),
.Y(n_1236)
);

INVxp67_ASAP7_75t_L g1237 ( 
.A(n_1015),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_765),
.Y(n_1238)
);

INVxp67_ASAP7_75t_L g1239 ( 
.A(n_1155),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_773),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_773),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_794),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_794),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_764),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_809),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_809),
.Y(n_1246)
);

INVxp67_ASAP7_75t_SL g1247 ( 
.A(n_730),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_812),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_720),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1070),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_859),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_812),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_730),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_818),
.Y(n_1254)
);

CKINVDCx16_ASAP7_75t_R g1255 ( 
.A(n_905),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_818),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_829),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_829),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_842),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_842),
.Y(n_1260)
);

CKINVDCx16_ASAP7_75t_R g1261 ( 
.A(n_905),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_720),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_811),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1155),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_729),
.Y(n_1265)
);

INVxp33_ASAP7_75t_SL g1266 ( 
.A(n_768),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_811),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_811),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_811),
.Y(n_1269)
);

CKINVDCx16_ASAP7_75t_R g1270 ( 
.A(n_1037),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_811),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_811),
.Y(n_1272)
);

INVxp67_ASAP7_75t_SL g1273 ( 
.A(n_820),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_783),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_820),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1037),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_876),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_820),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_820),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_876),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_820),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_881),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1043),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_774),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_768),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_881),
.Y(n_1286)
);

INVxp33_ASAP7_75t_SL g1287 ( 
.A(n_671),
.Y(n_1287)
);

CKINVDCx14_ASAP7_75t_R g1288 ( 
.A(n_1090),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_882),
.Y(n_1289)
);

CKINVDCx20_ASAP7_75t_R g1290 ( 
.A(n_781),
.Y(n_1290)
);

CKINVDCx16_ASAP7_75t_R g1291 ( 
.A(n_1043),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_882),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1057),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1057),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_907),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_907),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_919),
.Y(n_1297)
);

INVxp67_ASAP7_75t_SL g1298 ( 
.A(n_820),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_919),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_929),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_929),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_836),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_836),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1156),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1156),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_991),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_991),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_674),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_676),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_683),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_836),
.Y(n_1311)
);

INVxp33_ASAP7_75t_L g1312 ( 
.A(n_1071),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1001),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_688),
.Y(n_1314)
);

INVx1_ASAP7_75t_SL g1315 ( 
.A(n_796),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1001),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_693),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_836),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1045),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1045),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1150),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1150),
.Y(n_1322)
);

CKINVDCx16_ASAP7_75t_R g1323 ( 
.A(n_849),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1152),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_678),
.Y(n_1325)
);

INVxp33_ASAP7_75t_L g1326 ( 
.A(n_678),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1152),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_696),
.Y(n_1328)
);

CKINVDCx16_ASAP7_75t_R g1329 ( 
.A(n_849),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_708),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_708),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_708),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_745),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_745),
.Y(n_1334)
);

INVxp67_ASAP7_75t_L g1335 ( 
.A(n_679),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_697),
.Y(n_1336)
);

INVxp33_ASAP7_75t_L g1337 ( 
.A(n_679),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_745),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_756),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_756),
.Y(n_1340)
);

INVxp67_ASAP7_75t_SL g1341 ( 
.A(n_836),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_756),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_766),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_766),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_766),
.Y(n_1345)
);

INVxp67_ASAP7_75t_SL g1346 ( 
.A(n_836),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_729),
.Y(n_1347)
);

INVxp67_ASAP7_75t_SL g1348 ( 
.A(n_902),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_841),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_841),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_841),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_860),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_860),
.Y(n_1353)
);

INVxp67_ASAP7_75t_SL g1354 ( 
.A(n_902),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_860),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_940),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_940),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_940),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_698),
.Y(n_1359)
);

INVxp33_ASAP7_75t_SL g1360 ( 
.A(n_699),
.Y(n_1360)
);

INVxp33_ASAP7_75t_SL g1361 ( 
.A(n_701),
.Y(n_1361)
);

INVxp67_ASAP7_75t_L g1362 ( 
.A(n_681),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_966),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_966),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_966),
.Y(n_1365)
);

BUFx5_ASAP7_75t_L g1366 ( 
.A(n_729),
.Y(n_1366)
);

INVxp67_ASAP7_75t_SL g1367 ( 
.A(n_902),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_825),
.Y(n_1368)
);

INVxp33_ASAP7_75t_SL g1369 ( 
.A(n_702),
.Y(n_1369)
);

INVxp33_ASAP7_75t_L g1370 ( 
.A(n_681),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1005),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_827),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1005),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1005),
.Y(n_1374)
);

NOR2xp67_ASAP7_75t_L g1375 ( 
.A(n_838),
.B(n_0),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1034),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_707),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_861),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_709),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1034),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_902),
.Y(n_1381)
);

INVxp33_ASAP7_75t_SL g1382 ( 
.A(n_710),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1034),
.Y(n_1383)
);

INVxp33_ASAP7_75t_SL g1384 ( 
.A(n_714),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1048),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1048),
.Y(n_1386)
);

INVxp33_ASAP7_75t_SL g1387 ( 
.A(n_716),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1048),
.Y(n_1388)
);

INVxp67_ASAP7_75t_SL g1389 ( 
.A(n_902),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_717),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_718),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1089),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_884),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_898),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_725),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1089),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1089),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_727),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1104),
.Y(n_1399)
);

NOR2xp67_ASAP7_75t_L g1400 ( 
.A(n_932),
.B(n_1),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1104),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1104),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_731),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_723),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_723),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_723),
.Y(n_1406)
);

INVxp33_ASAP7_75t_L g1407 ( 
.A(n_684),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_804),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_804),
.Y(n_1409)
);

INVxp33_ASAP7_75t_L g1410 ( 
.A(n_684),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_732),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_733),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_804),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_902),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1167),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1167),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1167),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1167),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1167),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_909),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1167),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_685),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_685),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_690),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_690),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_692),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_692),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_736),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_706),
.Y(n_1429)
);

INVxp67_ASAP7_75t_SL g1430 ( 
.A(n_689),
.Y(n_1430)
);

INVxp33_ASAP7_75t_SL g1431 ( 
.A(n_739),
.Y(n_1431)
);

INVxp67_ASAP7_75t_SL g1432 ( 
.A(n_689),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_706),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_729),
.Y(n_1434)
);

CKINVDCx16_ASAP7_75t_R g1435 ( 
.A(n_849),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_916),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_711),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_711),
.Y(n_1438)
);

INVxp67_ASAP7_75t_SL g1439 ( 
.A(n_695),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_789),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_715),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_715),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1042),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_677),
.Y(n_1444)
);

INVxp67_ASAP7_75t_L g1445 ( 
.A(n_721),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_721),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_734),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_734),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1069),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_677),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_735),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_743),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_735),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_737),
.Y(n_1454)
);

CKINVDCx20_ASAP7_75t_R g1455 ( 
.A(n_1075),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_737),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_744),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_751),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_751),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_752),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_752),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_758),
.Y(n_1462)
);

CKINVDCx16_ASAP7_75t_R g1463 ( 
.A(n_893),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_758),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_746),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_748),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_759),
.Y(n_1467)
);

INVxp33_ASAP7_75t_SL g1468 ( 
.A(n_749),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_750),
.Y(n_1469)
);

INVxp67_ASAP7_75t_SL g1470 ( 
.A(n_695),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_759),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_1081),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_677),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_760),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_760),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_791),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_791),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_800),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_893),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_800),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_810),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_810),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_814),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_814),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_817),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_817),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_834),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_834),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_846),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_846),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_753),
.Y(n_1491)
);

CKINVDCx20_ASAP7_75t_R g1492 ( 
.A(n_1082),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_1095),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_847),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1111),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_847),
.Y(n_1496)
);

INVxp67_ASAP7_75t_L g1497 ( 
.A(n_851),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_851),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_852),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_680),
.Y(n_1500)
);

INVxp67_ASAP7_75t_SL g1501 ( 
.A(n_757),
.Y(n_1501)
);

CKINVDCx20_ASAP7_75t_R g1502 ( 
.A(n_1114),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_852),
.Y(n_1503)
);

CKINVDCx20_ASAP7_75t_R g1504 ( 
.A(n_1123),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1157),
.Y(n_1505)
);

INVxp67_ASAP7_75t_SL g1506 ( 
.A(n_757),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_855),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_855),
.Y(n_1508)
);

INVxp67_ASAP7_75t_L g1509 ( 
.A(n_856),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_856),
.Y(n_1510)
);

INVxp33_ASAP7_75t_SL g1511 ( 
.A(n_755),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_857),
.Y(n_1512)
);

INVxp33_ASAP7_75t_SL g1513 ( 
.A(n_762),
.Y(n_1513)
);

INVxp33_ASAP7_75t_L g1514 ( 
.A(n_857),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_767),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_680),
.Y(n_1516)
);

INVxp33_ASAP7_75t_L g1517 ( 
.A(n_864),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_864),
.Y(n_1518)
);

INVxp33_ASAP7_75t_SL g1519 ( 
.A(n_770),
.Y(n_1519)
);

CKINVDCx16_ASAP7_75t_R g1520 ( 
.A(n_893),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_680),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_789),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_865),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_865),
.Y(n_1524)
);

INVx1_ASAP7_75t_SL g1525 ( 
.A(n_670),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_871),
.Y(n_1526)
);

INVxp67_ASAP7_75t_SL g1527 ( 
.A(n_837),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_871),
.Y(n_1528)
);

CKINVDCx16_ASAP7_75t_R g1529 ( 
.A(n_893),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_878),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_878),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_885),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_885),
.Y(n_1533)
);

INVxp67_ASAP7_75t_L g1534 ( 
.A(n_887),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_887),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_891),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_891),
.Y(n_1537)
);

CKINVDCx16_ASAP7_75t_R g1538 ( 
.A(n_924),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_894),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_894),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_895),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_771),
.Y(n_1542)
);

CKINVDCx16_ASAP7_75t_R g1543 ( 
.A(n_924),
.Y(n_1543)
);

INVxp67_ASAP7_75t_SL g1544 ( 
.A(n_837),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_895),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_776),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_901),
.Y(n_1547)
);

BUFx8_ASAP7_75t_SL g1548 ( 
.A(n_906),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_901),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_913),
.B(n_1),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_687),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_913),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_779),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_780),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_782),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_687),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_918),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_687),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_784),
.Y(n_1559)
);

INVxp67_ASAP7_75t_SL g1560 ( 
.A(n_1087),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_724),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_724),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_918),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_935),
.Y(n_1564)
);

CKINVDCx16_ASAP7_75t_R g1565 ( 
.A(n_924),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_935),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_936),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_936),
.Y(n_1568)
);

INVxp67_ASAP7_75t_SL g1569 ( 
.A(n_1087),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_724),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_943),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_943),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_951),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_786),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_951),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_728),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_787),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_953),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_953),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_954),
.Y(n_1580)
);

INVxp67_ASAP7_75t_SL g1581 ( 
.A(n_850),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_954),
.Y(n_1582)
);

INVxp33_ASAP7_75t_SL g1583 ( 
.A(n_793),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_728),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1213),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1525),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1273),
.B(n_850),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1274),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1312),
.B(n_789),
.Y(n_1589)
);

INVx5_ASAP7_75t_L g1590 ( 
.A(n_1274),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1274),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_1274),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1213),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1251),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1216),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1216),
.Y(n_1596)
);

INVx5_ASAP7_75t_L g1597 ( 
.A(n_1274),
.Y(n_1597)
);

BUFx8_ASAP7_75t_L g1598 ( 
.A(n_1187),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1226),
.Y(n_1599)
);

INVx5_ASAP7_75t_L g1600 ( 
.A(n_1521),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1278),
.B(n_1144),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1265),
.B(n_1347),
.Y(n_1602)
);

BUFx6f_ASAP7_75t_L g1603 ( 
.A(n_1226),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1265),
.B(n_1144),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_1548),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1298),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1347),
.B(n_1434),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1251),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_L g1609 ( 
.A(n_1228),
.Y(n_1609)
);

BUFx3_ASAP7_75t_L g1610 ( 
.A(n_1215),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1302),
.Y(n_1611)
);

INVx2_ASAP7_75t_SL g1612 ( 
.A(n_1308),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_SL g1613 ( 
.A(n_1231),
.B(n_924),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1312),
.B(n_789),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1341),
.B(n_669),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1521),
.Y(n_1616)
);

BUFx8_ASAP7_75t_L g1617 ( 
.A(n_1187),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1346),
.B(n_675),
.Y(n_1618)
);

BUFx12f_ASAP7_75t_L g1619 ( 
.A(n_1194),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1581),
.B(n_948),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1288),
.B(n_950),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1348),
.B(n_686),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1215),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1171),
.B(n_1035),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1288),
.B(n_950),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1228),
.Y(n_1626)
);

INVx5_ASAP7_75t_L g1627 ( 
.A(n_1521),
.Y(n_1627)
);

BUFx6f_ASAP7_75t_L g1628 ( 
.A(n_1249),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1174),
.B(n_1085),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1354),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1367),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1389),
.B(n_694),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1430),
.B(n_704),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1434),
.B(n_1141),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1432),
.B(n_712),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1439),
.B(n_740),
.Y(n_1636)
);

BUFx6f_ASAP7_75t_L g1637 ( 
.A(n_1249),
.Y(n_1637)
);

AND2x6_ASAP7_75t_L g1638 ( 
.A(n_1180),
.B(n_783),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1470),
.B(n_747),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1177),
.B(n_1196),
.Y(n_1640)
);

BUFx8_ASAP7_75t_L g1641 ( 
.A(n_1479),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1501),
.B(n_754),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1506),
.B(n_763),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1293),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1414),
.Y(n_1645)
);

BUFx8_ASAP7_75t_SL g1646 ( 
.A(n_1548),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_SL g1647 ( 
.A(n_1255),
.B(n_950),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1440),
.B(n_728),
.Y(n_1648)
);

BUFx8_ASAP7_75t_L g1649 ( 
.A(n_1479),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1269),
.Y(n_1650)
);

BUFx6f_ASAP7_75t_L g1651 ( 
.A(n_1269),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1440),
.B(n_792),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_L g1653 ( 
.A(n_1279),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1390),
.B(n_950),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_L g1655 ( 
.A(n_1279),
.Y(n_1655)
);

INVx5_ASAP7_75t_L g1656 ( 
.A(n_1570),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1395),
.B(n_1145),
.Y(n_1657)
);

BUFx12f_ASAP7_75t_L g1658 ( 
.A(n_1194),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1398),
.B(n_1145),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_SL g1660 ( 
.A(n_1261),
.B(n_1145),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1522),
.B(n_792),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1281),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1527),
.B(n_769),
.Y(n_1663)
);

INVx5_ASAP7_75t_L g1664 ( 
.A(n_1570),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1522),
.B(n_792),
.Y(n_1665)
);

BUFx3_ASAP7_75t_L g1666 ( 
.A(n_1253),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1281),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1544),
.B(n_772),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1303),
.Y(n_1669)
);

INVx4_ASAP7_75t_L g1670 ( 
.A(n_1308),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1570),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1560),
.B(n_778),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1294),
.Y(n_1673)
);

INVx5_ASAP7_75t_L g1674 ( 
.A(n_1303),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1276),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1569),
.B(n_785),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1210),
.B(n_722),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1415),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1204),
.B(n_1145),
.Y(n_1679)
);

BUFx6f_ASAP7_75t_L g1680 ( 
.A(n_1311),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1311),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1304),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1247),
.B(n_867),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_1173),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1230),
.B(n_722),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1318),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1266),
.B(n_738),
.Y(n_1687)
);

INVx4_ASAP7_75t_L g1688 ( 
.A(n_1309),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1416),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1403),
.B(n_1428),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1266),
.B(n_738),
.Y(n_1691)
);

INVx2_ASAP7_75t_SL g1692 ( 
.A(n_1309),
.Y(n_1692)
);

INVx4_ASAP7_75t_L g1693 ( 
.A(n_1310),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1371),
.B(n_1164),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1371),
.B(n_1164),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1417),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1469),
.B(n_1164),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1253),
.B(n_1285),
.Y(n_1698)
);

BUFx3_ASAP7_75t_L g1699 ( 
.A(n_1330),
.Y(n_1699)
);

BUFx3_ASAP7_75t_L g1700 ( 
.A(n_1331),
.Y(n_1700)
);

AND2x6_ASAP7_75t_L g1701 ( 
.A(n_1180),
.B(n_783),
.Y(n_1701)
);

NOR2x1_ASAP7_75t_L g1702 ( 
.A(n_1262),
.B(n_783),
.Y(n_1702)
);

AND2x6_ASAP7_75t_L g1703 ( 
.A(n_1172),
.B(n_783),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1287),
.B(n_1583),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1287),
.B(n_741),
.Y(n_1705)
);

INVx5_ASAP7_75t_L g1706 ( 
.A(n_1381),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1469),
.B(n_1164),
.Y(n_1707)
);

INVx5_ASAP7_75t_L g1708 ( 
.A(n_1381),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1418),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1419),
.B(n_788),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1310),
.Y(n_1711)
);

BUFx3_ASAP7_75t_L g1712 ( 
.A(n_1332),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1204),
.B(n_1205),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1421),
.B(n_798),
.Y(n_1714)
);

INVx3_ASAP7_75t_L g1715 ( 
.A(n_1444),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1262),
.B(n_803),
.Y(n_1716)
);

INVx5_ASAP7_75t_L g1717 ( 
.A(n_1444),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1205),
.B(n_822),
.Y(n_1718)
);

CKINVDCx20_ASAP7_75t_R g1719 ( 
.A(n_1224),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1235),
.B(n_867),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1360),
.B(n_741),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1237),
.B(n_867),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1250),
.B(n_828),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1239),
.B(n_1333),
.Y(n_1724)
);

INVx5_ASAP7_75t_L g1725 ( 
.A(n_1450),
.Y(n_1725)
);

INVx5_ASAP7_75t_L g1726 ( 
.A(n_1450),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_SL g1727 ( 
.A(n_1270),
.B(n_775),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1250),
.B(n_831),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1263),
.B(n_832),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1263),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1267),
.B(n_843),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1267),
.B(n_844),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1268),
.B(n_845),
.Y(n_1733)
);

BUFx12f_ASAP7_75t_L g1734 ( 
.A(n_1173),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1276),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1283),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_L g1737 ( 
.A(n_1473),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_1473),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1268),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1516),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1271),
.B(n_862),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1360),
.B(n_826),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1334),
.B(n_1338),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1361),
.B(n_826),
.Y(n_1744)
);

BUFx3_ASAP7_75t_L g1745 ( 
.A(n_1339),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1271),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1361),
.B(n_1019),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1340),
.B(n_1342),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1343),
.B(n_874),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1272),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1272),
.B(n_869),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1275),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1344),
.B(n_874),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1283),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1305),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_SL g1756 ( 
.A(n_1291),
.B(n_873),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1275),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1345),
.B(n_874),
.Y(n_1758)
);

INVx5_ASAP7_75t_L g1759 ( 
.A(n_1516),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1551),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1175),
.Y(n_1761)
);

INVx5_ASAP7_75t_L g1762 ( 
.A(n_1551),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1556),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1305),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1176),
.B(n_888),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1193),
.Y(n_1766)
);

AND2x6_ASAP7_75t_L g1767 ( 
.A(n_1179),
.B(n_783),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1349),
.B(n_879),
.Y(n_1768)
);

BUFx6f_ASAP7_75t_L g1769 ( 
.A(n_1556),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1181),
.B(n_908),
.Y(n_1770)
);

BUFx12f_ASAP7_75t_L g1771 ( 
.A(n_1178),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1264),
.Y(n_1772)
);

INVx5_ASAP7_75t_L g1773 ( 
.A(n_1366),
.Y(n_1773)
);

INVx5_ASAP7_75t_L g1774 ( 
.A(n_1366),
.Y(n_1774)
);

BUFx6f_ASAP7_75t_L g1775 ( 
.A(n_1422),
.Y(n_1775)
);

INVx5_ASAP7_75t_L g1776 ( 
.A(n_1366),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1182),
.B(n_957),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1369),
.B(n_1019),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1350),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1183),
.Y(n_1780)
);

BUFx2_ASAP7_75t_L g1781 ( 
.A(n_1314),
.Y(n_1781)
);

BUFx8_ASAP7_75t_SL g1782 ( 
.A(n_1224),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1369),
.B(n_958),
.Y(n_1783)
);

BUFx12f_ASAP7_75t_L g1784 ( 
.A(n_1178),
.Y(n_1784)
);

INVx5_ASAP7_75t_L g1785 ( 
.A(n_1366),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1323),
.B(n_795),
.Y(n_1786)
);

INVx5_ASAP7_75t_L g1787 ( 
.A(n_1366),
.Y(n_1787)
);

INVxp67_ASAP7_75t_L g1788 ( 
.A(n_1351),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1314),
.Y(n_1789)
);

INVx3_ASAP7_75t_L g1790 ( 
.A(n_1423),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1424),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1184),
.B(n_972),
.Y(n_1792)
);

INVx5_ASAP7_75t_L g1793 ( 
.A(n_1366),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1317),
.B(n_985),
.Y(n_1794)
);

INVx5_ASAP7_75t_L g1795 ( 
.A(n_1366),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1352),
.B(n_879),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1353),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1355),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1185),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1425),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1188),
.Y(n_1801)
);

NOR2x1_ASAP7_75t_L g1802 ( 
.A(n_1404),
.B(n_879),
.Y(n_1802)
);

BUFx8_ASAP7_75t_SL g1803 ( 
.A(n_1227),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1426),
.Y(n_1804)
);

BUFx6f_ASAP7_75t_L g1805 ( 
.A(n_1427),
.Y(n_1805)
);

BUFx3_ASAP7_75t_L g1806 ( 
.A(n_1356),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1317),
.B(n_998),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1328),
.B(n_1336),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1429),
.Y(n_1809)
);

BUFx2_ASAP7_75t_L g1810 ( 
.A(n_1328),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1382),
.B(n_1384),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1189),
.B(n_1004),
.Y(n_1812)
);

BUFx12f_ASAP7_75t_L g1813 ( 
.A(n_1336),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1190),
.B(n_1018),
.Y(n_1814)
);

INVx3_ASAP7_75t_L g1815 ( 
.A(n_1433),
.Y(n_1815)
);

INVx4_ASAP7_75t_L g1816 ( 
.A(n_1359),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1191),
.B(n_1036),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1437),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1359),
.B(n_1052),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1377),
.B(n_1379),
.Y(n_1820)
);

INVx5_ASAP7_75t_L g1821 ( 
.A(n_1366),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1192),
.B(n_1047),
.Y(n_1822)
);

BUFx6f_ASAP7_75t_L g1823 ( 
.A(n_1438),
.Y(n_1823)
);

INVx5_ASAP7_75t_L g1824 ( 
.A(n_1329),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1435),
.B(n_1463),
.Y(n_1825)
);

BUFx6f_ASAP7_75t_L g1826 ( 
.A(n_1441),
.Y(n_1826)
);

BUFx12f_ASAP7_75t_L g1827 ( 
.A(n_1377),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1357),
.B(n_930),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_L g1829 ( 
.A(n_1382),
.B(n_1583),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1358),
.B(n_930),
.Y(n_1830)
);

BUFx3_ASAP7_75t_L g1831 ( 
.A(n_1363),
.Y(n_1831)
);

BUFx6f_ASAP7_75t_L g1832 ( 
.A(n_1442),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1195),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_L g1834 ( 
.A(n_1446),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1197),
.Y(n_1835)
);

INVx5_ASAP7_75t_L g1836 ( 
.A(n_1520),
.Y(n_1836)
);

AND2x4_ASAP7_75t_L g1837 ( 
.A(n_1364),
.B(n_930),
.Y(n_1837)
);

INVx6_ASAP7_75t_L g1838 ( 
.A(n_1529),
.Y(n_1838)
);

INVx5_ASAP7_75t_L g1839 ( 
.A(n_1538),
.Y(n_1839)
);

BUFx8_ASAP7_75t_SL g1840 ( 
.A(n_1227),
.Y(n_1840)
);

AND2x4_ASAP7_75t_L g1841 ( 
.A(n_1365),
.B(n_1010),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1373),
.Y(n_1842)
);

BUFx12f_ASAP7_75t_L g1843 ( 
.A(n_1379),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1198),
.B(n_1061),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1447),
.Y(n_1845)
);

BUFx12f_ASAP7_75t_L g1846 ( 
.A(n_1391),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1374),
.Y(n_1847)
);

BUFx6f_ASAP7_75t_L g1848 ( 
.A(n_1448),
.Y(n_1848)
);

BUFx12f_ASAP7_75t_L g1849 ( 
.A(n_1391),
.Y(n_1849)
);

AND2x4_ASAP7_75t_L g1850 ( 
.A(n_1376),
.B(n_1010),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1199),
.B(n_1079),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1380),
.B(n_1010),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1383),
.Y(n_1853)
);

INVx3_ASAP7_75t_L g1854 ( 
.A(n_1451),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1200),
.B(n_1083),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1411),
.B(n_1101),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1411),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1412),
.B(n_1102),
.Y(n_1858)
);

BUFx3_ASAP7_75t_L g1859 ( 
.A(n_1385),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1386),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_L g1861 ( 
.A(n_1453),
.Y(n_1861)
);

INVx5_ASAP7_75t_L g1862 ( 
.A(n_1543),
.Y(n_1862)
);

INVx3_ASAP7_75t_L g1863 ( 
.A(n_1454),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_L g1864 ( 
.A(n_1456),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1384),
.B(n_1387),
.Y(n_1865)
);

BUFx3_ASAP7_75t_L g1866 ( 
.A(n_1388),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1201),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_SL g1868 ( 
.A(n_1565),
.B(n_797),
.Y(n_1868)
);

INVx4_ASAP7_75t_L g1869 ( 
.A(n_1412),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1392),
.Y(n_1870)
);

AND2x6_ASAP7_75t_L g1871 ( 
.A(n_1202),
.B(n_1031),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1206),
.B(n_1133),
.Y(n_1872)
);

BUFx6f_ASAP7_75t_L g1873 ( 
.A(n_1458),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1387),
.B(n_799),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1207),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1208),
.B(n_1031),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1209),
.Y(n_1877)
);

INVx5_ASAP7_75t_L g1878 ( 
.A(n_1212),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1431),
.B(n_1468),
.Y(n_1879)
);

AND2x6_ASAP7_75t_L g1880 ( 
.A(n_1211),
.B(n_1031),
.Y(n_1880)
);

INVx4_ASAP7_75t_L g1881 ( 
.A(n_1452),
.Y(n_1881)
);

BUFx6f_ASAP7_75t_L g1882 ( 
.A(n_1459),
.Y(n_1882)
);

INVx5_ASAP7_75t_L g1883 ( 
.A(n_1214),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1431),
.B(n_801),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1396),
.Y(n_1885)
);

INVx4_ASAP7_75t_L g1886 ( 
.A(n_1452),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1468),
.B(n_805),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1397),
.B(n_1162),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1460),
.Y(n_1889)
);

INVx5_ASAP7_75t_L g1890 ( 
.A(n_1217),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1399),
.B(n_1162),
.Y(n_1891)
);

BUFx6f_ASAP7_75t_L g1892 ( 
.A(n_1461),
.Y(n_1892)
);

INVx6_ASAP7_75t_L g1893 ( 
.A(n_1550),
.Y(n_1893)
);

BUFx12f_ASAP7_75t_L g1894 ( 
.A(n_1457),
.Y(n_1894)
);

NAND2xp33_ASAP7_75t_L g1895 ( 
.A(n_1457),
.B(n_1153),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1401),
.B(n_1162),
.Y(n_1896)
);

BUFx6f_ASAP7_75t_L g1897 ( 
.A(n_1462),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1402),
.B(n_1110),
.Y(n_1898)
);

BUFx12f_ASAP7_75t_L g1899 ( 
.A(n_1465),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1465),
.B(n_806),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1511),
.B(n_808),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1511),
.B(n_813),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1375),
.B(n_1110),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1218),
.Y(n_1904)
);

INVx3_ASAP7_75t_L g1905 ( 
.A(n_1464),
.Y(n_1905)
);

INVx5_ASAP7_75t_L g1906 ( 
.A(n_1220),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1221),
.B(n_1110),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1400),
.B(n_1325),
.Y(n_1908)
);

BUFx6f_ASAP7_75t_L g1909 ( 
.A(n_1467),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1466),
.B(n_1491),
.Y(n_1910)
);

BUFx3_ASAP7_75t_L g1911 ( 
.A(n_1222),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1513),
.B(n_815),
.Y(n_1912)
);

BUFx6f_ASAP7_75t_L g1913 ( 
.A(n_1471),
.Y(n_1913)
);

HB1xp67_ASAP7_75t_L g1914 ( 
.A(n_1466),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1513),
.B(n_816),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1335),
.B(n_691),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1223),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1779),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1798),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1615),
.B(n_1618),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1842),
.Y(n_1921)
);

BUFx6f_ASAP7_75t_L g1922 ( 
.A(n_1588),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1683),
.B(n_1500),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1615),
.B(n_1225),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1586),
.Y(n_1925)
);

BUFx6f_ASAP7_75t_L g1926 ( 
.A(n_1588),
.Y(n_1926)
);

BUFx6f_ASAP7_75t_L g1927 ( 
.A(n_1588),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1737),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1634),
.B(n_1491),
.Y(n_1929)
);

HB1xp67_ASAP7_75t_L g1930 ( 
.A(n_1586),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_L g1931 ( 
.A(n_1606),
.B(n_1519),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1847),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1737),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1853),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1860),
.Y(n_1935)
);

INVx3_ASAP7_75t_L g1936 ( 
.A(n_1591),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1610),
.Y(n_1937)
);

HB1xp67_ASAP7_75t_L g1938 ( 
.A(n_1623),
.Y(n_1938)
);

BUFx2_ASAP7_75t_L g1939 ( 
.A(n_1589),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1870),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1885),
.Y(n_1941)
);

INVx3_ASAP7_75t_L g1942 ( 
.A(n_1591),
.Y(n_1942)
);

BUFx6f_ASAP7_75t_L g1943 ( 
.A(n_1591),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1618),
.B(n_1229),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1917),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1622),
.B(n_1234),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1683),
.B(n_1238),
.Y(n_1947)
);

BUFx6f_ASAP7_75t_L g1948 ( 
.A(n_1592),
.Y(n_1948)
);

BUFx2_ASAP7_75t_L g1949 ( 
.A(n_1614),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1904),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1699),
.Y(n_1951)
);

INVx5_ASAP7_75t_L g1952 ( 
.A(n_1638),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1666),
.B(n_1240),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1737),
.Y(n_1954)
);

INVx1_ASAP7_75t_SL g1955 ( 
.A(n_1782),
.Y(n_1955)
);

HB1xp67_ASAP7_75t_L g1956 ( 
.A(n_1644),
.Y(n_1956)
);

HB1xp67_ASAP7_75t_L g1957 ( 
.A(n_1644),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1648),
.B(n_1500),
.Y(n_1958)
);

BUFx6f_ASAP7_75t_L g1959 ( 
.A(n_1592),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1648),
.B(n_1558),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1738),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1700),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1622),
.B(n_1241),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1738),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1712),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1738),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1745),
.Y(n_1967)
);

HB1xp67_ASAP7_75t_L g1968 ( 
.A(n_1673),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1740),
.Y(n_1969)
);

BUFx6f_ASAP7_75t_L g1970 ( 
.A(n_1592),
.Y(n_1970)
);

INVx4_ASAP7_75t_L g1971 ( 
.A(n_1740),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1652),
.B(n_1558),
.Y(n_1972)
);

INVx3_ASAP7_75t_L g1973 ( 
.A(n_1603),
.Y(n_1973)
);

HB1xp67_ASAP7_75t_L g1974 ( 
.A(n_1673),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1797),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1632),
.B(n_1242),
.Y(n_1976)
);

BUFx2_ASAP7_75t_L g1977 ( 
.A(n_1634),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1740),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1806),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1760),
.Y(n_1980)
);

AND2x4_ASAP7_75t_L g1981 ( 
.A(n_1743),
.B(n_1243),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1831),
.Y(n_1982)
);

INVx3_ASAP7_75t_L g1983 ( 
.A(n_1603),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1652),
.B(n_1561),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1632),
.B(n_1245),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1760),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1611),
.B(n_1246),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1859),
.Y(n_1988)
);

HB1xp67_ASAP7_75t_L g1989 ( 
.A(n_1682),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1630),
.B(n_1248),
.Y(n_1990)
);

BUFx6f_ASAP7_75t_L g1991 ( 
.A(n_1603),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1866),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1911),
.Y(n_1993)
);

HB1xp67_ASAP7_75t_L g1994 ( 
.A(n_1682),
.Y(n_1994)
);

XNOR2xp5_ASAP7_75t_L g1995 ( 
.A(n_1719),
.B(n_1232),
.Y(n_1995)
);

INVx3_ASAP7_75t_L g1996 ( 
.A(n_1609),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1761),
.Y(n_1997)
);

INVx3_ASAP7_75t_L g1998 ( 
.A(n_1609),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1780),
.Y(n_1999)
);

AND2x4_ASAP7_75t_L g2000 ( 
.A(n_1743),
.B(n_1252),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1799),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1760),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1801),
.Y(n_2003)
);

INVxp67_ASAP7_75t_L g2004 ( 
.A(n_1874),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1763),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_1772),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1833),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1835),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1867),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1875),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1763),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1877),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1763),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1769),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1769),
.Y(n_2015)
);

INVxp67_ASAP7_75t_SL g2016 ( 
.A(n_1609),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_1748),
.B(n_1254),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1748),
.Y(n_2018)
);

AND2x4_ASAP7_75t_L g2019 ( 
.A(n_1661),
.B(n_1256),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1769),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1631),
.Y(n_2021)
);

INVx3_ASAP7_75t_L g2022 ( 
.A(n_1628),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1585),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1620),
.B(n_1257),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1645),
.Y(n_2025)
);

BUFx6f_ASAP7_75t_L g2026 ( 
.A(n_1628),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1593),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1678),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1595),
.Y(n_2029)
);

INVx3_ASAP7_75t_L g2030 ( 
.A(n_1628),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1689),
.Y(n_2031)
);

BUFx6f_ASAP7_75t_L g2032 ( 
.A(n_1637),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1661),
.B(n_1561),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1665),
.B(n_1562),
.Y(n_2034)
);

BUFx6f_ASAP7_75t_L g2035 ( 
.A(n_1637),
.Y(n_2035)
);

BUFx6f_ASAP7_75t_L g2036 ( 
.A(n_1637),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1633),
.B(n_1519),
.Y(n_2037)
);

BUFx8_ASAP7_75t_L g2038 ( 
.A(n_1619),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1803),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1620),
.B(n_1258),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1696),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_1633),
.B(n_1515),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1596),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1709),
.Y(n_2044)
);

INVxp67_ASAP7_75t_L g2045 ( 
.A(n_1874),
.Y(n_2045)
);

AND2x4_ASAP7_75t_L g2046 ( 
.A(n_1665),
.B(n_1259),
.Y(n_2046)
);

BUFx8_ASAP7_75t_L g2047 ( 
.A(n_1658),
.Y(n_2047)
);

AND2x4_ASAP7_75t_L g2048 ( 
.A(n_1749),
.B(n_1260),
.Y(n_2048)
);

NAND2xp33_ASAP7_75t_L g2049 ( 
.A(n_1871),
.B(n_863),
.Y(n_2049)
);

BUFx6f_ASAP7_75t_L g2050 ( 
.A(n_1650),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1775),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1775),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_L g2053 ( 
.A(n_1650),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1629),
.B(n_1515),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1599),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1626),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1662),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1775),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1650),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1791),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1791),
.Y(n_2061)
);

OAI22xp5_ASAP7_75t_SL g2062 ( 
.A1(n_1624),
.A2(n_1232),
.B1(n_1284),
.B2(n_1244),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1667),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1765),
.B(n_1770),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1791),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1730),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1750),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1739),
.Y(n_2068)
);

INVx3_ASAP7_75t_L g2069 ( 
.A(n_1651),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1765),
.B(n_1770),
.Y(n_2070)
);

BUFx6f_ASAP7_75t_L g2071 ( 
.A(n_1651),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1746),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1752),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1757),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1651),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1800),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1800),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1800),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1653),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1903),
.B(n_1698),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1777),
.B(n_1277),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1804),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_1653),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1653),
.Y(n_2084)
);

OR2x2_ASAP7_75t_L g2085 ( 
.A(n_1772),
.B(n_1315),
.Y(n_2085)
);

BUFx6f_ASAP7_75t_L g2086 ( 
.A(n_1655),
.Y(n_2086)
);

BUFx6f_ASAP7_75t_L g2087 ( 
.A(n_1655),
.Y(n_2087)
);

AND2x6_ASAP7_75t_L g2088 ( 
.A(n_1621),
.B(n_691),
.Y(n_2088)
);

CKINVDCx11_ASAP7_75t_R g2089 ( 
.A(n_1605),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1804),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1655),
.Y(n_2091)
);

INVx3_ASAP7_75t_L g2092 ( 
.A(n_1669),
.Y(n_2092)
);

BUFx6f_ASAP7_75t_L g2093 ( 
.A(n_1669),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1669),
.Y(n_2094)
);

BUFx6f_ASAP7_75t_L g2095 ( 
.A(n_1680),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1680),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1804),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1805),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1680),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1805),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1805),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1823),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1823),
.Y(n_2103)
);

BUFx6f_ASAP7_75t_L g2104 ( 
.A(n_1681),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1823),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1681),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1681),
.Y(n_2107)
);

BUFx6f_ASAP7_75t_L g2108 ( 
.A(n_1686),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_L g2109 ( 
.A(n_1686),
.Y(n_2109)
);

BUFx6f_ASAP7_75t_L g2110 ( 
.A(n_1686),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1616),
.Y(n_2111)
);

CKINVDCx16_ASAP7_75t_R g2112 ( 
.A(n_1613),
.Y(n_2112)
);

INVxp67_ASAP7_75t_L g2113 ( 
.A(n_1884),
.Y(n_2113)
);

HB1xp67_ASAP7_75t_L g2114 ( 
.A(n_1694),
.Y(n_2114)
);

INVxp67_ASAP7_75t_L g2115 ( 
.A(n_1884),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_1777),
.B(n_1280),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_1903),
.B(n_1562),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1698),
.B(n_1576),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1826),
.Y(n_2119)
);

BUFx8_ASAP7_75t_L g2120 ( 
.A(n_1771),
.Y(n_2120)
);

BUFx6f_ASAP7_75t_L g2121 ( 
.A(n_1826),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1616),
.Y(n_2122)
);

AND2x4_ASAP7_75t_L g2123 ( 
.A(n_1749),
.B(n_1282),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1826),
.Y(n_2124)
);

BUFx6f_ASAP7_75t_L g2125 ( 
.A(n_1832),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1832),
.Y(n_2126)
);

BUFx6f_ASAP7_75t_L g2127 ( 
.A(n_1832),
.Y(n_2127)
);

BUFx2_ASAP7_75t_L g2128 ( 
.A(n_1695),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1834),
.Y(n_2129)
);

XNOR2x2_ASAP7_75t_R g2130 ( 
.A(n_1646),
.B(n_777),
.Y(n_2130)
);

INVx5_ASAP7_75t_L g2131 ( 
.A(n_1638),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1671),
.Y(n_2132)
);

INVx3_ASAP7_75t_L g2133 ( 
.A(n_1590),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1671),
.Y(n_2134)
);

HB1xp67_ASAP7_75t_L g2135 ( 
.A(n_1735),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1834),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1834),
.Y(n_2137)
);

CKINVDCx5p33_ASAP7_75t_R g2138 ( 
.A(n_1840),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1845),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1715),
.Y(n_2140)
);

BUFx6f_ASAP7_75t_L g2141 ( 
.A(n_1845),
.Y(n_2141)
);

OA21x2_ASAP7_75t_L g2142 ( 
.A1(n_1876),
.A2(n_1406),
.B(n_1405),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1715),
.Y(n_2143)
);

INVx3_ASAP7_75t_L g2144 ( 
.A(n_1590),
.Y(n_2144)
);

BUFx3_ASAP7_75t_L g2145 ( 
.A(n_1602),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1792),
.B(n_1286),
.Y(n_2146)
);

BUFx3_ASAP7_75t_L g2147 ( 
.A(n_1602),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_SL g2148 ( 
.A(n_1624),
.B(n_1542),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_1753),
.B(n_1289),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_1889),
.Y(n_2150)
);

INVx3_ASAP7_75t_L g2151 ( 
.A(n_1590),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1845),
.Y(n_2152)
);

BUFx6f_ASAP7_75t_L g2153 ( 
.A(n_1848),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1792),
.B(n_1292),
.Y(n_2154)
);

BUFx6f_ASAP7_75t_L g2155 ( 
.A(n_1848),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1848),
.Y(n_2156)
);

BUFx6f_ASAP7_75t_L g2157 ( 
.A(n_1861),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_1788),
.B(n_1908),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1861),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1861),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_1753),
.B(n_1295),
.Y(n_2161)
);

OR2x6_ASAP7_75t_L g2162 ( 
.A(n_1813),
.B(n_1550),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_1812),
.B(n_1296),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_1812),
.B(n_1297),
.Y(n_2164)
);

NOR2xp33_ASAP7_75t_L g2165 ( 
.A(n_1635),
.B(n_1542),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1864),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1814),
.B(n_1299),
.Y(n_2167)
);

INVx3_ASAP7_75t_L g2168 ( 
.A(n_1590),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1876),
.Y(n_2169)
);

NAND2x1_ASAP7_75t_L g2170 ( 
.A(n_1638),
.B(n_1408),
.Y(n_2170)
);

XNOR2xp5_ASAP7_75t_L g2171 ( 
.A(n_1825),
.B(n_1244),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1864),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1864),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1873),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1873),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1873),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1882),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1882),
.Y(n_2178)
);

AND3x1_ASAP7_75t_L g2179 ( 
.A(n_1613),
.B(n_961),
.C(n_956),
.Y(n_2179)
);

BUFx6f_ASAP7_75t_L g2180 ( 
.A(n_1882),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1892),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1892),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1892),
.Y(n_2183)
);

HB1xp67_ASAP7_75t_L g2184 ( 
.A(n_1735),
.Y(n_2184)
);

INVx3_ASAP7_75t_L g2185 ( 
.A(n_1597),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1897),
.Y(n_2186)
);

BUFx6f_ASAP7_75t_L g2187 ( 
.A(n_1897),
.Y(n_2187)
);

HB1xp67_ASAP7_75t_L g2188 ( 
.A(n_1754),
.Y(n_2188)
);

BUFx6f_ASAP7_75t_L g2189 ( 
.A(n_1897),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1909),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1909),
.Y(n_2191)
);

BUFx3_ASAP7_75t_L g2192 ( 
.A(n_1607),
.Y(n_2192)
);

AND2x4_ASAP7_75t_L g2193 ( 
.A(n_1758),
.B(n_1300),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_1788),
.B(n_1576),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1909),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1814),
.B(n_1301),
.Y(n_2196)
);

BUFx6f_ASAP7_75t_L g2197 ( 
.A(n_1913),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_1817),
.B(n_1306),
.Y(n_2198)
);

CKINVDCx5p33_ASAP7_75t_R g2199 ( 
.A(n_1641),
.Y(n_2199)
);

BUFx3_ASAP7_75t_L g2200 ( 
.A(n_1607),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1913),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1913),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1790),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1790),
.Y(n_2204)
);

OAI22xp5_ASAP7_75t_SL g2205 ( 
.A1(n_1901),
.A2(n_1290),
.B1(n_1368),
.B2(n_1284),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_SL g2206 ( 
.A(n_1824),
.B(n_1546),
.Y(n_2206)
);

AND2x4_ASAP7_75t_L g2207 ( 
.A(n_1758),
.B(n_1307),
.Y(n_2207)
);

CKINVDCx6p67_ASAP7_75t_R g2208 ( 
.A(n_1824),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1817),
.B(n_1313),
.Y(n_2209)
);

BUFx6f_ASAP7_75t_L g2210 ( 
.A(n_1597),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1822),
.B(n_1316),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1822),
.B(n_1319),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1809),
.Y(n_2213)
);

BUFx6f_ASAP7_75t_L g2214 ( 
.A(n_1597),
.Y(n_2214)
);

BUFx2_ASAP7_75t_L g2215 ( 
.A(n_1598),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_1768),
.B(n_1320),
.Y(n_2216)
);

AND2x2_ASAP7_75t_SL g2217 ( 
.A(n_1647),
.B(n_941),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1809),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_1908),
.B(n_1584),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1815),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1815),
.Y(n_2221)
);

BUFx8_ASAP7_75t_L g2222 ( 
.A(n_1784),
.Y(n_2222)
);

HB1xp67_ASAP7_75t_L g2223 ( 
.A(n_1754),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1818),
.Y(n_2224)
);

HB1xp67_ASAP7_75t_L g2225 ( 
.A(n_1755),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_1818),
.Y(n_2226)
);

HB1xp67_ASAP7_75t_L g2227 ( 
.A(n_1755),
.Y(n_2227)
);

HB1xp67_ASAP7_75t_L g2228 ( 
.A(n_1764),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1844),
.B(n_1321),
.Y(n_2229)
);

BUFx6f_ASAP7_75t_L g2230 ( 
.A(n_1597),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1854),
.Y(n_2231)
);

OAI22xp5_ASAP7_75t_SL g2232 ( 
.A1(n_1901),
.A2(n_1368),
.B1(n_1372),
.B2(n_1290),
.Y(n_2232)
);

INVx3_ASAP7_75t_L g2233 ( 
.A(n_1717),
.Y(n_2233)
);

AND2x4_ASAP7_75t_L g2234 ( 
.A(n_1768),
.B(n_1322),
.Y(n_2234)
);

INVx2_ASAP7_75t_SL g2235 ( 
.A(n_1893),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1854),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1863),
.Y(n_2237)
);

BUFx6f_ASAP7_75t_L g2238 ( 
.A(n_1796),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1863),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1905),
.Y(n_2240)
);

INVx3_ASAP7_75t_L g2241 ( 
.A(n_1717),
.Y(n_2241)
);

INVx3_ASAP7_75t_L g2242 ( 
.A(n_1717),
.Y(n_2242)
);

NOR2xp33_ASAP7_75t_L g2243 ( 
.A(n_1635),
.B(n_1546),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_1905),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1796),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1828),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1828),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1717),
.Y(n_2248)
);

HB1xp67_ASAP7_75t_L g2249 ( 
.A(n_1764),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1830),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1830),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_SL g2252 ( 
.A(n_1824),
.B(n_1553),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1837),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1725),
.Y(n_2254)
);

BUFx3_ASAP7_75t_L g2255 ( 
.A(n_1871),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1837),
.Y(n_2256)
);

AND2x4_ASAP7_75t_L g2257 ( 
.A(n_1841),
.B(n_1324),
.Y(n_2257)
);

BUFx8_ASAP7_75t_L g2258 ( 
.A(n_1734),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1725),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1841),
.Y(n_2260)
);

CKINVDCx5p33_ASAP7_75t_R g2261 ( 
.A(n_1641),
.Y(n_2261)
);

INVx3_ASAP7_75t_L g2262 ( 
.A(n_1725),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_1824),
.B(n_1553),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_1640),
.A2(n_1203),
.B1(n_1236),
.B2(n_1554),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1725),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_1726),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1726),
.Y(n_2267)
);

INVx3_ASAP7_75t_L g2268 ( 
.A(n_1726),
.Y(n_2268)
);

OAI22xp5_ASAP7_75t_L g2269 ( 
.A1(n_1893),
.A2(n_1203),
.B1(n_1236),
.B2(n_1233),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_1844),
.B(n_1327),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1850),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1850),
.Y(n_2272)
);

NOR2xp33_ASAP7_75t_SL g2273 ( 
.A(n_1836),
.B(n_1378),
.Y(n_2273)
);

AND2x4_ASAP7_75t_L g2274 ( 
.A(n_1852),
.B(n_1584),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_1726),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1852),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1802),
.Y(n_2277)
);

HB1xp67_ASAP7_75t_L g2278 ( 
.A(n_1900),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_1851),
.B(n_1554),
.Y(n_2279)
);

CKINVDCx5p33_ASAP7_75t_R g2280 ( 
.A(n_1649),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1888),
.Y(n_2281)
);

BUFx3_ASAP7_75t_L g2282 ( 
.A(n_1871),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1888),
.Y(n_2283)
);

INVxp67_ASAP7_75t_L g2284 ( 
.A(n_1902),
.Y(n_2284)
);

INVx3_ASAP7_75t_L g2285 ( 
.A(n_1759),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1891),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1891),
.Y(n_2287)
);

INVx3_ASAP7_75t_L g2288 ( 
.A(n_1759),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_1604),
.B(n_1326),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_1759),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_1759),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_1604),
.B(n_1326),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_1762),
.Y(n_2293)
);

AOI22x1_ASAP7_75t_SL g2294 ( 
.A1(n_1684),
.A2(n_1393),
.B1(n_1394),
.B2(n_1372),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1896),
.Y(n_2295)
);

INVx3_ASAP7_75t_L g2296 ( 
.A(n_1762),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1896),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1898),
.Y(n_2298)
);

OR2x6_ASAP7_75t_L g2299 ( 
.A(n_1827),
.B(n_1362),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_1871),
.Y(n_2300)
);

OR2x2_ASAP7_75t_L g2301 ( 
.A(n_2085),
.B(n_1449),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_2111),
.Y(n_2302)
);

CKINVDCx6p67_ASAP7_75t_R g2303 ( 
.A(n_2089),
.Y(n_2303)
);

BUFx6f_ASAP7_75t_L g2304 ( 
.A(n_2300),
.Y(n_2304)
);

NAND2xp33_ASAP7_75t_L g2305 ( 
.A(n_2064),
.B(n_863),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2111),
.Y(n_2306)
);

NOR2xp33_ASAP7_75t_L g2307 ( 
.A(n_2004),
.B(n_1670),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2122),
.Y(n_2308)
);

AOI22xp33_ASAP7_75t_L g2309 ( 
.A1(n_2169),
.A2(n_1893),
.B1(n_1687),
.B2(n_1691),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2122),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2132),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_SL g2312 ( 
.A(n_2037),
.B(n_1836),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2132),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_1920),
.B(n_1851),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2134),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_SL g2316 ( 
.A(n_2037),
.B(n_1836),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2070),
.B(n_2169),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1958),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1958),
.Y(n_2319)
);

HB1xp67_ASAP7_75t_L g2320 ( 
.A(n_1925),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_2042),
.B(n_1836),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2281),
.B(n_2283),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_SL g2323 ( 
.A(n_2042),
.B(n_2165),
.Y(n_2323)
);

BUFx6f_ASAP7_75t_L g2324 ( 
.A(n_2300),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2134),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2142),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2142),
.Y(n_2327)
);

NOR2x1p5_ASAP7_75t_L g2328 ( 
.A(n_2208),
.B(n_1843),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1960),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_SL g2330 ( 
.A(n_2165),
.B(n_1839),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2286),
.B(n_1687),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2287),
.B(n_1691),
.Y(n_2332)
);

INVx4_ASAP7_75t_L g2333 ( 
.A(n_2300),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2142),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_SL g2335 ( 
.A(n_2243),
.B(n_1839),
.Y(n_2335)
);

BUFx10_ASAP7_75t_L g2336 ( 
.A(n_2243),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_1960),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2023),
.Y(n_2338)
);

INVx3_ASAP7_75t_L g2339 ( 
.A(n_2300),
.Y(n_2339)
);

CKINVDCx6p67_ASAP7_75t_R g2340 ( 
.A(n_2089),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2023),
.Y(n_2341)
);

INVx3_ASAP7_75t_L g2342 ( 
.A(n_2300),
.Y(n_2342)
);

NAND2xp33_ASAP7_75t_L g2343 ( 
.A(n_2088),
.B(n_2279),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2027),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_1972),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2027),
.Y(n_2346)
);

NAND3xp33_ASAP7_75t_L g2347 ( 
.A(n_1931),
.B(n_1640),
.C(n_1705),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2029),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_L g2349 ( 
.A(n_2045),
.B(n_2113),
.Y(n_2349)
);

BUFx6f_ASAP7_75t_L g2350 ( 
.A(n_2255),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2295),
.B(n_1677),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2029),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2043),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2043),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_SL g2355 ( 
.A(n_1939),
.B(n_1839),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_1939),
.B(n_1839),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2055),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2297),
.B(n_1855),
.Y(n_2358)
);

INVx1_ASAP7_75t_SL g2359 ( 
.A(n_1930),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2055),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_SL g2361 ( 
.A(n_1949),
.B(n_1862),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2056),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_2298),
.B(n_1677),
.Y(n_2363)
);

INVx2_ASAP7_75t_SL g2364 ( 
.A(n_2080),
.Y(n_2364)
);

INVx3_ASAP7_75t_L g2365 ( 
.A(n_2255),
.Y(n_2365)
);

NAND2xp33_ASAP7_75t_L g2366 ( 
.A(n_2088),
.B(n_863),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2056),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2057),
.Y(n_2368)
);

AOI21x1_ASAP7_75t_L g2369 ( 
.A1(n_2081),
.A2(n_1872),
.B(n_1855),
.Y(n_2369)
);

AO22x2_ASAP7_75t_L g2370 ( 
.A1(n_2115),
.A2(n_1707),
.B1(n_1697),
.B2(n_961),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2057),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_2289),
.B(n_1685),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2063),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2063),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2116),
.B(n_1872),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_SL g2376 ( 
.A(n_1949),
.B(n_1862),
.Y(n_2376)
);

HB1xp67_ASAP7_75t_L g2377 ( 
.A(n_1977),
.Y(n_2377)
);

OR2x2_ASAP7_75t_L g2378 ( 
.A(n_2085),
.B(n_1495),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2146),
.B(n_1636),
.Y(n_2379)
);

INVx8_ASAP7_75t_L g2380 ( 
.A(n_2088),
.Y(n_2380)
);

NOR2xp33_ASAP7_75t_L g2381 ( 
.A(n_2284),
.B(n_1670),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2154),
.B(n_1636),
.Y(n_2382)
);

INVx3_ASAP7_75t_L g2383 ( 
.A(n_2282),
.Y(n_2383)
);

AND2x2_ASAP7_75t_L g2384 ( 
.A(n_2289),
.B(n_1685),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2068),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2068),
.Y(n_2386)
);

BUFx3_ASAP7_75t_L g2387 ( 
.A(n_2145),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2163),
.B(n_1639),
.Y(n_2388)
);

CKINVDCx20_ASAP7_75t_R g2389 ( 
.A(n_1995),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2164),
.B(n_1639),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2218),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2167),
.B(n_1642),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2218),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2226),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_L g2395 ( 
.A(n_2148),
.B(n_1688),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2072),
.Y(n_2396)
);

INVx3_ASAP7_75t_L g2397 ( 
.A(n_2282),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2072),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_SL g2399 ( 
.A(n_2292),
.B(n_2128),
.Y(n_2399)
);

BUFx6f_ASAP7_75t_SL g2400 ( 
.A(n_2217),
.Y(n_2400)
);

NAND2xp33_ASAP7_75t_L g2401 ( 
.A(n_2088),
.B(n_863),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2073),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_SL g2403 ( 
.A(n_2292),
.B(n_1862),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2226),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_SL g2405 ( 
.A(n_2128),
.B(n_1862),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2196),
.B(n_1642),
.Y(n_2406)
);

BUFx4f_ASAP7_75t_L g2407 ( 
.A(n_2088),
.Y(n_2407)
);

AOI22xp33_ASAP7_75t_L g2408 ( 
.A1(n_1947),
.A2(n_1705),
.B1(n_1742),
.B2(n_1721),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2073),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_SL g2410 ( 
.A(n_1977),
.B(n_1688),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_2074),
.Y(n_2411)
);

BUFx6f_ASAP7_75t_L g2412 ( 
.A(n_2238),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2198),
.B(n_2209),
.Y(n_2413)
);

BUFx3_ASAP7_75t_L g2414 ( 
.A(n_2145),
.Y(n_2414)
);

BUFx6f_ASAP7_75t_L g2415 ( 
.A(n_2238),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2074),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2211),
.B(n_1643),
.Y(n_2417)
);

INVx1_ASAP7_75t_SL g2418 ( 
.A(n_2006),
.Y(n_2418)
);

INVx2_ASAP7_75t_SL g2419 ( 
.A(n_2080),
.Y(n_2419)
);

INVxp67_ASAP7_75t_SL g2420 ( 
.A(n_1991),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2066),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_SL g2422 ( 
.A(n_2217),
.B(n_1693),
.Y(n_2422)
);

NOR2x1p5_ASAP7_75t_L g2423 ( 
.A(n_2208),
.B(n_1846),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_1972),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2212),
.B(n_1643),
.Y(n_2425)
);

CKINVDCx6p67_ASAP7_75t_R g2426 ( 
.A(n_1955),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2066),
.Y(n_2427)
);

INVxp67_ASAP7_75t_SL g2428 ( 
.A(n_1991),
.Y(n_2428)
);

INVx3_ASAP7_75t_L g2429 ( 
.A(n_2170),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_L g2430 ( 
.A(n_2148),
.B(n_1693),
.Y(n_2430)
);

INVx1_ASAP7_75t_SL g2431 ( 
.A(n_1956),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2067),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_1984),
.Y(n_2433)
);

XNOR2xp5_ASAP7_75t_L g2434 ( 
.A(n_1995),
.B(n_2171),
.Y(n_2434)
);

INVx1_ASAP7_75t_SL g2435 ( 
.A(n_1957),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2067),
.Y(n_2436)
);

INVx6_ASAP7_75t_L g2437 ( 
.A(n_2238),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_1984),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_SL g2439 ( 
.A(n_2235),
.B(n_1886),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2033),
.Y(n_2440)
);

CKINVDCx20_ASAP7_75t_R g2441 ( 
.A(n_2205),
.Y(n_2441)
);

INVx3_ASAP7_75t_L g2442 ( 
.A(n_2170),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2140),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2033),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2034),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2034),
.Y(n_2446)
);

BUFx3_ASAP7_75t_L g2447 ( 
.A(n_2147),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_1923),
.Y(n_2448)
);

NAND3xp33_ASAP7_75t_L g2449 ( 
.A(n_1931),
.B(n_1742),
.C(n_1721),
.Y(n_2449)
);

INVxp67_ASAP7_75t_SL g2450 ( 
.A(n_1991),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_SL g2451 ( 
.A(n_2235),
.B(n_1816),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_SL g2452 ( 
.A(n_2158),
.B(n_1816),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2158),
.B(n_1869),
.Y(n_2453)
);

BUFx3_ASAP7_75t_L g2454 ( 
.A(n_2147),
.Y(n_2454)
);

NOR2xp33_ASAP7_75t_L g2455 ( 
.A(n_2054),
.B(n_1869),
.Y(n_2455)
);

CKINVDCx5p33_ASAP7_75t_R g2456 ( 
.A(n_2039),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2229),
.B(n_1663),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_2024),
.B(n_2040),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2140),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2143),
.Y(n_2460)
);

AO21x2_ASAP7_75t_L g2461 ( 
.A1(n_2270),
.A2(n_1729),
.B(n_1716),
.Y(n_2461)
);

BUFx10_ASAP7_75t_L g2462 ( 
.A(n_2039),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_1924),
.B(n_1663),
.Y(n_2463)
);

OAI22xp33_ASAP7_75t_L g2464 ( 
.A1(n_1944),
.A2(n_1756),
.B1(n_1727),
.B2(n_1660),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_1923),
.Y(n_2465)
);

BUFx3_ASAP7_75t_L g2466 ( 
.A(n_2192),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2237),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2143),
.Y(n_2468)
);

CKINVDCx6p67_ASAP7_75t_R g2469 ( 
.A(n_2299),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2237),
.Y(n_2470)
);

BUFx6f_ASAP7_75t_L g2471 ( 
.A(n_2238),
.Y(n_2471)
);

NOR2xp33_ASAP7_75t_L g2472 ( 
.A(n_2054),
.B(n_1881),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2244),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2244),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2274),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2274),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_1946),
.B(n_1668),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2274),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2150),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2150),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2203),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_1928),
.Y(n_2482)
);

BUFx10_ASAP7_75t_L g2483 ( 
.A(n_2138),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_1963),
.B(n_1668),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_1928),
.Y(n_2485)
);

INVxp33_ASAP7_75t_L g2486 ( 
.A(n_1968),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2204),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_SL g2488 ( 
.A(n_2114),
.B(n_1881),
.Y(n_2488)
);

INVxp33_ASAP7_75t_L g2489 ( 
.A(n_1974),
.Y(n_2489)
);

NOR2xp33_ASAP7_75t_SL g2490 ( 
.A(n_2199),
.B(n_1849),
.Y(n_2490)
);

NAND3xp33_ASAP7_75t_L g2491 ( 
.A(n_2264),
.B(n_1747),
.C(n_1744),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_1976),
.B(n_1672),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_1933),
.Y(n_2493)
);

NOR2xp33_ASAP7_75t_L g2494 ( 
.A(n_1929),
.B(n_1886),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_SL g2495 ( 
.A(n_1947),
.B(n_1612),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2213),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_1985),
.B(n_1672),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_1933),
.Y(n_2498)
);

BUFx3_ASAP7_75t_L g2499 ( 
.A(n_2192),
.Y(n_2499)
);

OAI22xp33_ASAP7_75t_L g2500 ( 
.A1(n_2273),
.A2(n_1756),
.B1(n_1727),
.B2(n_1660),
.Y(n_2500)
);

AND2x2_ASAP7_75t_L g2501 ( 
.A(n_2219),
.B(n_1724),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_1954),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2220),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2221),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_1954),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_1961),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_1961),
.Y(n_2507)
);

OR2x6_ASAP7_75t_L g2508 ( 
.A(n_2162),
.B(n_1894),
.Y(n_2508)
);

BUFx6f_ASAP7_75t_L g2509 ( 
.A(n_2200),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_1964),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_1964),
.Y(n_2511)
);

AOI21x1_ASAP7_75t_L g2512 ( 
.A1(n_1997),
.A2(n_1729),
.B(n_1716),
.Y(n_2512)
);

NOR2xp33_ASAP7_75t_L g2513 ( 
.A(n_1929),
.B(n_1692),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_1947),
.B(n_1711),
.Y(n_2514)
);

INVx3_ASAP7_75t_L g2515 ( 
.A(n_2075),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_1966),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2021),
.B(n_1676),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_1966),
.Y(n_2518)
);

OAI22xp33_ASAP7_75t_L g2519 ( 
.A1(n_2278),
.A2(n_1647),
.B1(n_1219),
.B2(n_1233),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2224),
.Y(n_2520)
);

AND2x2_ASAP7_75t_SL g2521 ( 
.A(n_2179),
.B(n_1704),
.Y(n_2521)
);

NAND2xp33_ASAP7_75t_L g2522 ( 
.A(n_2088),
.B(n_863),
.Y(n_2522)
);

INVx4_ASAP7_75t_L g2523 ( 
.A(n_2086),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_1969),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_1969),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_1978),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_1978),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_SL g2528 ( 
.A(n_2200),
.B(n_1808),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_1980),
.Y(n_2529)
);

INVx2_ASAP7_75t_SL g2530 ( 
.A(n_1953),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_1999),
.B(n_1676),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_SL g2532 ( 
.A(n_2019),
.B(n_1820),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_1980),
.Y(n_2533)
);

INVx2_ASAP7_75t_SL g2534 ( 
.A(n_1953),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_1986),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_1986),
.Y(n_2536)
);

BUFx6f_ASAP7_75t_L g2537 ( 
.A(n_2086),
.Y(n_2537)
);

INVx3_ASAP7_75t_L g2538 ( 
.A(n_2075),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2002),
.Y(n_2539)
);

INVx2_ASAP7_75t_SL g2540 ( 
.A(n_1953),
.Y(n_2540)
);

INVx8_ASAP7_75t_L g2541 ( 
.A(n_2019),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2002),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2001),
.B(n_1783),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2005),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2231),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2005),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2236),
.Y(n_2547)
);

INVx2_ASAP7_75t_SL g2548 ( 
.A(n_2117),
.Y(n_2548)
);

INVxp67_ASAP7_75t_L g2549 ( 
.A(n_1989),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2003),
.B(n_1731),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2011),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2007),
.B(n_1731),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_1945),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_1950),
.Y(n_2554)
);

BUFx2_ASAP7_75t_L g2555 ( 
.A(n_1994),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_1918),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_1919),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_SL g2558 ( 
.A(n_2019),
.B(n_1910),
.Y(n_2558)
);

INVx2_ASAP7_75t_SL g2559 ( 
.A(n_2117),
.Y(n_2559)
);

INVx3_ASAP7_75t_L g2560 ( 
.A(n_2079),
.Y(n_2560)
);

NOR2xp33_ASAP7_75t_L g2561 ( 
.A(n_2269),
.B(n_1887),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_SL g2562 ( 
.A(n_2046),
.B(n_1704),
.Y(n_2562)
);

INVx2_ASAP7_75t_SL g2563 ( 
.A(n_2219),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_1921),
.Y(n_2564)
);

NOR2xp33_ASAP7_75t_L g2565 ( 
.A(n_2206),
.B(n_1902),
.Y(n_2565)
);

AOI22xp5_ASAP7_75t_L g2566 ( 
.A1(n_2118),
.A2(n_1829),
.B1(n_1865),
.B2(n_1811),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2011),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2013),
.Y(n_2568)
);

AND3x2_ASAP7_75t_L g2569 ( 
.A(n_2215),
.B(n_1608),
.C(n_1594),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2008),
.B(n_1732),
.Y(n_2570)
);

INVx3_ASAP7_75t_L g2571 ( 
.A(n_2079),
.Y(n_2571)
);

BUFx2_ASAP7_75t_L g2572 ( 
.A(n_2135),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_1932),
.Y(n_2573)
);

CKINVDCx6p67_ASAP7_75t_R g2574 ( 
.A(n_2299),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_2013),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_1934),
.Y(n_2576)
);

INVx4_ASAP7_75t_L g2577 ( 
.A(n_2086),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_1935),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2014),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2009),
.B(n_1732),
.Y(n_2580)
);

AND2x2_ASAP7_75t_L g2581 ( 
.A(n_2118),
.B(n_1724),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_SL g2582 ( 
.A(n_2046),
.B(n_1811),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2014),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_2015),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_1940),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2015),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2020),
.Y(n_2587)
);

AOI22xp33_ASAP7_75t_L g2588 ( 
.A1(n_2046),
.A2(n_1744),
.B1(n_1778),
.B2(n_1747),
.Y(n_2588)
);

INVx4_ASAP7_75t_L g2589 ( 
.A(n_2086),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2020),
.Y(n_2590)
);

NOR2xp33_ASAP7_75t_L g2591 ( 
.A(n_2206),
.B(n_1912),
.Y(n_2591)
);

INVx4_ASAP7_75t_L g2592 ( 
.A(n_2086),
.Y(n_2592)
);

NOR2xp33_ASAP7_75t_L g2593 ( 
.A(n_2252),
.B(n_1912),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_1941),
.Y(n_2594)
);

AOI22xp5_ASAP7_75t_L g2595 ( 
.A1(n_2018),
.A2(n_1865),
.B1(n_1879),
.B2(n_1829),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2239),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2010),
.B(n_1733),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2012),
.B(n_1733),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2240),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2025),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2083),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2028),
.Y(n_2602)
);

NAND3xp33_ASAP7_75t_L g2603 ( 
.A(n_2245),
.B(n_1778),
.C(n_1895),
.Y(n_2603)
);

INVx3_ASAP7_75t_L g2604 ( 
.A(n_2083),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2084),
.Y(n_2605)
);

INVx2_ASAP7_75t_SL g2606 ( 
.A(n_1981),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2084),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_SL g2608 ( 
.A(n_1981),
.B(n_1879),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2031),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2041),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2091),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2091),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2094),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2044),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2246),
.Y(n_2615)
);

INVx2_ASAP7_75t_SL g2616 ( 
.A(n_1981),
.Y(n_2616)
);

AOI22xp33_ASAP7_75t_L g2617 ( 
.A1(n_2048),
.A2(n_1871),
.B1(n_1880),
.B2(n_1915),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2247),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2250),
.Y(n_2619)
);

AOI22xp33_ASAP7_75t_L g2620 ( 
.A1(n_2048),
.A2(n_2149),
.B1(n_2161),
.B2(n_2123),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2251),
.Y(n_2621)
);

BUFx6f_ASAP7_75t_L g2622 ( 
.A(n_2087),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2253),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2256),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2094),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2260),
.Y(n_2626)
);

INVx2_ASAP7_75t_SL g2627 ( 
.A(n_2000),
.Y(n_2627)
);

INVx2_ASAP7_75t_SL g2628 ( 
.A(n_2000),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2096),
.Y(n_2629)
);

INVx4_ASAP7_75t_L g2630 ( 
.A(n_2087),
.Y(n_2630)
);

OR2x6_ASAP7_75t_L g2631 ( 
.A(n_2162),
.B(n_1899),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2271),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2272),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_SL g2634 ( 
.A(n_2000),
.B(n_1649),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2277),
.B(n_1741),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_SL g2636 ( 
.A(n_2017),
.B(n_1794),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2276),
.Y(n_2637)
);

INVx3_ASAP7_75t_L g2638 ( 
.A(n_2096),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2099),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2099),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_SL g2641 ( 
.A(n_2017),
.B(n_1807),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2106),
.Y(n_2642)
);

BUFx6f_ASAP7_75t_L g2643 ( 
.A(n_2087),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2106),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2107),
.Y(n_2645)
);

AOI22xp33_ASAP7_75t_L g2646 ( 
.A1(n_2048),
.A2(n_1880),
.B1(n_1915),
.B2(n_1690),
.Y(n_2646)
);

AND2x2_ASAP7_75t_SL g2647 ( 
.A(n_2112),
.B(n_1781),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2107),
.Y(n_2648)
);

AND2x4_ASAP7_75t_L g2649 ( 
.A(n_2017),
.B(n_1720),
.Y(n_2649)
);

NOR2xp33_ASAP7_75t_L g2650 ( 
.A(n_2252),
.B(n_1857),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2123),
.Y(n_2651)
);

BUFx6f_ASAP7_75t_L g2652 ( 
.A(n_2087),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2172),
.Y(n_2653)
);

INVx4_ASAP7_75t_L g2654 ( 
.A(n_2087),
.Y(n_2654)
);

INVx3_ASAP7_75t_L g2655 ( 
.A(n_2093),
.Y(n_2655)
);

INVx4_ASAP7_75t_L g2656 ( 
.A(n_2093),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2172),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2174),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2174),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2194),
.B(n_1654),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2178),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2123),
.Y(n_2662)
);

AND3x2_ASAP7_75t_L g2663 ( 
.A(n_2215),
.B(n_1736),
.C(n_1675),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_SL g2664 ( 
.A(n_2149),
.B(n_1819),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2149),
.Y(n_2665)
);

NOR2xp33_ASAP7_75t_L g2666 ( 
.A(n_2263),
.B(n_1857),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2178),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2161),
.Y(n_2668)
);

CKINVDCx5p33_ASAP7_75t_R g2669 ( 
.A(n_2138),
.Y(n_2669)
);

OR2x6_ASAP7_75t_L g2670 ( 
.A(n_2162),
.B(n_1838),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2182),
.B(n_1741),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2194),
.B(n_1657),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2161),
.Y(n_2673)
);

CKINVDCx5p33_ASAP7_75t_R g2674 ( 
.A(n_2258),
.Y(n_2674)
);

AO21x2_ASAP7_75t_L g2675 ( 
.A1(n_2049),
.A2(n_1751),
.B(n_1714),
.Y(n_2675)
);

INVx5_ASAP7_75t_L g2676 ( 
.A(n_2210),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2193),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2182),
.Y(n_2678)
);

NOR2xp33_ASAP7_75t_L g2679 ( 
.A(n_2263),
.B(n_1914),
.Y(n_2679)
);

CKINVDCx5p33_ASAP7_75t_R g2680 ( 
.A(n_2258),
.Y(n_2680)
);

NOR2x1p5_ASAP7_75t_L g2681 ( 
.A(n_2199),
.B(n_1625),
.Y(n_2681)
);

BUFx6f_ASAP7_75t_SL g2682 ( 
.A(n_2299),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_SL g2683 ( 
.A(n_2193),
.B(n_1856),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2193),
.B(n_1659),
.Y(n_2684)
);

BUFx3_ASAP7_75t_L g2685 ( 
.A(n_1993),
.Y(n_2685)
);

INVx3_ASAP7_75t_L g2686 ( 
.A(n_2093),
.Y(n_2686)
);

INVx3_ASAP7_75t_L g2687 ( 
.A(n_2093),
.Y(n_2687)
);

INVx3_ASAP7_75t_L g2688 ( 
.A(n_2093),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_SL g2689 ( 
.A(n_2207),
.B(n_1858),
.Y(n_2689)
);

BUFx3_ASAP7_75t_L g2690 ( 
.A(n_1951),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_SL g2691 ( 
.A(n_2261),
.B(n_1914),
.Y(n_2691)
);

AOI21x1_ASAP7_75t_L g2692 ( 
.A1(n_1987),
.A2(n_1751),
.B(n_1714),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2195),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2195),
.Y(n_2694)
);

AND2x2_ASAP7_75t_SL g2695 ( 
.A(n_2049),
.B(n_1789),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2207),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2207),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_1973),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2306),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2306),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2660),
.B(n_1810),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2391),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2391),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2393),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2393),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2394),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2394),
.Y(n_2707)
);

XNOR2xp5_ASAP7_75t_L g2708 ( 
.A(n_2434),
.B(n_2171),
.Y(n_2708)
);

INVxp33_ASAP7_75t_SL g2709 ( 
.A(n_2456),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2404),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2404),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2443),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2473),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2473),
.Y(n_2714)
);

NOR2xp33_ASAP7_75t_L g2715 ( 
.A(n_2349),
.B(n_2184),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2474),
.Y(n_2716)
);

INVxp67_ASAP7_75t_SL g2717 ( 
.A(n_2412),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2474),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2475),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2475),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2346),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2346),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2660),
.B(n_1505),
.Y(n_2723)
);

AND2x2_ASAP7_75t_L g2724 ( 
.A(n_2672),
.B(n_2188),
.Y(n_2724)
);

INVx2_ASAP7_75t_SL g2725 ( 
.A(n_2555),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2352),
.Y(n_2726)
);

AND2x2_ASAP7_75t_L g2727 ( 
.A(n_2672),
.B(n_2372),
.Y(n_2727)
);

INVxp67_ASAP7_75t_L g2728 ( 
.A(n_2301),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_2456),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2352),
.Y(n_2730)
);

NOR2xp33_ASAP7_75t_L g2731 ( 
.A(n_2323),
.B(n_2223),
.Y(n_2731)
);

CKINVDCx5p33_ASAP7_75t_R g2732 ( 
.A(n_2669),
.Y(n_2732)
);

XOR2x2_ASAP7_75t_L g2733 ( 
.A(n_2434),
.B(n_2232),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2353),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2353),
.Y(n_2735)
);

NOR2xp33_ASAP7_75t_L g2736 ( 
.A(n_2449),
.B(n_2225),
.Y(n_2736)
);

OR2x6_ASAP7_75t_L g2737 ( 
.A(n_2541),
.B(n_2299),
.Y(n_2737)
);

NOR2xp33_ASAP7_75t_L g2738 ( 
.A(n_2314),
.B(n_2227),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2354),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2443),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2354),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2362),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2459),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2372),
.B(n_2384),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2362),
.Y(n_2745)
);

XOR2xp5_ASAP7_75t_L g2746 ( 
.A(n_2389),
.B(n_2294),
.Y(n_2746)
);

NOR2xp33_ASAP7_75t_L g2747 ( 
.A(n_2566),
.B(n_2228),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2459),
.Y(n_2748)
);

BUFx6f_ASAP7_75t_L g2749 ( 
.A(n_2350),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_SL g2750 ( 
.A(n_2565),
.B(n_2121),
.Y(n_2750)
);

NOR2xp33_ASAP7_75t_L g2751 ( 
.A(n_2347),
.B(n_2249),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2368),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2368),
.Y(n_2753)
);

BUFx6f_ASAP7_75t_SL g2754 ( 
.A(n_2462),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2373),
.Y(n_2755)
);

XOR2xp5_ASAP7_75t_L g2756 ( 
.A(n_2389),
.B(n_2294),
.Y(n_2756)
);

OAI21xp5_ASAP7_75t_L g2757 ( 
.A1(n_2326),
.A2(n_1990),
.B(n_2216),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2384),
.B(n_1766),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2373),
.Y(n_2759)
);

XNOR2xp5_ASAP7_75t_L g2760 ( 
.A(n_2669),
.B(n_2062),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2374),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2374),
.Y(n_2762)
);

NAND2xp33_ASAP7_75t_R g2763 ( 
.A(n_2572),
.B(n_2261),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2476),
.Y(n_2764)
);

INVx4_ASAP7_75t_SL g2765 ( 
.A(n_2304),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2460),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2476),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2478),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2478),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2460),
.Y(n_2770)
);

CKINVDCx16_ASAP7_75t_R g2771 ( 
.A(n_2462),
.Y(n_2771)
);

NAND2x1p5_ASAP7_75t_L g2772 ( 
.A(n_2333),
.B(n_1952),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2421),
.Y(n_2773)
);

HB1xp67_ASAP7_75t_L g2774 ( 
.A(n_2377),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2421),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2427),
.Y(n_2776)
);

AND2x4_ASAP7_75t_L g2777 ( 
.A(n_2387),
.B(n_1962),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2427),
.Y(n_2778)
);

BUFx6f_ASAP7_75t_L g2779 ( 
.A(n_2350),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2432),
.Y(n_2780)
);

NAND2x1p5_ASAP7_75t_L g2781 ( 
.A(n_2333),
.B(n_1952),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2432),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2468),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2436),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2436),
.Y(n_2785)
);

CKINVDCx14_ASAP7_75t_R g2786 ( 
.A(n_2303),
.Y(n_2786)
);

XNOR2xp5_ASAP7_75t_L g2787 ( 
.A(n_2647),
.B(n_1393),
.Y(n_2787)
);

AND2x2_ASAP7_75t_L g2788 ( 
.A(n_2331),
.B(n_1766),
.Y(n_2788)
);

XOR2xp5_ASAP7_75t_L g2789 ( 
.A(n_2674),
.B(n_1394),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2331),
.B(n_1937),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2385),
.Y(n_2791)
);

CKINVDCx16_ASAP7_75t_R g2792 ( 
.A(n_2462),
.Y(n_2792)
);

AND2x2_ASAP7_75t_L g2793 ( 
.A(n_2332),
.B(n_1938),
.Y(n_2793)
);

AND2x4_ASAP7_75t_L g2794 ( 
.A(n_2387),
.B(n_1965),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2385),
.Y(n_2795)
);

OR2x2_ASAP7_75t_L g2796 ( 
.A(n_2301),
.B(n_1555),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2317),
.B(n_2216),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2386),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2386),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2396),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2396),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2375),
.B(n_2216),
.Y(n_2802)
);

AND2x6_ASAP7_75t_L g2803 ( 
.A(n_2326),
.B(n_2327),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2398),
.Y(n_2804)
);

INVxp67_ASAP7_75t_L g2805 ( 
.A(n_2378),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2463),
.B(n_2234),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2468),
.Y(n_2807)
);

CKINVDCx20_ASAP7_75t_R g2808 ( 
.A(n_2303),
.Y(n_2808)
);

BUFx2_ASAP7_75t_L g2809 ( 
.A(n_2555),
.Y(n_2809)
);

INVx4_ASAP7_75t_SL g2810 ( 
.A(n_2304),
.Y(n_2810)
);

INVx1_ASAP7_75t_SL g2811 ( 
.A(n_2359),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2302),
.Y(n_2812)
);

CKINVDCx20_ASAP7_75t_R g2813 ( 
.A(n_2340),
.Y(n_2813)
);

OR2x2_ASAP7_75t_L g2814 ( 
.A(n_2378),
.B(n_1555),
.Y(n_2814)
);

AND2x2_ASAP7_75t_L g2815 ( 
.A(n_2332),
.B(n_1713),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2398),
.Y(n_2816)
);

XNOR2xp5_ASAP7_75t_L g2817 ( 
.A(n_2647),
.B(n_1420),
.Y(n_2817)
);

BUFx2_ASAP7_75t_L g2818 ( 
.A(n_2572),
.Y(n_2818)
);

CKINVDCx20_ASAP7_75t_R g2819 ( 
.A(n_2340),
.Y(n_2819)
);

CKINVDCx20_ASAP7_75t_R g2820 ( 
.A(n_2426),
.Y(n_2820)
);

XOR2xp5_ASAP7_75t_L g2821 ( 
.A(n_2674),
.B(n_1420),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2402),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2351),
.B(n_1219),
.Y(n_2823)
);

BUFx6f_ASAP7_75t_L g2824 ( 
.A(n_2350),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2402),
.Y(n_2825)
);

INVx3_ASAP7_75t_L g2826 ( 
.A(n_2350),
.Y(n_2826)
);

HB1xp67_ASAP7_75t_L g2827 ( 
.A(n_2320),
.Y(n_2827)
);

INVxp67_ASAP7_75t_SL g2828 ( 
.A(n_2412),
.Y(n_2828)
);

INVx2_ASAP7_75t_SL g2829 ( 
.A(n_2418),
.Y(n_2829)
);

AND2x2_ASAP7_75t_L g2830 ( 
.A(n_2351),
.B(n_1838),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2409),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_SL g2832 ( 
.A(n_2695),
.B(n_1952),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2302),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2409),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2308),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2411),
.Y(n_2836)
);

HB1xp67_ASAP7_75t_L g2837 ( 
.A(n_2431),
.Y(n_2837)
);

XNOR2xp5_ASAP7_75t_L g2838 ( 
.A(n_2500),
.B(n_1436),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2411),
.Y(n_2839)
);

NOR2xp33_ASAP7_75t_L g2840 ( 
.A(n_2561),
.B(n_2595),
.Y(n_2840)
);

AND2x2_ASAP7_75t_L g2841 ( 
.A(n_2363),
.B(n_1838),
.Y(n_2841)
);

NOR2xp33_ASAP7_75t_SL g2842 ( 
.A(n_2400),
.B(n_2280),
.Y(n_2842)
);

INVxp33_ASAP7_75t_SL g2843 ( 
.A(n_2490),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2308),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2416),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2416),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2310),
.Y(n_2847)
);

XOR2xp5_ASAP7_75t_L g2848 ( 
.A(n_2680),
.B(n_1436),
.Y(n_2848)
);

NOR2xp33_ASAP7_75t_L g2849 ( 
.A(n_2477),
.B(n_1786),
.Y(n_2849)
);

HB1xp67_ASAP7_75t_L g2850 ( 
.A(n_2435),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2310),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2311),
.Y(n_2852)
);

INVxp33_ASAP7_75t_L g2853 ( 
.A(n_2486),
.Y(n_2853)
);

NOR2xp33_ASAP7_75t_L g2854 ( 
.A(n_2484),
.B(n_1868),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2311),
.Y(n_2855)
);

BUFx2_ASAP7_75t_L g2856 ( 
.A(n_2549),
.Y(n_2856)
);

AND2x2_ASAP7_75t_L g2857 ( 
.A(n_2363),
.B(n_1720),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2313),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2313),
.Y(n_2859)
);

NOR2xp33_ASAP7_75t_L g2860 ( 
.A(n_2492),
.B(n_1967),
.Y(n_2860)
);

AND2x2_ASAP7_75t_L g2861 ( 
.A(n_2309),
.B(n_1722),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2315),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2315),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2325),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2497),
.B(n_1975),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2325),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2338),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2479),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2479),
.Y(n_2869)
);

CKINVDCx5p33_ASAP7_75t_R g2870 ( 
.A(n_2426),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2480),
.Y(n_2871)
);

HB1xp67_ASAP7_75t_L g2872 ( 
.A(n_2649),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2338),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2480),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2615),
.Y(n_2875)
);

AND2x2_ASAP7_75t_L g2876 ( 
.A(n_2581),
.B(n_1722),
.Y(n_2876)
);

NOR2xp67_ASAP7_75t_L g2877 ( 
.A(n_2494),
.B(n_2280),
.Y(n_2877)
);

AND2x4_ASAP7_75t_L g2878 ( 
.A(n_2414),
.B(n_2447),
.Y(n_2878)
);

OR2x2_ASAP7_75t_L g2879 ( 
.A(n_2408),
.B(n_1559),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2615),
.Y(n_2880)
);

NOR2xp67_ASAP7_75t_L g2881 ( 
.A(n_2395),
.B(n_1979),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2618),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2618),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2619),
.Y(n_2884)
);

OAI21xp5_ASAP7_75t_L g2885 ( 
.A1(n_2327),
.A2(n_2257),
.B(n_2234),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2341),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2619),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2621),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2341),
.Y(n_2889)
);

NOR2xp33_ASAP7_75t_L g2890 ( 
.A(n_2379),
.B(n_1982),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2344),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2581),
.B(n_1559),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2621),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2623),
.Y(n_2894)
);

CKINVDCx20_ASAP7_75t_R g2895 ( 
.A(n_2483),
.Y(n_2895)
);

NOR2xp33_ASAP7_75t_L g2896 ( 
.A(n_2382),
.B(n_1988),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2623),
.Y(n_2897)
);

XOR2x2_ASAP7_75t_L g2898 ( 
.A(n_2491),
.B(n_2513),
.Y(n_2898)
);

OR2x2_ASAP7_75t_L g2899 ( 
.A(n_2399),
.B(n_1574),
.Y(n_2899)
);

XOR2xp5_ASAP7_75t_L g2900 ( 
.A(n_2680),
.B(n_1443),
.Y(n_2900)
);

INVx2_ASAP7_75t_SL g2901 ( 
.A(n_2501),
.Y(n_2901)
);

XOR2xp5_ASAP7_75t_L g2902 ( 
.A(n_2441),
.B(n_1443),
.Y(n_2902)
);

AND2x2_ASAP7_75t_L g2903 ( 
.A(n_2501),
.B(n_1574),
.Y(n_2903)
);

XOR2xp5_ASAP7_75t_L g2904 ( 
.A(n_2441),
.B(n_1455),
.Y(n_2904)
);

AND2x4_ASAP7_75t_L g2905 ( 
.A(n_2414),
.B(n_2447),
.Y(n_2905)
);

INVx3_ASAP7_75t_L g2906 ( 
.A(n_2350),
.Y(n_2906)
);

CKINVDCx5p33_ASAP7_75t_R g2907 ( 
.A(n_2483),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2624),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2358),
.B(n_2388),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2624),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2626),
.Y(n_2911)
);

INVxp67_ASAP7_75t_L g2912 ( 
.A(n_2322),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2626),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2632),
.Y(n_2914)
);

AND2x2_ASAP7_75t_L g2915 ( 
.A(n_2413),
.B(n_1577),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2632),
.Y(n_2916)
);

CKINVDCx20_ASAP7_75t_R g2917 ( 
.A(n_2483),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2633),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2633),
.Y(n_2919)
);

INVx2_ASAP7_75t_SL g2920 ( 
.A(n_2685),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2637),
.Y(n_2921)
);

NOR2xp33_ASAP7_75t_L g2922 ( 
.A(n_2390),
.B(n_1992),
.Y(n_2922)
);

XOR2xp5_ASAP7_75t_L g2923 ( 
.A(n_2486),
.B(n_1455),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2637),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2588),
.B(n_1577),
.Y(n_2925)
);

NAND2xp33_ASAP7_75t_R g2926 ( 
.A(n_2591),
.B(n_2162),
.Y(n_2926)
);

CKINVDCx20_ASAP7_75t_R g2927 ( 
.A(n_2469),
.Y(n_2927)
);

INVxp33_ASAP7_75t_SL g2928 ( 
.A(n_2691),
.Y(n_2928)
);

XNOR2xp5_ASAP7_75t_L g2929 ( 
.A(n_2328),
.B(n_1472),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2344),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2348),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2348),
.Y(n_2932)
);

AND2x2_ASAP7_75t_L g2933 ( 
.A(n_2684),
.B(n_2234),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2357),
.Y(n_2934)
);

NOR2xp33_ASAP7_75t_L g2935 ( 
.A(n_2392),
.B(n_1679),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2357),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2360),
.Y(n_2937)
);

INVx1_ASAP7_75t_SL g2938 ( 
.A(n_2649),
.Y(n_2938)
);

CKINVDCx20_ASAP7_75t_R g2939 ( 
.A(n_2469),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2360),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2367),
.Y(n_2941)
);

BUFx6f_ASAP7_75t_L g2942 ( 
.A(n_2304),
.Y(n_2942)
);

AND2x4_ASAP7_75t_L g2943 ( 
.A(n_2454),
.B(n_2257),
.Y(n_2943)
);

CKINVDCx20_ASAP7_75t_R g2944 ( 
.A(n_2574),
.Y(n_2944)
);

XOR2xp5_ASAP7_75t_L g2945 ( 
.A(n_2489),
.B(n_1472),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2367),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2371),
.Y(n_2947)
);

XOR2xp5_ASAP7_75t_L g2948 ( 
.A(n_2489),
.B(n_1492),
.Y(n_2948)
);

INVxp67_ASAP7_75t_SL g2949 ( 
.A(n_2412),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2371),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2467),
.Y(n_2951)
);

AND2x2_ASAP7_75t_L g2952 ( 
.A(n_2684),
.B(n_2257),
.Y(n_2952)
);

NOR2xp33_ASAP7_75t_L g2953 ( 
.A(n_2406),
.B(n_1718),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2470),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2645),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2645),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2600),
.Y(n_2957)
);

NOR2xp33_ASAP7_75t_L g2958 ( 
.A(n_2417),
.B(n_1723),
.Y(n_2958)
);

AND2x2_ASAP7_75t_L g2959 ( 
.A(n_2425),
.B(n_1186),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2457),
.B(n_1587),
.Y(n_2960)
);

BUFx2_ASAP7_75t_L g2961 ( 
.A(n_2649),
.Y(n_2961)
);

NOR2xp67_ASAP7_75t_L g2962 ( 
.A(n_2430),
.B(n_1728),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2482),
.Y(n_2963)
);

AND2x2_ASAP7_75t_L g2964 ( 
.A(n_2563),
.B(n_1186),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2458),
.B(n_1587),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2600),
.Y(n_2966)
);

INVx8_ASAP7_75t_L g2967 ( 
.A(n_2541),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2602),
.Y(n_2968)
);

INVxp33_ASAP7_75t_L g2969 ( 
.A(n_2650),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2602),
.Y(n_2970)
);

XOR2xp5_ASAP7_75t_L g2971 ( 
.A(n_2603),
.B(n_1492),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2609),
.Y(n_2972)
);

INVxp33_ASAP7_75t_L g2973 ( 
.A(n_2666),
.Y(n_2973)
);

AND2x2_ASAP7_75t_L g2974 ( 
.A(n_2563),
.B(n_1337),
.Y(n_2974)
);

INVx3_ASAP7_75t_L g2975 ( 
.A(n_2412),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2482),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2461),
.B(n_1601),
.Y(n_2977)
);

CKINVDCx20_ASAP7_75t_R g2978 ( 
.A(n_2574),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2609),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2610),
.Y(n_2980)
);

NOR2xp33_ASAP7_75t_L g2981 ( 
.A(n_2593),
.B(n_777),
.Y(n_2981)
);

INVxp33_ASAP7_75t_L g2982 ( 
.A(n_2679),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2610),
.Y(n_2983)
);

NOR2xp33_ASAP7_75t_SL g2984 ( 
.A(n_2400),
.B(n_2258),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2614),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2614),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2318),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2319),
.Y(n_2988)
);

AOI21xp5_ASAP7_75t_L g2989 ( 
.A1(n_2671),
.A2(n_2016),
.B(n_1952),
.Y(n_2989)
);

XOR2x2_ASAP7_75t_L g2990 ( 
.A(n_2455),
.B(n_2130),
.Y(n_2990)
);

XOR2x2_ASAP7_75t_L g2991 ( 
.A(n_2472),
.B(n_2130),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2329),
.Y(n_2992)
);

NOR2x1_ASAP7_75t_L g2993 ( 
.A(n_2422),
.B(n_1710),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2485),
.Y(n_2994)
);

NOR2xp33_ASAP7_75t_L g2995 ( 
.A(n_2336),
.B(n_2307),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2337),
.Y(n_2996)
);

INVx1_ASAP7_75t_SL g2997 ( 
.A(n_2521),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2345),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2461),
.B(n_1601),
.Y(n_2999)
);

INVxp67_ASAP7_75t_SL g3000 ( 
.A(n_2412),
.Y(n_3000)
);

CKINVDCx5p33_ASAP7_75t_R g3001 ( 
.A(n_2336),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2424),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2433),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2438),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2440),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2444),
.Y(n_3006)
);

CKINVDCx5p33_ASAP7_75t_R g3007 ( 
.A(n_2336),
.Y(n_3007)
);

AND2x2_ASAP7_75t_L g3008 ( 
.A(n_2448),
.B(n_1337),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2445),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_SL g3010 ( 
.A(n_2606),
.B(n_2121),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2446),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2485),
.Y(n_3012)
);

AND2x6_ASAP7_75t_L g3013 ( 
.A(n_2334),
.B(n_2051),
.Y(n_3013)
);

XOR2xp5_ASAP7_75t_L g3014 ( 
.A(n_2608),
.B(n_1493),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2548),
.Y(n_3015)
);

XNOR2xp5_ASAP7_75t_L g3016 ( 
.A(n_2423),
.B(n_1493),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_SL g3017 ( 
.A(n_2695),
.B(n_1952),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2548),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_SL g3019 ( 
.A(n_2606),
.B(n_2616),
.Y(n_3019)
);

NOR2xp33_ASAP7_75t_SL g3020 ( 
.A(n_2400),
.B(n_2120),
.Y(n_3020)
);

XOR2x2_ASAP7_75t_L g3021 ( 
.A(n_2521),
.B(n_1502),
.Y(n_3021)
);

NOR2xp33_ASAP7_75t_L g3022 ( 
.A(n_2381),
.B(n_2052),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2559),
.Y(n_3023)
);

NOR2xp33_ASAP7_75t_L g3024 ( 
.A(n_2517),
.B(n_2058),
.Y(n_3024)
);

AND2x2_ASAP7_75t_L g3025 ( 
.A(n_2465),
.B(n_1370),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2559),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2696),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2696),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2697),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2493),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2697),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2553),
.Y(n_3032)
);

CKINVDCx5p33_ASAP7_75t_R g3033 ( 
.A(n_2670),
.Y(n_3033)
);

NOR2xp67_ASAP7_75t_L g3034 ( 
.A(n_2364),
.B(n_2060),
.Y(n_3034)
);

CKINVDCx20_ASAP7_75t_R g3035 ( 
.A(n_2670),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2554),
.Y(n_3036)
);

CKINVDCx20_ASAP7_75t_R g3037 ( 
.A(n_2670),
.Y(n_3037)
);

AOI21xp5_ASAP7_75t_L g3038 ( 
.A1(n_2407),
.A2(n_2131),
.B(n_1774),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2556),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2461),
.B(n_2121),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2557),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2564),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2573),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2576),
.Y(n_3044)
);

AND2x4_ASAP7_75t_L g3045 ( 
.A(n_2454),
.B(n_2061),
.Y(n_3045)
);

NOR2xp33_ASAP7_75t_L g3046 ( 
.A(n_2464),
.B(n_2065),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2578),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2585),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2594),
.Y(n_3049)
);

NAND2x1p5_ASAP7_75t_L g3050 ( 
.A(n_2333),
.B(n_2131),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2481),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2481),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2487),
.Y(n_3053)
);

AND2x2_ASAP7_75t_L g3054 ( 
.A(n_2364),
.B(n_2419),
.Y(n_3054)
);

AND2x4_ASAP7_75t_L g3055 ( 
.A(n_2466),
.B(n_2076),
.Y(n_3055)
);

NOR2xp33_ASAP7_75t_L g3056 ( 
.A(n_2562),
.B(n_2077),
.Y(n_3056)
);

INVx2_ASAP7_75t_SL g3057 ( 
.A(n_2685),
.Y(n_3057)
);

INVx2_ASAP7_75t_SL g3058 ( 
.A(n_2690),
.Y(n_3058)
);

AND2x2_ASAP7_75t_L g3059 ( 
.A(n_2419),
.B(n_1370),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2487),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2496),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2496),
.Y(n_3062)
);

XNOR2xp5_ASAP7_75t_L g3063 ( 
.A(n_2681),
.B(n_1502),
.Y(n_3063)
);

BUFx2_ASAP7_75t_L g3064 ( 
.A(n_2670),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2503),
.Y(n_3065)
);

NOR2xp33_ASAP7_75t_L g3066 ( 
.A(n_2582),
.B(n_2078),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2503),
.Y(n_3067)
);

CKINVDCx20_ASAP7_75t_R g3068 ( 
.A(n_2508),
.Y(n_3068)
);

NOR2xp33_ASAP7_75t_L g3069 ( 
.A(n_2519),
.B(n_2082),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2493),
.Y(n_3070)
);

AND2x2_ASAP7_75t_L g3071 ( 
.A(n_2616),
.B(n_1407),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2504),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2504),
.Y(n_3073)
);

HB1xp67_ASAP7_75t_L g3074 ( 
.A(n_2509),
.Y(n_3074)
);

OR2x6_ASAP7_75t_L g3075 ( 
.A(n_2541),
.B(n_2120),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2520),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2520),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2498),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2545),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2545),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_2498),
.Y(n_3081)
);

CKINVDCx16_ASAP7_75t_R g3082 ( 
.A(n_2682),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2547),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_2627),
.B(n_2628),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2502),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2547),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2653),
.Y(n_3087)
);

NOR2xp33_ASAP7_75t_SL g3088 ( 
.A(n_2407),
.B(n_2120),
.Y(n_3088)
);

INVxp67_ASAP7_75t_SL g3089 ( 
.A(n_2415),
.Y(n_3089)
);

AND2x6_ASAP7_75t_L g3090 ( 
.A(n_2334),
.B(n_2304),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2653),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2657),
.Y(n_3092)
);

INVxp67_ASAP7_75t_SL g3093 ( 
.A(n_2415),
.Y(n_3093)
);

CKINVDCx20_ASAP7_75t_R g3094 ( 
.A(n_2508),
.Y(n_3094)
);

XOR2x2_ASAP7_75t_L g3095 ( 
.A(n_2634),
.B(n_1504),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2657),
.Y(n_3096)
);

AND2x6_ASAP7_75t_L g3097 ( 
.A(n_2304),
.B(n_2090),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2658),
.Y(n_3098)
);

HB1xp67_ASAP7_75t_L g3099 ( 
.A(n_2509),
.Y(n_3099)
);

INVx2_ASAP7_75t_L g3100 ( 
.A(n_2712),
.Y(n_3100)
);

AOI22xp33_ASAP7_75t_L g3101 ( 
.A1(n_2840),
.A2(n_2662),
.B1(n_2665),
.B2(n_2651),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_L g3102 ( 
.A(n_2969),
.B(n_1504),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2764),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2909),
.B(n_2635),
.Y(n_3104)
);

OR2x2_ASAP7_75t_L g3105 ( 
.A(n_2840),
.B(n_2543),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2767),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2909),
.B(n_2531),
.Y(n_3107)
);

NAND2xp33_ASAP7_75t_L g3108 ( 
.A(n_2967),
.B(n_2380),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_2740),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2953),
.B(n_2550),
.Y(n_3110)
);

OAI21xp5_ASAP7_75t_L g3111 ( 
.A1(n_3040),
.A2(n_2343),
.B(n_2305),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_SL g3112 ( 
.A(n_2849),
.B(n_2627),
.Y(n_3112)
);

AND2x4_ASAP7_75t_SL g3113 ( 
.A(n_2837),
.B(n_2850),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2953),
.B(n_2552),
.Y(n_3114)
);

NOR2xp33_ASAP7_75t_L g3115 ( 
.A(n_2973),
.B(n_2452),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_SL g3116 ( 
.A(n_2849),
.B(n_2628),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2743),
.Y(n_3117)
);

NOR2xp33_ASAP7_75t_L g3118 ( 
.A(n_2982),
.B(n_2453),
.Y(n_3118)
);

INVx2_ASAP7_75t_SL g3119 ( 
.A(n_2829),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2958),
.B(n_2570),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2958),
.B(n_2580),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2912),
.B(n_2597),
.Y(n_3122)
);

INVxp67_ASAP7_75t_SL g3123 ( 
.A(n_2717),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2912),
.B(n_2598),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_SL g3125 ( 
.A(n_2854),
.B(n_2620),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2960),
.B(n_2646),
.Y(n_3126)
);

NOR2xp33_ASAP7_75t_L g3127 ( 
.A(n_2715),
.B(n_2935),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_SL g3128 ( 
.A(n_2854),
.B(n_2509),
.Y(n_3128)
);

NAND2xp33_ASAP7_75t_SL g3129 ( 
.A(n_2754),
.B(n_2682),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2768),
.Y(n_3130)
);

INVx2_ASAP7_75t_L g3131 ( 
.A(n_2748),
.Y(n_3131)
);

BUFx5_ASAP7_75t_L g3132 ( 
.A(n_3090),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2766),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_SL g3134 ( 
.A(n_2935),
.B(n_2509),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2770),
.Y(n_3135)
);

OR2x2_ASAP7_75t_L g3136 ( 
.A(n_2728),
.B(n_2532),
.Y(n_3136)
);

AND2x2_ASAP7_75t_L g3137 ( 
.A(n_2959),
.B(n_2370),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_2783),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2960),
.B(n_2370),
.Y(n_3139)
);

AOI22xp33_ASAP7_75t_L g3140 ( 
.A1(n_2898),
.A2(n_2305),
.B1(n_2370),
.B2(n_2366),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2769),
.Y(n_3141)
);

AOI22xp5_ASAP7_75t_L g3142 ( 
.A1(n_2915),
.A2(n_2744),
.B1(n_2997),
.B2(n_2727),
.Y(n_3142)
);

AOI22xp5_ASAP7_75t_L g3143 ( 
.A1(n_2997),
.A2(n_2558),
.B1(n_2641),
.B2(n_2636),
.Y(n_3143)
);

INVx3_ASAP7_75t_L g3144 ( 
.A(n_2749),
.Y(n_3144)
);

AOI22xp5_ASAP7_75t_L g3145 ( 
.A1(n_2815),
.A2(n_2689),
.B1(n_2683),
.B2(n_2664),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2860),
.B(n_2370),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_2860),
.B(n_2530),
.Y(n_3147)
);

AOI22xp5_ASAP7_75t_L g3148 ( 
.A1(n_2738),
.A2(n_2528),
.B1(n_2495),
.B2(n_2514),
.Y(n_3148)
);

AND2x6_ASAP7_75t_SL g3149 ( 
.A(n_2981),
.B(n_2508),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2699),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_2807),
.Y(n_3151)
);

NAND2xp33_ASAP7_75t_SL g3152 ( 
.A(n_2754),
.B(n_2682),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2865),
.B(n_2530),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2865),
.B(n_2534),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2700),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_2890),
.B(n_2534),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2890),
.B(n_2896),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2812),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2896),
.B(n_2540),
.Y(n_3159)
);

NOR3xp33_ASAP7_75t_L g3160 ( 
.A(n_2981),
.B(n_2316),
.C(n_2312),
.Y(n_3160)
);

AOI21xp5_ASAP7_75t_L g3161 ( 
.A1(n_2806),
.A2(n_2802),
.B(n_2797),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_SL g3162 ( 
.A(n_2802),
.B(n_2509),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2922),
.B(n_2540),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2833),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_2806),
.B(n_2415),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2922),
.B(n_2668),
.Y(n_3166)
);

INVxp67_ASAP7_75t_L g3167 ( 
.A(n_2837),
.Y(n_3167)
);

NOR2xp33_ASAP7_75t_L g3168 ( 
.A(n_2715),
.B(n_2410),
.Y(n_3168)
);

BUFx2_ASAP7_75t_L g3169 ( 
.A(n_2850),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_2738),
.B(n_2673),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2702),
.Y(n_3171)
);

OAI22xp33_ASAP7_75t_L g3172 ( 
.A1(n_2797),
.A2(n_2966),
.B1(n_2968),
.B2(n_2957),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2703),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_3024),
.B(n_2965),
.Y(n_3174)
);

NOR2xp33_ASAP7_75t_L g3175 ( 
.A(n_2995),
.B(n_2488),
.Y(n_3175)
);

NAND2xp33_ASAP7_75t_L g3176 ( 
.A(n_2967),
.B(n_2380),
.Y(n_3176)
);

NAND2xp33_ASAP7_75t_L g3177 ( 
.A(n_2967),
.B(n_2380),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_2835),
.Y(n_3178)
);

NOR2xp33_ASAP7_75t_L g3179 ( 
.A(n_2995),
.B(n_2355),
.Y(n_3179)
);

INVx3_ASAP7_75t_L g3180 ( 
.A(n_2749),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_2844),
.Y(n_3181)
);

NOR2xp33_ASAP7_75t_L g3182 ( 
.A(n_2728),
.B(n_2356),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_3024),
.B(n_2677),
.Y(n_3183)
);

OR2x6_ASAP7_75t_L g3184 ( 
.A(n_3075),
.B(n_2541),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_SL g3185 ( 
.A(n_2938),
.B(n_2701),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_SL g3186 ( 
.A(n_2938),
.B(n_2415),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2965),
.B(n_2415),
.Y(n_3187)
);

AOI22xp5_ASAP7_75t_L g3188 ( 
.A1(n_2901),
.A2(n_2343),
.B1(n_2403),
.B2(n_2330),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2704),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2857),
.B(n_2471),
.Y(n_3190)
);

NOR3xp33_ASAP7_75t_L g3191 ( 
.A(n_2747),
.B(n_2335),
.C(n_2321),
.Y(n_3191)
);

INVxp67_ASAP7_75t_L g3192 ( 
.A(n_2827),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_2758),
.B(n_2471),
.Y(n_3193)
);

NOR2x1p5_ASAP7_75t_L g3194 ( 
.A(n_2870),
.B(n_2466),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_SL g3195 ( 
.A(n_2811),
.B(n_2962),
.Y(n_3195)
);

INVx2_ASAP7_75t_SL g3196 ( 
.A(n_2809),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2861),
.B(n_2471),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_2963),
.Y(n_3198)
);

NOR2xp33_ASAP7_75t_SL g3199 ( 
.A(n_2709),
.B(n_2222),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2788),
.B(n_2471),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_2976),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_SL g3202 ( 
.A(n_2811),
.B(n_2471),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2705),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2706),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_2974),
.B(n_2499),
.Y(n_3205)
);

OAI221xp5_ASAP7_75t_L g3206 ( 
.A1(n_2838),
.A2(n_2405),
.B1(n_2376),
.B2(n_2361),
.C(n_2690),
.Y(n_3206)
);

NOR2xp33_ASAP7_75t_L g3207 ( 
.A(n_2805),
.B(n_2853),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_3059),
.B(n_2499),
.Y(n_3208)
);

INVxp67_ASAP7_75t_L g3209 ( 
.A(n_2827),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_2970),
.B(n_2596),
.Y(n_3210)
);

NOR2xp33_ASAP7_75t_L g3211 ( 
.A(n_2805),
.B(n_2599),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2972),
.B(n_2369),
.Y(n_3212)
);

HB1xp67_ASAP7_75t_L g3213 ( 
.A(n_2818),
.Y(n_3213)
);

NOR2x1p5_ASAP7_75t_L g3214 ( 
.A(n_2729),
.B(n_2222),
.Y(n_3214)
);

INVx6_ASAP7_75t_L g3215 ( 
.A(n_2878),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_2979),
.B(n_2369),
.Y(n_3216)
);

NOR2xp33_ASAP7_75t_L g3217 ( 
.A(n_2928),
.B(n_2451),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2980),
.B(n_2365),
.Y(n_3218)
);

O2A1O1Ixp33_ASAP7_75t_L g3219 ( 
.A1(n_3046),
.A2(n_1710),
.B(n_2401),
.C(n_2366),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2983),
.B(n_2365),
.Y(n_3220)
);

INVx2_ASAP7_75t_L g3221 ( 
.A(n_2994),
.Y(n_3221)
);

AOI22xp5_ASAP7_75t_L g3222 ( 
.A1(n_2747),
.A2(n_2439),
.B1(n_2437),
.B2(n_2617),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2985),
.B(n_2365),
.Y(n_3223)
);

AOI22xp5_ASAP7_75t_L g3224 ( 
.A1(n_2926),
.A2(n_2437),
.B1(n_2675),
.B2(n_2522),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_2986),
.B(n_2383),
.Y(n_3225)
);

OAI21xp33_ASAP7_75t_L g3226 ( 
.A1(n_2823),
.A2(n_1410),
.B(n_1407),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_SL g3227 ( 
.A(n_2830),
.B(n_2407),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_L g3228 ( 
.A(n_3022),
.B(n_2383),
.Y(n_3228)
);

INVx2_ASAP7_75t_SL g3229 ( 
.A(n_2725),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_SL g3230 ( 
.A(n_2841),
.B(n_2324),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_SL g3231 ( 
.A(n_2920),
.B(n_2324),
.Y(n_3231)
);

AND2x2_ASAP7_75t_L g3232 ( 
.A(n_2723),
.B(n_1916),
.Y(n_3232)
);

INVxp67_ASAP7_75t_L g3233 ( 
.A(n_2774),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_SL g3234 ( 
.A(n_3057),
.B(n_2324),
.Y(n_3234)
);

NOR2xp33_ASAP7_75t_L g3235 ( 
.A(n_2796),
.B(n_1598),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_SL g3236 ( 
.A(n_3058),
.B(n_2324),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_3022),
.B(n_2383),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_SL g3238 ( 
.A(n_2943),
.B(n_2324),
.Y(n_3238)
);

INVxp33_ASAP7_75t_L g3239 ( 
.A(n_2923),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_2876),
.B(n_2397),
.Y(n_3240)
);

INVx2_ASAP7_75t_SL g3241 ( 
.A(n_2774),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_2875),
.B(n_2397),
.Y(n_3242)
);

NAND2xp33_ASAP7_75t_SL g3243 ( 
.A(n_2926),
.B(n_2397),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_2880),
.B(n_2658),
.Y(n_3244)
);

BUFx5_ASAP7_75t_L g3245 ( 
.A(n_3090),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_2882),
.B(n_2659),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2707),
.Y(n_3247)
);

AND2x2_ASAP7_75t_L g3248 ( 
.A(n_2724),
.B(n_1916),
.Y(n_3248)
);

NOR2xp33_ASAP7_75t_L g3249 ( 
.A(n_2814),
.B(n_1617),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_SL g3250 ( 
.A(n_2943),
.B(n_2121),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2883),
.B(n_2659),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_SL g3252 ( 
.A(n_2790),
.B(n_2793),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_2884),
.B(n_2661),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_2887),
.B(n_2661),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_2888),
.B(n_2667),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_SL g3256 ( 
.A(n_2731),
.B(n_2125),
.Y(n_3256)
);

HB1xp67_ASAP7_75t_L g3257 ( 
.A(n_3074),
.Y(n_3257)
);

AND2x2_ASAP7_75t_SL g3258 ( 
.A(n_3088),
.B(n_2401),
.Y(n_3258)
);

INVx3_ASAP7_75t_L g3259 ( 
.A(n_2749),
.Y(n_3259)
);

NOR2xp33_ASAP7_75t_L g3260 ( 
.A(n_2856),
.B(n_1617),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_3012),
.Y(n_3261)
);

NOR2x1p5_ASAP7_75t_L g3262 ( 
.A(n_2732),
.B(n_2222),
.Y(n_3262)
);

AOI21xp5_ASAP7_75t_L g3263 ( 
.A1(n_2757),
.A2(n_2522),
.B(n_2380),
.Y(n_3263)
);

A2O1A1Ixp33_ASAP7_75t_L g3264 ( 
.A1(n_3069),
.A2(n_2678),
.B(n_2693),
.C(n_2667),
.Y(n_3264)
);

NOR2xp33_ASAP7_75t_L g3265 ( 
.A(n_2879),
.B(n_2569),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_2710),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_2893),
.B(n_2678),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_SL g3268 ( 
.A(n_2731),
.B(n_2125),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_SL g3269 ( 
.A(n_2878),
.B(n_2125),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_2894),
.B(n_2693),
.Y(n_3270)
);

INVx2_ASAP7_75t_L g3271 ( 
.A(n_3030),
.Y(n_3271)
);

AOI22xp5_ASAP7_75t_L g3272 ( 
.A1(n_2925),
.A2(n_2437),
.B1(n_2675),
.B2(n_2097),
.Y(n_3272)
);

O2A1O1Ixp5_ASAP7_75t_L g3273 ( 
.A1(n_2750),
.A2(n_2512),
.B(n_2692),
.C(n_2505),
.Y(n_3273)
);

AOI22xp5_ASAP7_75t_L g3274 ( 
.A1(n_2751),
.A2(n_2736),
.B1(n_2952),
.B2(n_2933),
.Y(n_3274)
);

INVx3_ASAP7_75t_L g3275 ( 
.A(n_2779),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_SL g3276 ( 
.A(n_2905),
.B(n_2125),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_2897),
.B(n_2908),
.Y(n_3277)
);

AOI22xp33_ASAP7_75t_L g3278 ( 
.A1(n_3046),
.A2(n_3069),
.B1(n_2999),
.B2(n_2977),
.Y(n_3278)
);

INVx1_ASAP7_75t_SL g3279 ( 
.A(n_2964),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_2910),
.B(n_2694),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2911),
.B(n_2694),
.Y(n_3281)
);

NAND2xp33_ASAP7_75t_L g3282 ( 
.A(n_3090),
.B(n_2537),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_3070),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_2913),
.B(n_2437),
.Y(n_3284)
);

AOI21xp5_ASAP7_75t_L g3285 ( 
.A1(n_2757),
.A2(n_2885),
.B(n_3040),
.Y(n_3285)
);

AOI22xp5_ASAP7_75t_L g3286 ( 
.A1(n_2751),
.A2(n_2675),
.B1(n_2098),
.B2(n_2101),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_2711),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_2914),
.B(n_2502),
.Y(n_3288)
);

AOI22xp5_ASAP7_75t_L g3289 ( 
.A1(n_2736),
.A2(n_2100),
.B1(n_2103),
.B2(n_2102),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_2916),
.B(n_2505),
.Y(n_3290)
);

AO221x1_ASAP7_75t_L g3291 ( 
.A1(n_2826),
.A2(n_2560),
.B1(n_2571),
.B2(n_2538),
.C(n_2515),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_2918),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_SL g3293 ( 
.A(n_2905),
.B(n_2127),
.Y(n_3293)
);

INVx2_ASAP7_75t_SL g3294 ( 
.A(n_2777),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_2919),
.B(n_2921),
.Y(n_3295)
);

AND2x6_ASAP7_75t_SL g3296 ( 
.A(n_3075),
.B(n_2508),
.Y(n_3296)
);

NAND2xp33_ASAP7_75t_L g3297 ( 
.A(n_3090),
.B(n_2643),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_3078),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_3081),
.Y(n_3299)
);

AOI22xp5_ASAP7_75t_L g3300 ( 
.A1(n_2892),
.A2(n_2105),
.B1(n_2124),
.B2(n_2119),
.Y(n_3300)
);

BUFx8_ASAP7_75t_L g3301 ( 
.A(n_3064),
.Y(n_3301)
);

HB1xp67_ASAP7_75t_L g3302 ( 
.A(n_3074),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_2924),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_3085),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3027),
.Y(n_3305)
);

HB1xp67_ASAP7_75t_L g3306 ( 
.A(n_3099),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_SL g3307 ( 
.A(n_2877),
.B(n_2127),
.Y(n_3307)
);

OAI22xp33_ASAP7_75t_L g3308 ( 
.A1(n_2987),
.A2(n_1514),
.B1(n_1517),
.B2(n_1410),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3071),
.B(n_2506),
.Y(n_3309)
);

INVxp33_ASAP7_75t_SL g3310 ( 
.A(n_2789),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3054),
.B(n_3051),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_SL g3312 ( 
.A(n_2881),
.B(n_2127),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_SL g3313 ( 
.A(n_2903),
.B(n_2127),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_3052),
.B(n_2506),
.Y(n_3314)
);

AND2x2_ASAP7_75t_L g3315 ( 
.A(n_3008),
.B(n_3025),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_SL g3316 ( 
.A(n_2872),
.B(n_2141),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3028),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3029),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_2867),
.Y(n_3319)
);

OR2x2_ASAP7_75t_L g3320 ( 
.A(n_2899),
.B(n_2708),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_3053),
.B(n_3060),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_SL g3322 ( 
.A(n_2872),
.B(n_2141),
.Y(n_3322)
);

NOR2xp33_ASAP7_75t_L g3323 ( 
.A(n_2945),
.B(n_2663),
.Y(n_3323)
);

NOR2xp33_ASAP7_75t_L g3324 ( 
.A(n_2948),
.B(n_2692),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_SL g3325 ( 
.A(n_2961),
.B(n_2141),
.Y(n_3325)
);

OR2x6_ASAP7_75t_L g3326 ( 
.A(n_3075),
.B(n_2631),
.Y(n_3326)
);

NOR2xp33_ASAP7_75t_L g3327 ( 
.A(n_2971),
.B(n_2631),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3061),
.B(n_2507),
.Y(n_3328)
);

AOI22xp33_ASAP7_75t_L g3329 ( 
.A1(n_2977),
.A2(n_968),
.B1(n_975),
.B2(n_956),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_2873),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_3062),
.B(n_2507),
.Y(n_3331)
);

NOR2xp33_ASAP7_75t_L g3332 ( 
.A(n_3014),
.B(n_2631),
.Y(n_3332)
);

NOR2xp33_ASAP7_75t_L g3333 ( 
.A(n_3001),
.B(n_2631),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3031),
.Y(n_3334)
);

OAI221xp5_ASAP7_75t_L g3335 ( 
.A1(n_3021),
.A2(n_969),
.B1(n_1009),
.B2(n_923),
.C(n_886),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_3065),
.B(n_2510),
.Y(n_3336)
);

OR2x6_ASAP7_75t_L g3337 ( 
.A(n_2737),
.B(n_2339),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_SL g3338 ( 
.A(n_3084),
.B(n_2141),
.Y(n_3338)
);

INVx2_ASAP7_75t_SL g3339 ( 
.A(n_2777),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_SL g3340 ( 
.A(n_2794),
.B(n_2153),
.Y(n_3340)
);

AND2x2_ASAP7_75t_L g3341 ( 
.A(n_2988),
.B(n_1514),
.Y(n_3341)
);

O2A1O1Ixp33_ASAP7_75t_L g3342 ( 
.A1(n_2999),
.A2(n_1907),
.B(n_1898),
.C(n_2510),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_2721),
.Y(n_3343)
);

AOI21xp5_ASAP7_75t_L g3344 ( 
.A1(n_2885),
.A2(n_2577),
.B(n_2523),
.Y(n_3344)
);

INVxp67_ASAP7_75t_SL g3345 ( 
.A(n_2717),
.Y(n_3345)
);

OR2x6_ASAP7_75t_L g3346 ( 
.A(n_2737),
.B(n_2339),
.Y(n_3346)
);

HB1xp67_ASAP7_75t_L g3347 ( 
.A(n_3099),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_2886),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_SL g3349 ( 
.A(n_2794),
.B(n_2153),
.Y(n_3349)
);

AOI22xp33_ASAP7_75t_L g3350 ( 
.A1(n_2719),
.A2(n_2126),
.B1(n_2136),
.B2(n_2129),
.Y(n_3350)
);

OR2x6_ASAP7_75t_L g3351 ( 
.A(n_2737),
.B(n_2339),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_SL g3352 ( 
.A(n_3032),
.B(n_2153),
.Y(n_3352)
);

AND2x6_ASAP7_75t_SL g3353 ( 
.A(n_2746),
.B(n_2038),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_3067),
.B(n_2511),
.Y(n_3354)
);

INVx2_ASAP7_75t_L g3355 ( 
.A(n_2889),
.Y(n_3355)
);

BUFx3_ASAP7_75t_L g3356 ( 
.A(n_2820),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_L g3357 ( 
.A(n_3072),
.B(n_2511),
.Y(n_3357)
);

BUFx8_ASAP7_75t_L g3358 ( 
.A(n_2992),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3073),
.B(n_2516),
.Y(n_3359)
);

CKINVDCx5p33_ASAP7_75t_R g3360 ( 
.A(n_2786),
.Y(n_3360)
);

NOR2xp33_ASAP7_75t_L g3361 ( 
.A(n_3007),
.B(n_2342),
.Y(n_3361)
);

NOR3xp33_ASAP7_75t_L g3362 ( 
.A(n_3056),
.B(n_2139),
.C(n_2137),
.Y(n_3362)
);

AOI22xp33_ASAP7_75t_L g3363 ( 
.A1(n_2996),
.A2(n_975),
.B1(n_977),
.B2(n_968),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_SL g3364 ( 
.A(n_3036),
.B(n_2153),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_3076),
.B(n_2516),
.Y(n_3365)
);

NOR2xp33_ASAP7_75t_L g3366 ( 
.A(n_3015),
.B(n_2342),
.Y(n_3366)
);

INVx2_ASAP7_75t_L g3367 ( 
.A(n_2891),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_3077),
.B(n_2518),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3079),
.B(n_2518),
.Y(n_3369)
);

BUFx8_ASAP7_75t_L g3370 ( 
.A(n_2998),
.Y(n_3370)
);

NOR2xp33_ASAP7_75t_L g3371 ( 
.A(n_3018),
.B(n_3023),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_2722),
.Y(n_3372)
);

AOI22xp5_ASAP7_75t_L g3373 ( 
.A1(n_3056),
.A2(n_2152),
.B1(n_2159),
.B2(n_2156),
.Y(n_3373)
);

NAND2xp33_ASAP7_75t_L g3374 ( 
.A(n_3090),
.B(n_2643),
.Y(n_3374)
);

NOR2xp33_ASAP7_75t_L g3375 ( 
.A(n_3026),
.B(n_2342),
.Y(n_3375)
);

OR2x2_ASAP7_75t_L g3376 ( 
.A(n_2787),
.B(n_2529),
.Y(n_3376)
);

AOI22xp5_ASAP7_75t_L g3377 ( 
.A1(n_3066),
.A2(n_2166),
.B1(n_2173),
.B2(n_2160),
.Y(n_3377)
);

OAI22xp33_ASAP7_75t_L g3378 ( 
.A1(n_3002),
.A2(n_3004),
.B1(n_3005),
.B2(n_3003),
.Y(n_3378)
);

AOI221xp5_ASAP7_75t_L g3379 ( 
.A1(n_3039),
.A2(n_1509),
.B1(n_1534),
.B2(n_1497),
.C(n_1445),
.Y(n_3379)
);

AND2x2_ASAP7_75t_L g3380 ( 
.A(n_3006),
.B(n_1517),
.Y(n_3380)
);

AND2x4_ASAP7_75t_L g3381 ( 
.A(n_3045),
.B(n_2429),
.Y(n_3381)
);

BUFx6f_ASAP7_75t_SL g3382 ( 
.A(n_3009),
.Y(n_3382)
);

INVx4_ASAP7_75t_L g3383 ( 
.A(n_2779),
.Y(n_3383)
);

BUFx6f_ASAP7_75t_L g3384 ( 
.A(n_2779),
.Y(n_3384)
);

AOI22xp33_ASAP7_75t_L g3385 ( 
.A1(n_3011),
.A2(n_978),
.B1(n_994),
.B2(n_977),
.Y(n_3385)
);

NOR2xp33_ASAP7_75t_L g3386 ( 
.A(n_2817),
.B(n_2843),
.Y(n_3386)
);

NOR2xp33_ASAP7_75t_L g3387 ( 
.A(n_2902),
.B(n_2512),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_SL g3388 ( 
.A(n_3041),
.B(n_2155),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3080),
.B(n_2524),
.Y(n_3389)
);

INVx2_ASAP7_75t_L g3390 ( 
.A(n_2934),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3083),
.B(n_2524),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_SL g3392 ( 
.A(n_3042),
.B(n_2155),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_2726),
.Y(n_3393)
);

AOI22xp33_ASAP7_75t_L g3394 ( 
.A1(n_3086),
.A2(n_994),
.B1(n_999),
.B2(n_978),
.Y(n_3394)
);

INVx5_ASAP7_75t_L g3395 ( 
.A(n_2803),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3066),
.B(n_2639),
.Y(n_3396)
);

NOR2xp33_ASAP7_75t_L g3397 ( 
.A(n_2904),
.B(n_2515),
.Y(n_3397)
);

NOR2xp67_ASAP7_75t_L g3398 ( 
.A(n_2907),
.B(n_3043),
.Y(n_3398)
);

INVx2_ASAP7_75t_L g3399 ( 
.A(n_2720),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3044),
.B(n_2639),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_3047),
.B(n_3048),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_2713),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3049),
.B(n_2640),
.Y(n_3403)
);

HB1xp67_ASAP7_75t_L g3404 ( 
.A(n_2765),
.Y(n_3404)
);

NOR2xp33_ASAP7_75t_L g3405 ( 
.A(n_2842),
.B(n_2515),
.Y(n_3405)
);

NAND2xp33_ASAP7_75t_L g3406 ( 
.A(n_2824),
.B(n_2942),
.Y(n_3406)
);

INVx3_ASAP7_75t_L g3407 ( 
.A(n_2824),
.Y(n_3407)
);

NOR2xp33_ASAP7_75t_L g3408 ( 
.A(n_2842),
.B(n_2538),
.Y(n_3408)
);

OR2x2_ASAP7_75t_L g3409 ( 
.A(n_2733),
.B(n_2526),
.Y(n_3409)
);

INVx2_ASAP7_75t_SL g3410 ( 
.A(n_3045),
.Y(n_3410)
);

AOI22xp5_ASAP7_75t_L g3411 ( 
.A1(n_2993),
.A2(n_2176),
.B1(n_2177),
.B2(n_2175),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_2828),
.B(n_2648),
.Y(n_3412)
);

O2A1O1Ixp33_ASAP7_75t_L g3413 ( 
.A1(n_2730),
.A2(n_1907),
.B(n_2526),
.C(n_2525),
.Y(n_3413)
);

INVx3_ASAP7_75t_L g3414 ( 
.A(n_2824),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_SL g3415 ( 
.A(n_3088),
.B(n_2155),
.Y(n_3415)
);

NOR2x1p5_ASAP7_75t_L g3416 ( 
.A(n_3033),
.B(n_3055),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_2828),
.B(n_2525),
.Y(n_3417)
);

BUFx6f_ASAP7_75t_L g3418 ( 
.A(n_2942),
.Y(n_3418)
);

INVxp67_ASAP7_75t_L g3419 ( 
.A(n_2763),
.Y(n_3419)
);

A2O1A1Ixp33_ASAP7_75t_L g3420 ( 
.A1(n_2951),
.A2(n_2442),
.B(n_2429),
.C(n_2527),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_2734),
.Y(n_3421)
);

INVx2_ASAP7_75t_L g3422 ( 
.A(n_2714),
.Y(n_3422)
);

AND2x2_ASAP7_75t_L g3423 ( 
.A(n_3055),
.B(n_1474),
.Y(n_3423)
);

INVx4_ASAP7_75t_L g3424 ( 
.A(n_2942),
.Y(n_3424)
);

OAI21xp5_ASAP7_75t_L g3425 ( 
.A1(n_2832),
.A2(n_2529),
.B(n_2527),
.Y(n_3425)
);

O2A1O1Ixp5_ASAP7_75t_L g3426 ( 
.A1(n_2832),
.A2(n_2535),
.B(n_2536),
.C(n_2533),
.Y(n_3426)
);

NOR2xp33_ASAP7_75t_L g3427 ( 
.A(n_2821),
.B(n_2848),
.Y(n_3427)
);

NOR2xp33_ASAP7_75t_L g3428 ( 
.A(n_2900),
.B(n_2538),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_2949),
.B(n_2533),
.Y(n_3429)
);

AOI22xp33_ASAP7_75t_L g3430 ( 
.A1(n_2735),
.A2(n_1000),
.B1(n_1011),
.B2(n_999),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_2949),
.B(n_2535),
.Y(n_3431)
);

INVxp33_ASAP7_75t_L g3432 ( 
.A(n_3063),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3000),
.B(n_2536),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_2739),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_2741),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3000),
.B(n_2640),
.Y(n_3436)
);

AND2x2_ASAP7_75t_L g3437 ( 
.A(n_2771),
.B(n_1475),
.Y(n_3437)
);

CKINVDCx5p33_ASAP7_75t_R g3438 ( 
.A(n_2763),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_2716),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_2742),
.Y(n_3440)
);

NOR3xp33_ASAP7_75t_L g3441 ( 
.A(n_2792),
.B(n_2183),
.C(n_2181),
.Y(n_3441)
);

NAND2xp33_ASAP7_75t_L g3442 ( 
.A(n_3097),
.B(n_2652),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_3089),
.B(n_2644),
.Y(n_3443)
);

O2A1O1Ixp33_ASAP7_75t_L g3444 ( 
.A1(n_2745),
.A2(n_2542),
.B(n_2544),
.C(n_2539),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_SL g3445 ( 
.A(n_3034),
.B(n_2155),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3089),
.B(n_2648),
.Y(n_3446)
);

AND2x2_ASAP7_75t_L g3447 ( 
.A(n_2990),
.B(n_1476),
.Y(n_3447)
);

NOR2xp33_ASAP7_75t_L g3448 ( 
.A(n_2760),
.B(n_2560),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_2752),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_2753),
.Y(n_3450)
);

NOR3xp33_ASAP7_75t_L g3451 ( 
.A(n_3019),
.B(n_2190),
.C(n_2186),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_SL g3452 ( 
.A(n_2984),
.B(n_2157),
.Y(n_3452)
);

INVx2_ASAP7_75t_L g3453 ( 
.A(n_2718),
.Y(n_3453)
);

INVx2_ASAP7_75t_L g3454 ( 
.A(n_2847),
.Y(n_3454)
);

INVxp67_ASAP7_75t_SL g3455 ( 
.A(n_3093),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3093),
.B(n_2539),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_2755),
.B(n_2542),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_2759),
.B(n_2544),
.Y(n_3458)
);

O2A1O1Ixp5_ASAP7_75t_L g3459 ( 
.A1(n_3017),
.A2(n_2956),
.B(n_2955),
.C(n_2762),
.Y(n_3459)
);

AOI22xp33_ASAP7_75t_L g3460 ( 
.A1(n_2761),
.A2(n_1011),
.B1(n_1014),
.B2(n_1000),
.Y(n_3460)
);

INVx4_ASAP7_75t_L g3461 ( 
.A(n_2765),
.Y(n_3461)
);

INVx5_ASAP7_75t_L g3462 ( 
.A(n_2803),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_2851),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_2868),
.B(n_2546),
.Y(n_3464)
);

OAI22xp33_ASAP7_75t_L g3465 ( 
.A1(n_2984),
.A2(n_1088),
.B1(n_1117),
.B2(n_1038),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_2869),
.B(n_2642),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_SL g3467 ( 
.A(n_3020),
.B(n_2157),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_2954),
.B(n_2642),
.Y(n_3468)
);

BUFx6f_ASAP7_75t_L g3469 ( 
.A(n_3097),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_2791),
.B(n_2644),
.Y(n_3470)
);

INVx2_ASAP7_75t_SL g3471 ( 
.A(n_3095),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_SL g3472 ( 
.A(n_3020),
.B(n_2157),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_2795),
.Y(n_3473)
);

INVx2_ASAP7_75t_L g3474 ( 
.A(n_2852),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_SL g3475 ( 
.A(n_2765),
.B(n_2157),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_SL g3476 ( 
.A(n_2810),
.B(n_2975),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_2798),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_2799),
.Y(n_3478)
);

HB1xp67_ASAP7_75t_L g3479 ( 
.A(n_2810),
.Y(n_3479)
);

INVx2_ASAP7_75t_SL g3480 ( 
.A(n_2991),
.Y(n_3480)
);

NOR2xp33_ASAP7_75t_L g3481 ( 
.A(n_3017),
.B(n_2929),
.Y(n_3481)
);

INVx3_ASAP7_75t_L g3482 ( 
.A(n_2826),
.Y(n_3482)
);

NOR2xp33_ASAP7_75t_L g3483 ( 
.A(n_3127),
.B(n_3016),
.Y(n_3483)
);

NOR3xp33_ASAP7_75t_L g3484 ( 
.A(n_3335),
.B(n_3249),
.C(n_3235),
.Y(n_3484)
);

O2A1O1Ixp33_ASAP7_75t_L g3485 ( 
.A1(n_3157),
.A2(n_2201),
.B(n_2202),
.C(n_2191),
.Y(n_3485)
);

AND2x4_ASAP7_75t_L g3486 ( 
.A(n_3416),
.B(n_2810),
.Y(n_3486)
);

OR2x2_ASAP7_75t_L g3487 ( 
.A(n_3105),
.B(n_3082),
.Y(n_3487)
);

AOI21xp5_ASAP7_75t_L g3488 ( 
.A1(n_3263),
.A2(n_3038),
.B(n_2781),
.Y(n_3488)
);

BUFx2_ASAP7_75t_SL g3489 ( 
.A(n_3119),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3292),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3107),
.B(n_2800),
.Y(n_3491)
);

NOR2xp33_ASAP7_75t_L g3492 ( 
.A(n_3168),
.B(n_2895),
.Y(n_3492)
);

A2O1A1Ixp33_ASAP7_75t_L g3493 ( 
.A1(n_3104),
.A2(n_2989),
.B(n_2804),
.C(n_2816),
.Y(n_3493)
);

AOI21xp5_ASAP7_75t_L g3494 ( 
.A1(n_3263),
.A2(n_3161),
.B(n_3038),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3303),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3315),
.B(n_3035),
.Y(n_3496)
);

INVx2_ASAP7_75t_SL g3497 ( 
.A(n_3113),
.Y(n_3497)
);

OAI21xp33_ASAP7_75t_L g3498 ( 
.A1(n_3122),
.A2(n_1151),
.B(n_1135),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3110),
.B(n_2801),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3114),
.B(n_2822),
.Y(n_3500)
);

AO21x1_ASAP7_75t_L g3501 ( 
.A1(n_3172),
.A2(n_3134),
.B(n_3128),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3120),
.B(n_2825),
.Y(n_3502)
);

BUFx12f_ASAP7_75t_L g3503 ( 
.A(n_3296),
.Y(n_3503)
);

AOI21x1_ASAP7_75t_L g3504 ( 
.A1(n_3161),
.A2(n_2989),
.B(n_3010),
.Y(n_3504)
);

INVx4_ASAP7_75t_L g3505 ( 
.A(n_3461),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3121),
.B(n_2831),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3124),
.B(n_2834),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3174),
.B(n_2836),
.Y(n_3508)
);

INVx4_ASAP7_75t_L g3509 ( 
.A(n_3461),
.Y(n_3509)
);

AOI21xp5_ASAP7_75t_L g3510 ( 
.A1(n_3282),
.A2(n_3374),
.B(n_3297),
.Y(n_3510)
);

AOI21xp5_ASAP7_75t_L g3511 ( 
.A1(n_3344),
.A2(n_2781),
.B(n_2772),
.Y(n_3511)
);

AOI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_3344),
.A2(n_3050),
.B(n_2772),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3402),
.Y(n_3513)
);

AO21x1_ASAP7_75t_L g3514 ( 
.A1(n_3172),
.A2(n_3091),
.B(n_3087),
.Y(n_3514)
);

AOI21xp5_ASAP7_75t_L g3515 ( 
.A1(n_3442),
.A2(n_3050),
.B(n_2577),
.Y(n_3515)
);

INVx3_ASAP7_75t_L g3516 ( 
.A(n_3469),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3150),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_3170),
.B(n_3278),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3278),
.B(n_2839),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3155),
.Y(n_3520)
);

NOR2xp33_ASAP7_75t_L g3521 ( 
.A(n_3102),
.B(n_2917),
.Y(n_3521)
);

NAND2xp33_ASAP7_75t_L g3522 ( 
.A(n_3191),
.B(n_3097),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_3166),
.B(n_2845),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3171),
.Y(n_3524)
);

AOI21xp5_ASAP7_75t_L g3525 ( 
.A1(n_3228),
.A2(n_2577),
.B(n_2523),
.Y(n_3525)
);

AOI22xp5_ASAP7_75t_L g3526 ( 
.A1(n_3387),
.A2(n_3037),
.B1(n_2846),
.B2(n_3068),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_3175),
.B(n_2803),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3274),
.B(n_2803),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3147),
.B(n_2803),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3153),
.B(n_2773),
.Y(n_3530)
);

INVxp67_ASAP7_75t_L g3531 ( 
.A(n_3169),
.Y(n_3531)
);

BUFx12f_ASAP7_75t_L g3532 ( 
.A(n_3358),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_3154),
.B(n_2775),
.Y(n_3533)
);

AOI21xp5_ASAP7_75t_L g3534 ( 
.A1(n_3237),
.A2(n_2589),
.B(n_2523),
.Y(n_3534)
);

OAI21xp5_ASAP7_75t_L g3535 ( 
.A1(n_3125),
.A2(n_2778),
.B(n_2776),
.Y(n_3535)
);

NAND3xp33_ASAP7_75t_L g3536 ( 
.A(n_3160),
.B(n_2047),
.C(n_2038),
.Y(n_3536)
);

OR2x2_ASAP7_75t_L g3537 ( 
.A(n_3320),
.B(n_2780),
.Y(n_3537)
);

AND2x2_ASAP7_75t_L g3538 ( 
.A(n_3232),
.B(n_2855),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3173),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3422),
.Y(n_3540)
);

NAND2x1_ASAP7_75t_L g3541 ( 
.A(n_3469),
.B(n_3097),
.Y(n_3541)
);

A2O1A1Ixp33_ASAP7_75t_L g3542 ( 
.A1(n_3219),
.A2(n_2784),
.B(n_2785),
.C(n_2782),
.Y(n_3542)
);

NOR2xp33_ASAP7_75t_L g3543 ( 
.A(n_3179),
.B(n_2756),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_3156),
.B(n_2871),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3159),
.B(n_2874),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3189),
.Y(n_3546)
);

AOI21xp5_ASAP7_75t_L g3547 ( 
.A1(n_3285),
.A2(n_2592),
.B(n_2589),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3203),
.Y(n_3548)
);

NOR2xp33_ASAP7_75t_L g3549 ( 
.A(n_3419),
.B(n_2927),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3163),
.B(n_2930),
.Y(n_3550)
);

INVx2_ASAP7_75t_L g3551 ( 
.A(n_3439),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3200),
.B(n_2931),
.Y(n_3552)
);

NOR2xp33_ASAP7_75t_L g3553 ( 
.A(n_3419),
.B(n_2939),
.Y(n_3553)
);

OAI21xp5_ASAP7_75t_L g3554 ( 
.A1(n_3126),
.A2(n_2936),
.B(n_2932),
.Y(n_3554)
);

AOI21xp5_ASAP7_75t_L g3555 ( 
.A1(n_3285),
.A2(n_2592),
.B(n_2589),
.Y(n_3555)
);

OAI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_3219),
.A2(n_2940),
.B(n_2937),
.Y(n_3556)
);

AOI21xp5_ASAP7_75t_L g3557 ( 
.A1(n_3111),
.A2(n_3345),
.B(n_3123),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3204),
.Y(n_3558)
);

AOI21xp5_ASAP7_75t_L g3559 ( 
.A1(n_3123),
.A2(n_2630),
.B(n_2592),
.Y(n_3559)
);

AOI21xp5_ASAP7_75t_L g3560 ( 
.A1(n_3345),
.A2(n_3455),
.B(n_3258),
.Y(n_3560)
);

A2O1A1Ixp33_ASAP7_75t_L g3561 ( 
.A1(n_3145),
.A2(n_2946),
.B(n_2947),
.C(n_2941),
.Y(n_3561)
);

NOR3xp33_ASAP7_75t_L g3562 ( 
.A(n_3465),
.B(n_3217),
.C(n_3206),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3142),
.B(n_2950),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3193),
.B(n_2858),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3183),
.B(n_2859),
.Y(n_3565)
);

HB1xp67_ASAP7_75t_L g3566 ( 
.A(n_3213),
.Y(n_3566)
);

AOI21xp5_ASAP7_75t_L g3567 ( 
.A1(n_3455),
.A2(n_2654),
.B(n_2630),
.Y(n_3567)
);

OR2x6_ASAP7_75t_L g3568 ( 
.A(n_3184),
.B(n_2906),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3247),
.Y(n_3569)
);

INVx3_ASAP7_75t_L g3570 ( 
.A(n_3469),
.Y(n_3570)
);

NOR2xp33_ASAP7_75t_L g3571 ( 
.A(n_3376),
.B(n_2944),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3266),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3287),
.Y(n_3573)
);

AOI21xp5_ASAP7_75t_L g3574 ( 
.A1(n_3258),
.A2(n_2654),
.B(n_2630),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3248),
.B(n_2862),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3343),
.Y(n_3576)
);

O2A1O1Ixp5_ASAP7_75t_L g3577 ( 
.A1(n_3415),
.A2(n_2906),
.B(n_2975),
.C(n_3092),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_SL g3578 ( 
.A(n_3207),
.B(n_2978),
.Y(n_3578)
);

NAND2xp33_ASAP7_75t_L g3579 ( 
.A(n_3191),
.B(n_3097),
.Y(n_3579)
);

OAI21xp33_ASAP7_75t_L g3580 ( 
.A1(n_3226),
.A2(n_3148),
.B(n_3341),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3311),
.B(n_2863),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3372),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3205),
.B(n_2864),
.Y(n_3583)
);

AOI21xp5_ASAP7_75t_L g3584 ( 
.A1(n_3108),
.A2(n_2656),
.B(n_2654),
.Y(n_3584)
);

OR2x6_ASAP7_75t_L g3585 ( 
.A(n_3184),
.B(n_2866),
.Y(n_3585)
);

AOI21xp5_ASAP7_75t_L g3586 ( 
.A1(n_3176),
.A2(n_2656),
.B(n_2622),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3208),
.B(n_3096),
.Y(n_3587)
);

AOI21xp5_ASAP7_75t_L g3588 ( 
.A1(n_3177),
.A2(n_2656),
.B(n_2622),
.Y(n_3588)
);

AOI21xp5_ASAP7_75t_L g3589 ( 
.A1(n_3112),
.A2(n_2622),
.B(n_2537),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3393),
.Y(n_3590)
);

BUFx6f_ASAP7_75t_L g3591 ( 
.A(n_3418),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3421),
.Y(n_3592)
);

INVx2_ASAP7_75t_L g3593 ( 
.A(n_3453),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3380),
.B(n_3098),
.Y(n_3594)
);

AOI21xp5_ASAP7_75t_L g3595 ( 
.A1(n_3116),
.A2(n_2622),
.B(n_2537),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3252),
.B(n_2546),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3212),
.A2(n_2622),
.B(n_2537),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3434),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3216),
.A2(n_2643),
.B(n_2537),
.Y(n_3599)
);

HB1xp67_ASAP7_75t_L g3600 ( 
.A(n_3213),
.Y(n_3600)
);

OAI21xp5_ASAP7_75t_L g3601 ( 
.A1(n_3459),
.A2(n_2567),
.B(n_2551),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_SL g3602 ( 
.A(n_3279),
.B(n_3094),
.Y(n_3602)
);

AOI22xp33_ASAP7_75t_SL g3603 ( 
.A1(n_3471),
.A2(n_3481),
.B1(n_3199),
.B2(n_3386),
.Y(n_3603)
);

AOI21xp5_ASAP7_75t_L g3604 ( 
.A1(n_3187),
.A2(n_2652),
.B(n_2643),
.Y(n_3604)
);

O2A1O1Ixp33_ASAP7_75t_L g3605 ( 
.A1(n_3465),
.A2(n_1159),
.B(n_1017),
.C(n_1020),
.Y(n_3605)
);

NOR2xp67_ASAP7_75t_L g3606 ( 
.A(n_3143),
.B(n_2560),
.Y(n_3606)
);

BUFx6f_ASAP7_75t_L g3607 ( 
.A(n_3418),
.Y(n_3607)
);

AOI21xp5_ASAP7_75t_L g3608 ( 
.A1(n_3240),
.A2(n_2652),
.B(n_2643),
.Y(n_3608)
);

O2A1O1Ixp5_ASAP7_75t_L g3609 ( 
.A1(n_3452),
.A2(n_2567),
.B(n_2568),
.C(n_2551),
.Y(n_3609)
);

AOI21xp5_ASAP7_75t_L g3610 ( 
.A1(n_3243),
.A2(n_2652),
.B(n_2676),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_3139),
.B(n_3137),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_3115),
.B(n_2568),
.Y(n_3612)
);

O2A1O1Ixp33_ASAP7_75t_L g3613 ( 
.A1(n_3160),
.A2(n_1017),
.B(n_1020),
.C(n_1014),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3118),
.B(n_2575),
.Y(n_3614)
);

AOI21xp5_ASAP7_75t_L g3615 ( 
.A1(n_3227),
.A2(n_2652),
.B(n_2676),
.Y(n_3615)
);

NOR3xp33_ASAP7_75t_L g3616 ( 
.A(n_3265),
.B(n_1026),
.C(n_1023),
.Y(n_3616)
);

BUFx6f_ASAP7_75t_L g3617 ( 
.A(n_3418),
.Y(n_3617)
);

NOR2xp33_ASAP7_75t_SL g3618 ( 
.A(n_3360),
.B(n_2808),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_3447),
.B(n_1477),
.Y(n_3619)
);

AOI21xp5_ASAP7_75t_L g3620 ( 
.A1(n_3162),
.A2(n_2676),
.B(n_2428),
.Y(n_3620)
);

INVx2_ASAP7_75t_L g3621 ( 
.A(n_3454),
.Y(n_3621)
);

AOI33xp33_ASAP7_75t_L g3622 ( 
.A1(n_3379),
.A2(n_1482),
.A3(n_1480),
.B1(n_1483),
.B2(n_1481),
.B3(n_1478),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3435),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_SL g3624 ( 
.A(n_3438),
.B(n_2180),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_SL g3625 ( 
.A(n_3167),
.B(n_2180),
.Y(n_3625)
);

NAND2x1p5_ASAP7_75t_L g3626 ( 
.A(n_3395),
.B(n_2571),
.Y(n_3626)
);

AND2x2_ASAP7_75t_SL g3627 ( 
.A(n_3140),
.B(n_1023),
.Y(n_3627)
);

INVx11_ASAP7_75t_L g3628 ( 
.A(n_3301),
.Y(n_3628)
);

BUFx6f_ASAP7_75t_L g3629 ( 
.A(n_3384),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_SL g3630 ( 
.A(n_3167),
.B(n_2180),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_3371),
.B(n_3146),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3440),
.Y(n_3632)
);

OAI21xp5_ASAP7_75t_L g3633 ( 
.A1(n_3459),
.A2(n_2579),
.B(n_2575),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3423),
.B(n_1484),
.Y(n_3634)
);

AOI21xp5_ASAP7_75t_L g3635 ( 
.A1(n_3224),
.A2(n_2676),
.B(n_2450),
.Y(n_3635)
);

BUFx6f_ASAP7_75t_L g3636 ( 
.A(n_3384),
.Y(n_3636)
);

CKINVDCx5p33_ASAP7_75t_R g3637 ( 
.A(n_3353),
.Y(n_3637)
);

OAI22xp5_ASAP7_75t_L g3638 ( 
.A1(n_3222),
.A2(n_2420),
.B1(n_2686),
.B2(n_2655),
.Y(n_3638)
);

HB1xp67_ASAP7_75t_L g3639 ( 
.A(n_3241),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_SL g3640 ( 
.A(n_3196),
.B(n_2180),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_3463),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3309),
.B(n_2579),
.Y(n_3642)
);

AOI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_3165),
.A2(n_2676),
.B(n_1774),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3401),
.B(n_2583),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_SL g3645 ( 
.A(n_3448),
.B(n_2187),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3449),
.Y(n_3646)
);

BUFx2_ASAP7_75t_L g3647 ( 
.A(n_3192),
.Y(n_3647)
);

HB1xp67_ASAP7_75t_L g3648 ( 
.A(n_3192),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_3185),
.B(n_2583),
.Y(n_3649)
);

AOI21xp5_ASAP7_75t_L g3650 ( 
.A1(n_3396),
.A2(n_1774),
.B(n_1773),
.Y(n_3650)
);

OAI22xp5_ASAP7_75t_L g3651 ( 
.A1(n_3140),
.A2(n_2686),
.B1(n_2687),
.B2(n_2655),
.Y(n_3651)
);

AOI21x1_ASAP7_75t_L g3652 ( 
.A1(n_3256),
.A2(n_2586),
.B(n_2584),
.Y(n_3652)
);

AOI21xp5_ASAP7_75t_L g3653 ( 
.A1(n_3406),
.A2(n_1774),
.B(n_1773),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3211),
.B(n_2584),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_SL g3655 ( 
.A(n_3409),
.B(n_2187),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3378),
.B(n_3277),
.Y(n_3656)
);

BUFx2_ASAP7_75t_L g3657 ( 
.A(n_3209),
.Y(n_3657)
);

BUFx8_ASAP7_75t_L g3658 ( 
.A(n_3382),
.Y(n_3658)
);

OR2x2_ASAP7_75t_L g3659 ( 
.A(n_3324),
.B(n_2586),
.Y(n_3659)
);

INVx3_ASAP7_75t_L g3660 ( 
.A(n_3395),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3378),
.B(n_2587),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3295),
.B(n_2587),
.Y(n_3662)
);

HB1xp67_ASAP7_75t_L g3663 ( 
.A(n_3209),
.Y(n_3663)
);

AOI21xp5_ASAP7_75t_L g3664 ( 
.A1(n_3395),
.A2(n_1776),
.B(n_1773),
.Y(n_3664)
);

AOI21xp5_ASAP7_75t_L g3665 ( 
.A1(n_3395),
.A2(n_1776),
.B(n_1773),
.Y(n_3665)
);

NOR2xp33_ASAP7_75t_L g3666 ( 
.A(n_3432),
.B(n_2813),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3474),
.Y(n_3667)
);

AOI21xp5_ASAP7_75t_L g3668 ( 
.A1(n_3462),
.A2(n_1785),
.B(n_1776),
.Y(n_3668)
);

NOR2xp33_ASAP7_75t_L g3669 ( 
.A(n_3239),
.B(n_2819),
.Y(n_3669)
);

O2A1O1Ixp33_ASAP7_75t_L g3670 ( 
.A1(n_3195),
.A2(n_1027),
.B(n_1029),
.C(n_1026),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3399),
.Y(n_3671)
);

AOI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_3462),
.A2(n_1785),
.B(n_1776),
.Y(n_3672)
);

OAI22xp5_ASAP7_75t_L g3673 ( 
.A1(n_3101),
.A2(n_2686),
.B1(n_2687),
.B2(n_2655),
.Y(n_3673)
);

BUFx6f_ASAP7_75t_L g3674 ( 
.A(n_3384),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_3321),
.B(n_2590),
.Y(n_3675)
);

AOI22xp5_ASAP7_75t_L g3676 ( 
.A1(n_3182),
.A2(n_3013),
.B1(n_821),
.B2(n_830),
.Y(n_3676)
);

AOI21xp5_ASAP7_75t_L g3677 ( 
.A1(n_3462),
.A2(n_3420),
.B(n_3197),
.Y(n_3677)
);

OR2x2_ASAP7_75t_L g3678 ( 
.A(n_3136),
.B(n_2625),
.Y(n_3678)
);

BUFx3_ASAP7_75t_L g3679 ( 
.A(n_3301),
.Y(n_3679)
);

INVx2_ASAP7_75t_L g3680 ( 
.A(n_3103),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3190),
.B(n_2590),
.Y(n_3681)
);

INVxp67_ASAP7_75t_L g3682 ( 
.A(n_3437),
.Y(n_3682)
);

NOR2xp33_ASAP7_75t_L g3683 ( 
.A(n_3397),
.B(n_2698),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_L g3684 ( 
.A(n_3106),
.B(n_2601),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_L g3685 ( 
.A(n_3130),
.B(n_2601),
.Y(n_3685)
);

BUFx3_ASAP7_75t_L g3686 ( 
.A(n_3229),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_SL g3687 ( 
.A(n_3398),
.B(n_2187),
.Y(n_3687)
);

OAI22xp5_ASAP7_75t_L g3688 ( 
.A1(n_3381),
.A2(n_2688),
.B1(n_2687),
.B2(n_2442),
.Y(n_3688)
);

AOI21xp5_ASAP7_75t_L g3689 ( 
.A1(n_3462),
.A2(n_3342),
.B(n_3412),
.Y(n_3689)
);

NOR2xp33_ASAP7_75t_L g3690 ( 
.A(n_3428),
.B(n_2698),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_SL g3691 ( 
.A(n_3233),
.B(n_2187),
.Y(n_3691)
);

OAI21xp5_ASAP7_75t_L g3692 ( 
.A1(n_3272),
.A2(n_2607),
.B(n_2605),
.Y(n_3692)
);

NOR2x1p5_ASAP7_75t_L g3693 ( 
.A(n_3356),
.B(n_2038),
.Y(n_3693)
);

AOI21xp5_ASAP7_75t_L g3694 ( 
.A1(n_3342),
.A2(n_1787),
.B(n_1785),
.Y(n_3694)
);

INVxp67_ASAP7_75t_L g3695 ( 
.A(n_3233),
.Y(n_3695)
);

NOR2x1_ASAP7_75t_L g3696 ( 
.A(n_3383),
.B(n_3424),
.Y(n_3696)
);

AOI21xp5_ASAP7_75t_L g3697 ( 
.A1(n_3417),
.A2(n_1787),
.B(n_1785),
.Y(n_3697)
);

BUFx5_ASAP7_75t_L g3698 ( 
.A(n_3473),
.Y(n_3698)
);

AOI21xp5_ASAP7_75t_L g3699 ( 
.A1(n_3429),
.A2(n_1793),
.B(n_1787),
.Y(n_3699)
);

AOI21xp5_ASAP7_75t_L g3700 ( 
.A1(n_3431),
.A2(n_1793),
.B(n_1787),
.Y(n_3700)
);

INVx4_ASAP7_75t_L g3701 ( 
.A(n_3215),
.Y(n_3701)
);

A2O1A1Ixp33_ASAP7_75t_L g3702 ( 
.A1(n_3188),
.A2(n_2607),
.B(n_2611),
.C(n_2605),
.Y(n_3702)
);

AOI21xp5_ASAP7_75t_L g3703 ( 
.A1(n_3433),
.A2(n_1795),
.B(n_1793),
.Y(n_3703)
);

CKINVDCx10_ASAP7_75t_R g3704 ( 
.A(n_3382),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3141),
.Y(n_3705)
);

AOI21xp5_ASAP7_75t_L g3706 ( 
.A1(n_3436),
.A2(n_1795),
.B(n_1793),
.Y(n_3706)
);

OAI21xp5_ASAP7_75t_L g3707 ( 
.A1(n_3286),
.A2(n_2612),
.B(n_2611),
.Y(n_3707)
);

AOI21x1_ASAP7_75t_L g3708 ( 
.A1(n_3268),
.A2(n_2613),
.B(n_2612),
.Y(n_3708)
);

INVx3_ASAP7_75t_L g3709 ( 
.A(n_3381),
.Y(n_3709)
);

AOI21xp5_ASAP7_75t_L g3710 ( 
.A1(n_3443),
.A2(n_1821),
.B(n_1795),
.Y(n_3710)
);

AOI21x1_ASAP7_75t_L g3711 ( 
.A1(n_3312),
.A2(n_2625),
.B(n_2613),
.Y(n_3711)
);

AOI21xp5_ASAP7_75t_L g3712 ( 
.A1(n_3446),
.A2(n_1821),
.B(n_1795),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3305),
.B(n_3317),
.Y(n_3713)
);

AOI22xp5_ASAP7_75t_L g3714 ( 
.A1(n_3480),
.A2(n_3013),
.B1(n_2189),
.B2(n_2197),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3294),
.B(n_1485),
.Y(n_3715)
);

INVx3_ASAP7_75t_L g3716 ( 
.A(n_3337),
.Y(n_3716)
);

HB1xp67_ASAP7_75t_L g3717 ( 
.A(n_3257),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_SL g3718 ( 
.A(n_3308),
.B(n_2189),
.Y(n_3718)
);

INVx2_ASAP7_75t_L g3719 ( 
.A(n_3318),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3334),
.B(n_3210),
.Y(n_3720)
);

BUFx6f_ASAP7_75t_L g3721 ( 
.A(n_3215),
.Y(n_3721)
);

INVx5_ASAP7_75t_L g3722 ( 
.A(n_3337),
.Y(n_3722)
);

NOR2xp67_ASAP7_75t_L g3723 ( 
.A(n_3482),
.B(n_2571),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3450),
.Y(n_3724)
);

NOR2xp33_ASAP7_75t_L g3725 ( 
.A(n_3310),
.B(n_2604),
.Y(n_3725)
);

AOI21xp5_ASAP7_75t_L g3726 ( 
.A1(n_3456),
.A2(n_1821),
.B(n_1971),
.Y(n_3726)
);

INVx2_ASAP7_75t_L g3727 ( 
.A(n_3100),
.Y(n_3727)
);

A2O1A1Ixp33_ASAP7_75t_L g3728 ( 
.A1(n_3300),
.A2(n_2629),
.B(n_2638),
.C(n_2604),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3329),
.B(n_2629),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3329),
.B(n_3013),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3308),
.B(n_3013),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3339),
.B(n_1486),
.Y(n_3732)
);

AOI21xp5_ASAP7_75t_L g3733 ( 
.A1(n_3273),
.A2(n_1821),
.B(n_1971),
.Y(n_3733)
);

AOI21xp5_ASAP7_75t_L g3734 ( 
.A1(n_3273),
.A2(n_1971),
.B(n_2131),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3363),
.B(n_3013),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3363),
.B(n_2604),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3385),
.B(n_2638),
.Y(n_3737)
);

AND2x6_ASAP7_75t_SL g3738 ( 
.A(n_3427),
.B(n_3323),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_3385),
.B(n_2638),
.Y(n_3739)
);

AOI21xp5_ASAP7_75t_L g3740 ( 
.A1(n_3444),
.A2(n_2131),
.B(n_2688),
.Y(n_3740)
);

AOI21xp5_ASAP7_75t_L g3741 ( 
.A1(n_3444),
.A2(n_2131),
.B(n_2688),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3477),
.Y(n_3742)
);

NOR2xp33_ASAP7_75t_L g3743 ( 
.A(n_3361),
.B(n_2189),
.Y(n_3743)
);

INVx3_ASAP7_75t_L g3744 ( 
.A(n_3337),
.Y(n_3744)
);

AOI21xp5_ASAP7_75t_L g3745 ( 
.A1(n_3413),
.A2(n_2197),
.B(n_2189),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3478),
.Y(n_3746)
);

NOR2xp33_ASAP7_75t_L g3747 ( 
.A(n_3260),
.B(n_2197),
.Y(n_3747)
);

AOI22xp33_ASAP7_75t_L g3748 ( 
.A1(n_3410),
.A2(n_2429),
.B1(n_2442),
.B2(n_2197),
.Y(n_3748)
);

OAI21xp5_ASAP7_75t_L g3749 ( 
.A1(n_3264),
.A2(n_1983),
.B(n_1973),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_L g3750 ( 
.A(n_3257),
.B(n_1973),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_SL g3751 ( 
.A(n_3327),
.B(n_2047),
.Y(n_3751)
);

O2A1O1Ixp5_ASAP7_75t_L g3752 ( 
.A1(n_3467),
.A2(n_1996),
.B(n_1998),
.C(n_1983),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_SL g3753 ( 
.A(n_3332),
.B(n_2047),
.Y(n_3753)
);

O2A1O1Ixp33_ASAP7_75t_L g3754 ( 
.A1(n_3313),
.A2(n_1029),
.B(n_1055),
.C(n_1027),
.Y(n_3754)
);

NOR2xp33_ASAP7_75t_L g3755 ( 
.A(n_3215),
.B(n_819),
.Y(n_3755)
);

AND2x2_ASAP7_75t_L g3756 ( 
.A(n_3302),
.B(n_1487),
.Y(n_3756)
);

INVx2_ASAP7_75t_SL g3757 ( 
.A(n_3194),
.Y(n_3757)
);

OAI22xp5_ASAP7_75t_L g3758 ( 
.A1(n_3346),
.A2(n_1996),
.B1(n_1998),
.B2(n_1983),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_3302),
.B(n_1996),
.Y(n_3759)
);

AOI21xp5_ASAP7_75t_L g3760 ( 
.A1(n_3413),
.A2(n_2109),
.B(n_2095),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3400),
.Y(n_3761)
);

AOI21xp33_ASAP7_75t_L g3762 ( 
.A1(n_3405),
.A2(n_835),
.B(n_833),
.Y(n_3762)
);

AOI21xp5_ASAP7_75t_L g3763 ( 
.A1(n_3218),
.A2(n_2109),
.B(n_2095),
.Y(n_3763)
);

INVx2_ASAP7_75t_L g3764 ( 
.A(n_3109),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3403),
.Y(n_3765)
);

NAND2x1_ASAP7_75t_L g3766 ( 
.A(n_3383),
.B(n_1998),
.Y(n_3766)
);

A2O1A1Ixp33_ASAP7_75t_L g3767 ( 
.A1(n_3408),
.A2(n_1086),
.B(n_1099),
.C(n_1055),
.Y(n_3767)
);

NAND2x1p5_ASAP7_75t_L g3768 ( 
.A(n_3424),
.B(n_2022),
.Y(n_3768)
);

AOI21xp5_ASAP7_75t_L g3769 ( 
.A1(n_3220),
.A2(n_2109),
.B(n_2095),
.Y(n_3769)
);

HB1xp67_ASAP7_75t_L g3770 ( 
.A(n_3566),
.Y(n_3770)
);

O2A1O1Ixp33_ASAP7_75t_L g3771 ( 
.A1(n_3562),
.A2(n_3472),
.B(n_3441),
.C(n_3202),
.Y(n_3771)
);

BUFx6f_ASAP7_75t_L g3772 ( 
.A(n_3591),
.Y(n_3772)
);

AOI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_3557),
.A2(n_3307),
.B(n_3426),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3631),
.B(n_3306),
.Y(n_3774)
);

NAND3xp33_ASAP7_75t_L g3775 ( 
.A(n_3484),
.B(n_3441),
.C(n_3379),
.Y(n_3775)
);

INVx4_ASAP7_75t_L g3776 ( 
.A(n_3505),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3713),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3494),
.A2(n_3426),
.B(n_3225),
.Y(n_3778)
);

NOR2xp33_ASAP7_75t_L g3779 ( 
.A(n_3483),
.B(n_3149),
.Y(n_3779)
);

NOR2xp33_ASAP7_75t_L g3780 ( 
.A(n_3492),
.B(n_3333),
.Y(n_3780)
);

NOR2xp33_ASAP7_75t_L g3781 ( 
.A(n_3487),
.B(n_3306),
.Y(n_3781)
);

INVx3_ASAP7_75t_SL g3782 ( 
.A(n_3637),
.Y(n_3782)
);

NOR3xp33_ASAP7_75t_L g3783 ( 
.A(n_3536),
.B(n_3605),
.C(n_3580),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_3761),
.B(n_3347),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3765),
.B(n_3347),
.Y(n_3785)
);

NAND3xp33_ASAP7_75t_L g3786 ( 
.A(n_3616),
.B(n_3370),
.C(n_3358),
.Y(n_3786)
);

AOI21xp5_ASAP7_75t_L g3787 ( 
.A1(n_3510),
.A2(n_3242),
.B(n_3223),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_3507),
.B(n_3394),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3680),
.Y(n_3789)
);

NAND2x1p5_ASAP7_75t_L g3790 ( 
.A(n_3701),
.B(n_3144),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_SL g3791 ( 
.A(n_3526),
.B(n_3289),
.Y(n_3791)
);

AOI21xp5_ASAP7_75t_L g3792 ( 
.A1(n_3488),
.A2(n_3425),
.B(n_3186),
.Y(n_3792)
);

AOI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_3560),
.A2(n_3445),
.B(n_3475),
.Y(n_3793)
);

BUFx4_ASAP7_75t_SL g3794 ( 
.A(n_3679),
.Y(n_3794)
);

AOI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_3511),
.A2(n_3230),
.B(n_3338),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_SL g3796 ( 
.A(n_3526),
.B(n_3370),
.Y(n_3796)
);

A2O1A1Ixp33_ASAP7_75t_L g3797 ( 
.A1(n_3613),
.A2(n_3362),
.B(n_3377),
.C(n_3373),
.Y(n_3797)
);

INVx3_ASAP7_75t_L g3798 ( 
.A(n_3505),
.Y(n_3798)
);

AOI21xp5_ASAP7_75t_L g3799 ( 
.A1(n_3512),
.A2(n_3234),
.B(n_3231),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_3619),
.B(n_3394),
.Y(n_3800)
);

O2A1O1Ixp33_ASAP7_75t_L g3801 ( 
.A1(n_3655),
.A2(n_3349),
.B(n_3340),
.C(n_1099),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_SL g3802 ( 
.A(n_3603),
.B(n_3129),
.Y(n_3802)
);

INVx3_ASAP7_75t_L g3803 ( 
.A(n_3509),
.Y(n_3803)
);

O2A1O1Ixp33_ASAP7_75t_SL g3804 ( 
.A1(n_3656),
.A2(n_3476),
.B(n_3479),
.C(n_3404),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_L g3805 ( 
.A(n_3634),
.B(n_3430),
.Y(n_3805)
);

O2A1O1Ixp33_ASAP7_75t_L g3806 ( 
.A1(n_3762),
.A2(n_1100),
.B(n_1106),
.C(n_1086),
.Y(n_3806)
);

INVxp67_ASAP7_75t_L g3807 ( 
.A(n_3600),
.Y(n_3807)
);

AOI33xp33_ASAP7_75t_L g3808 ( 
.A1(n_3715),
.A2(n_1124),
.A3(n_1106),
.B1(n_1127),
.B2(n_1107),
.B3(n_1100),
.Y(n_3808)
);

NOR2xp33_ASAP7_75t_SL g3809 ( 
.A(n_3618),
.B(n_3326),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3538),
.B(n_3430),
.Y(n_3810)
);

AND2x2_ASAP7_75t_L g3811 ( 
.A(n_3496),
.B(n_3460),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3537),
.B(n_3460),
.Y(n_3812)
);

AOI21xp5_ASAP7_75t_L g3813 ( 
.A1(n_3515),
.A2(n_3236),
.B(n_3346),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3705),
.Y(n_3814)
);

AOI21xp5_ASAP7_75t_L g3815 ( 
.A1(n_3584),
.A2(n_3351),
.B(n_3346),
.Y(n_3815)
);

AOI22xp5_ASAP7_75t_L g3816 ( 
.A1(n_3627),
.A2(n_3362),
.B1(n_3152),
.B2(n_3326),
.Y(n_3816)
);

CKINVDCx20_ASAP7_75t_R g3817 ( 
.A(n_3658),
.Y(n_3817)
);

OAI22xp5_ASAP7_75t_L g3818 ( 
.A1(n_3543),
.A2(n_3351),
.B1(n_3350),
.B2(n_3326),
.Y(n_3818)
);

AOI22xp5_ASAP7_75t_L g3819 ( 
.A1(n_3521),
.A2(n_3214),
.B1(n_3262),
.B2(n_3184),
.Y(n_3819)
);

A2O1A1Ixp33_ASAP7_75t_L g3820 ( 
.A1(n_3676),
.A2(n_3411),
.B(n_3375),
.C(n_3366),
.Y(n_3820)
);

INVx5_ASAP7_75t_L g3821 ( 
.A(n_3591),
.Y(n_3821)
);

O2A1O1Ixp33_ASAP7_75t_L g3822 ( 
.A1(n_3767),
.A2(n_1124),
.B(n_1127),
.C(n_1107),
.Y(n_3822)
);

A2O1A1Ixp33_ASAP7_75t_SL g3823 ( 
.A1(n_3747),
.A2(n_3451),
.B(n_3482),
.C(n_3180),
.Y(n_3823)
);

AOI21xp5_ASAP7_75t_L g3824 ( 
.A1(n_3689),
.A2(n_3351),
.B(n_3457),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3594),
.B(n_3117),
.Y(n_3825)
);

HB1xp67_ASAP7_75t_L g3826 ( 
.A(n_3647),
.Y(n_3826)
);

AND2x2_ASAP7_75t_L g3827 ( 
.A(n_3690),
.B(n_3131),
.Y(n_3827)
);

NOR2xp33_ASAP7_75t_R g3828 ( 
.A(n_3704),
.B(n_3144),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3720),
.B(n_3498),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3683),
.B(n_3133),
.Y(n_3830)
);

AOI21x1_ASAP7_75t_L g3831 ( 
.A1(n_3733),
.A2(n_3364),
.B(n_3352),
.Y(n_3831)
);

AOI21x1_ASAP7_75t_L g3832 ( 
.A1(n_3760),
.A2(n_3745),
.B(n_3555),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3518),
.B(n_3135),
.Y(n_3833)
);

AND2x2_ASAP7_75t_L g3834 ( 
.A(n_3756),
.B(n_3138),
.Y(n_3834)
);

AOI22xp5_ASAP7_75t_L g3835 ( 
.A1(n_3682),
.A2(n_3451),
.B1(n_3325),
.B2(n_3250),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_3491),
.B(n_3151),
.Y(n_3836)
);

AOI21xp5_ASAP7_75t_L g3837 ( 
.A1(n_3559),
.A2(n_3567),
.B(n_3522),
.Y(n_3837)
);

AOI22xp33_ASAP7_75t_L g3838 ( 
.A1(n_3645),
.A2(n_3291),
.B1(n_3322),
.B2(n_3316),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_3499),
.B(n_3500),
.Y(n_3839)
);

AOI21xp5_ASAP7_75t_L g3840 ( 
.A1(n_3579),
.A2(n_3464),
.B(n_3458),
.Y(n_3840)
);

INVx2_ASAP7_75t_L g3841 ( 
.A(n_3719),
.Y(n_3841)
);

BUFx2_ASAP7_75t_L g3842 ( 
.A(n_3686),
.Y(n_3842)
);

NAND2x1p5_ASAP7_75t_L g3843 ( 
.A(n_3701),
.B(n_3180),
.Y(n_3843)
);

AO21x1_ASAP7_75t_L g3844 ( 
.A1(n_3731),
.A2(n_3392),
.B(n_3388),
.Y(n_3844)
);

NOR2xp33_ASAP7_75t_L g3845 ( 
.A(n_3725),
.B(n_3158),
.Y(n_3845)
);

A2O1A1Ixp33_ASAP7_75t_L g3846 ( 
.A1(n_3676),
.A2(n_3284),
.B(n_3238),
.C(n_3276),
.Y(n_3846)
);

A2O1A1Ixp33_ASAP7_75t_L g3847 ( 
.A1(n_3622),
.A2(n_3293),
.B(n_3269),
.C(n_3468),
.Y(n_3847)
);

BUFx2_ASAP7_75t_L g3848 ( 
.A(n_3657),
.Y(n_3848)
);

BUFx12f_ASAP7_75t_L g3849 ( 
.A(n_3658),
.Y(n_3849)
);

AND2x4_ASAP7_75t_L g3850 ( 
.A(n_3486),
.B(n_3259),
.Y(n_3850)
);

AOI21xp5_ASAP7_75t_L g3851 ( 
.A1(n_3586),
.A2(n_3466),
.B(n_3470),
.Y(n_3851)
);

AND2x2_ASAP7_75t_L g3852 ( 
.A(n_3732),
.B(n_3164),
.Y(n_3852)
);

INVxp67_ASAP7_75t_L g3853 ( 
.A(n_3639),
.Y(n_3853)
);

OAI22xp5_ASAP7_75t_L g3854 ( 
.A1(n_3531),
.A2(n_3246),
.B1(n_3251),
.B2(n_3244),
.Y(n_3854)
);

NOR2xp33_ASAP7_75t_L g3855 ( 
.A(n_3549),
.B(n_3178),
.Y(n_3855)
);

AOI21xp5_ASAP7_75t_L g3856 ( 
.A1(n_3588),
.A2(n_3254),
.B(n_3253),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3502),
.B(n_3181),
.Y(n_3857)
);

O2A1O1Ixp33_ASAP7_75t_L g3858 ( 
.A1(n_3753),
.A2(n_1137),
.B(n_1139),
.C(n_1136),
.Y(n_3858)
);

AOI22xp5_ASAP7_75t_L g3859 ( 
.A1(n_3751),
.A2(n_3201),
.B1(n_3221),
.B2(n_3198),
.Y(n_3859)
);

NOR2xp33_ASAP7_75t_L g3860 ( 
.A(n_3553),
.B(n_3261),
.Y(n_3860)
);

NOR2xp33_ASAP7_75t_L g3861 ( 
.A(n_3578),
.B(n_3271),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_SL g3862 ( 
.A(n_3575),
.B(n_3132),
.Y(n_3862)
);

OAI21xp5_ASAP7_75t_L g3863 ( 
.A1(n_3554),
.A2(n_3485),
.B(n_3677),
.Y(n_3863)
);

AND2x2_ASAP7_75t_L g3864 ( 
.A(n_3611),
.B(n_3283),
.Y(n_3864)
);

CKINVDCx5p33_ASAP7_75t_R g3865 ( 
.A(n_3704),
.Y(n_3865)
);

A2O1A1Ixp33_ASAP7_75t_L g3866 ( 
.A1(n_3563),
.A2(n_3267),
.B(n_3270),
.C(n_3255),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3513),
.Y(n_3867)
);

AND2x4_ASAP7_75t_L g3868 ( 
.A(n_3486),
.B(n_3259),
.Y(n_3868)
);

AOI21x1_ASAP7_75t_L g3869 ( 
.A1(n_3547),
.A2(n_3281),
.B(n_3280),
.Y(n_3869)
);

INVx8_ASAP7_75t_L g3870 ( 
.A(n_3568),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_L g3871 ( 
.A(n_3506),
.B(n_3298),
.Y(n_3871)
);

AOI21xp5_ASAP7_75t_L g3872 ( 
.A1(n_3574),
.A2(n_3290),
.B(n_3288),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_SL g3873 ( 
.A(n_3527),
.B(n_3132),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3540),
.Y(n_3874)
);

AOI21xp5_ASAP7_75t_L g3875 ( 
.A1(n_3525),
.A2(n_3328),
.B(n_3314),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_3581),
.B(n_3299),
.Y(n_3876)
);

AOI21xp5_ASAP7_75t_L g3877 ( 
.A1(n_3534),
.A2(n_3694),
.B(n_3493),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_L g3878 ( 
.A(n_3508),
.B(n_3304),
.Y(n_3878)
);

INVx3_ASAP7_75t_L g3879 ( 
.A(n_3509),
.Y(n_3879)
);

AOI22xp5_ASAP7_75t_L g3880 ( 
.A1(n_3528),
.A2(n_840),
.B1(n_848),
.B2(n_839),
.Y(n_3880)
);

NOR2xp33_ASAP7_75t_L g3881 ( 
.A(n_3602),
.B(n_3319),
.Y(n_3881)
);

AOI21xp5_ASAP7_75t_L g3882 ( 
.A1(n_3635),
.A2(n_3336),
.B(n_3331),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3583),
.B(n_3330),
.Y(n_3883)
);

AOI21xp5_ASAP7_75t_L g3884 ( 
.A1(n_3597),
.A2(n_3357),
.B(n_3354),
.Y(n_3884)
);

AND2x2_ASAP7_75t_L g3885 ( 
.A(n_3709),
.B(n_3717),
.Y(n_3885)
);

INVx2_ASAP7_75t_L g3886 ( 
.A(n_3551),
.Y(n_3886)
);

BUFx6f_ASAP7_75t_L g3887 ( 
.A(n_3591),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_SL g3888 ( 
.A(n_3678),
.B(n_3132),
.Y(n_3888)
);

AOI21xp5_ASAP7_75t_L g3889 ( 
.A1(n_3599),
.A2(n_3365),
.B(n_3359),
.Y(n_3889)
);

AND2x4_ASAP7_75t_L g3890 ( 
.A(n_3716),
.B(n_3275),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_L g3891 ( 
.A(n_3587),
.B(n_3348),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_3530),
.B(n_3355),
.Y(n_3892)
);

NOR2xp33_ASAP7_75t_L g3893 ( 
.A(n_3571),
.B(n_3367),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_L g3894 ( 
.A(n_3533),
.B(n_3390),
.Y(n_3894)
);

NOR2xp33_ASAP7_75t_L g3895 ( 
.A(n_3738),
.B(n_3275),
.Y(n_3895)
);

AOI22xp33_ASAP7_75t_L g3896 ( 
.A1(n_3503),
.A2(n_3755),
.B1(n_3716),
.B2(n_3744),
.Y(n_3896)
);

NOR2xp33_ASAP7_75t_SL g3897 ( 
.A(n_3532),
.B(n_3404),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3544),
.B(n_3545),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_L g3899 ( 
.A(n_3550),
.B(n_3368),
.Y(n_3899)
);

OAI22xp5_ASAP7_75t_L g3900 ( 
.A1(n_3695),
.A2(n_3389),
.B1(n_3391),
.B2(n_3369),
.Y(n_3900)
);

AOI21xp5_ASAP7_75t_L g3901 ( 
.A1(n_3523),
.A2(n_3245),
.B(n_3132),
.Y(n_3901)
);

AOI21xp5_ASAP7_75t_L g3902 ( 
.A1(n_3565),
.A2(n_3245),
.B(n_3132),
.Y(n_3902)
);

AOI21xp5_ASAP7_75t_L g3903 ( 
.A1(n_3556),
.A2(n_3245),
.B(n_3132),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3648),
.B(n_3407),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3490),
.Y(n_3905)
);

AOI21xp5_ASAP7_75t_L g3906 ( 
.A1(n_3734),
.A2(n_3245),
.B(n_3479),
.Y(n_3906)
);

INVx2_ASAP7_75t_L g3907 ( 
.A(n_3593),
.Y(n_3907)
);

AOI21xp5_ASAP7_75t_L g3908 ( 
.A1(n_3610),
.A2(n_3245),
.B(n_3407),
.Y(n_3908)
);

AND2x4_ASAP7_75t_L g3909 ( 
.A(n_3744),
.B(n_3414),
.Y(n_3909)
);

INVx2_ASAP7_75t_L g3910 ( 
.A(n_3621),
.Y(n_3910)
);

CKINVDCx20_ASAP7_75t_R g3911 ( 
.A(n_3669),
.Y(n_3911)
);

NOR2xp33_ASAP7_75t_L g3912 ( 
.A(n_3666),
.B(n_3414),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_L g3913 ( 
.A(n_3663),
.B(n_853),
.Y(n_3913)
);

OAI22xp5_ASAP7_75t_L g3914 ( 
.A1(n_3743),
.A2(n_3585),
.B1(n_3722),
.B2(n_3497),
.Y(n_3914)
);

NOR2xp33_ASAP7_75t_L g3915 ( 
.A(n_3709),
.B(n_854),
.Y(n_3915)
);

AOI221xp5_ASAP7_75t_L g3916 ( 
.A1(n_3670),
.A2(n_870),
.B1(n_875),
.B2(n_872),
.C(n_868),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_L g3917 ( 
.A(n_3612),
.B(n_877),
.Y(n_3917)
);

OR2x2_ASAP7_75t_L g3918 ( 
.A(n_3659),
.B(n_1488),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3641),
.Y(n_3919)
);

NOR2xp33_ASAP7_75t_L g3920 ( 
.A(n_3721),
.B(n_880),
.Y(n_3920)
);

CKINVDCx16_ASAP7_75t_R g3921 ( 
.A(n_3489),
.Y(n_3921)
);

AOI21xp5_ASAP7_75t_L g3922 ( 
.A1(n_3692),
.A2(n_3245),
.B(n_2109),
.Y(n_3922)
);

AND2x2_ASAP7_75t_SL g3923 ( 
.A(n_3519),
.B(n_858),
.Y(n_3923)
);

AOI21x1_ASAP7_75t_L g3924 ( 
.A1(n_3711),
.A2(n_1413),
.B(n_1409),
.Y(n_3924)
);

NAND2xp5_ASAP7_75t_L g3925 ( 
.A(n_3614),
.B(n_883),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_3667),
.Y(n_3926)
);

OAI21xp5_ASAP7_75t_L g3927 ( 
.A1(n_3606),
.A2(n_2030),
.B(n_2022),
.Y(n_3927)
);

AOI21xp5_ASAP7_75t_L g3928 ( 
.A1(n_3707),
.A2(n_2109),
.B(n_2095),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3654),
.B(n_889),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_SL g3930 ( 
.A(n_3722),
.B(n_890),
.Y(n_3930)
);

INVx2_ASAP7_75t_SL g3931 ( 
.A(n_3628),
.Y(n_3931)
);

O2A1O1Ixp5_ASAP7_75t_L g3932 ( 
.A1(n_3514),
.A2(n_1137),
.B(n_1139),
.C(n_1136),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3671),
.B(n_892),
.Y(n_3933)
);

NOR2xp33_ASAP7_75t_L g3934 ( 
.A(n_3721),
.B(n_896),
.Y(n_3934)
);

AOI21xp5_ASAP7_75t_L g3935 ( 
.A1(n_3604),
.A2(n_2095),
.B(n_2030),
.Y(n_3935)
);

HB1xp67_ASAP7_75t_L g3936 ( 
.A(n_3721),
.Y(n_3936)
);

AOI21xp5_ASAP7_75t_L g3937 ( 
.A1(n_3542),
.A2(n_3608),
.B(n_3529),
.Y(n_3937)
);

NOR2x1_ASAP7_75t_L g3938 ( 
.A(n_3568),
.B(n_1936),
.Y(n_3938)
);

AOI21xp5_ASAP7_75t_L g3939 ( 
.A1(n_3561),
.A2(n_2030),
.B(n_2022),
.Y(n_3939)
);

BUFx2_ASAP7_75t_L g3940 ( 
.A(n_3607),
.Y(n_3940)
);

AOI21x1_ASAP7_75t_L g3941 ( 
.A1(n_3504),
.A2(n_1490),
.B(n_1489),
.Y(n_3941)
);

CKINVDCx5p33_ASAP7_75t_R g3942 ( 
.A(n_3693),
.Y(n_3942)
);

AO22x1_ASAP7_75t_L g3943 ( 
.A1(n_3722),
.A2(n_897),
.B1(n_900),
.B2(n_899),
.Y(n_3943)
);

A2O1A1Ixp33_ASAP7_75t_L g3944 ( 
.A1(n_3606),
.A2(n_3754),
.B(n_3730),
.C(n_3535),
.Y(n_3944)
);

AOI21xp5_ASAP7_75t_L g3945 ( 
.A1(n_3726),
.A2(n_2092),
.B(n_2069),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_SL g3946 ( 
.A(n_3698),
.B(n_903),
.Y(n_3946)
);

INVx3_ASAP7_75t_SL g3947 ( 
.A(n_3757),
.Y(n_3947)
);

OAI22xp5_ASAP7_75t_L g3948 ( 
.A1(n_3585),
.A2(n_904),
.B1(n_911),
.B2(n_910),
.Y(n_3948)
);

CKINVDCx11_ASAP7_75t_R g3949 ( 
.A(n_3607),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_3495),
.B(n_912),
.Y(n_3950)
);

O2A1O1Ixp33_ASAP7_75t_L g3951 ( 
.A1(n_3718),
.A2(n_1149),
.B(n_1158),
.C(n_1143),
.Y(n_3951)
);

O2A1O1Ixp5_ASAP7_75t_L g3952 ( 
.A1(n_3501),
.A2(n_1149),
.B(n_1158),
.C(n_1143),
.Y(n_3952)
);

OR2x2_ASAP7_75t_L g3953 ( 
.A(n_3517),
.B(n_1494),
.Y(n_3953)
);

INVx3_ASAP7_75t_L g3954 ( 
.A(n_3568),
.Y(n_3954)
);

INVx2_ASAP7_75t_L g3955 ( 
.A(n_3727),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3520),
.B(n_914),
.Y(n_3956)
);

AOI21x1_ASAP7_75t_L g3957 ( 
.A1(n_3652),
.A2(n_1498),
.B(n_1496),
.Y(n_3957)
);

OAI21xp33_ASAP7_75t_L g3958 ( 
.A1(n_3596),
.A2(n_917),
.B(n_915),
.Y(n_3958)
);

AOI21xp5_ASAP7_75t_L g3959 ( 
.A1(n_3763),
.A2(n_2092),
.B(n_2069),
.Y(n_3959)
);

NOR2xp33_ASAP7_75t_L g3960 ( 
.A(n_3764),
.B(n_920),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3524),
.B(n_921),
.Y(n_3961)
);

NAND2x1p5_ASAP7_75t_L g3962 ( 
.A(n_3696),
.B(n_2069),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_L g3963 ( 
.A(n_3539),
.B(n_922),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_SL g3964 ( 
.A(n_3698),
.B(n_925),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_3546),
.B(n_926),
.Y(n_3965)
);

AOI21xp5_ASAP7_75t_L g3966 ( 
.A1(n_3769),
.A2(n_2092),
.B(n_2026),
.Y(n_3966)
);

O2A1O1Ixp5_ASAP7_75t_L g3967 ( 
.A1(n_3624),
.A2(n_1170),
.B(n_1168),
.C(n_941),
.Y(n_3967)
);

NOR2xp33_ASAP7_75t_L g3968 ( 
.A(n_3687),
.B(n_927),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3548),
.B(n_3558),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_L g3970 ( 
.A(n_3569),
.B(n_928),
.Y(n_3970)
);

NOR2x1p5_ASAP7_75t_L g3971 ( 
.A(n_3516),
.B(n_1499),
.Y(n_3971)
);

O2A1O1Ixp33_ASAP7_75t_L g3972 ( 
.A1(n_3640),
.A2(n_1170),
.B(n_1168),
.C(n_945),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3572),
.B(n_931),
.Y(n_3973)
);

AND2x4_ASAP7_75t_L g3974 ( 
.A(n_3585),
.B(n_1936),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_3573),
.B(n_933),
.Y(n_3975)
);

AOI21xp5_ASAP7_75t_L g3976 ( 
.A1(n_3601),
.A2(n_2026),
.B(n_1991),
.Y(n_3976)
);

AOI21xp5_ASAP7_75t_L g3977 ( 
.A1(n_3633),
.A2(n_2032),
.B(n_2026),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3576),
.Y(n_3978)
);

AOI22x1_ASAP7_75t_SL g3979 ( 
.A1(n_3516),
.A2(n_934),
.B1(n_939),
.B2(n_937),
.Y(n_3979)
);

OAI21xp5_ASAP7_75t_L g3980 ( 
.A1(n_3577),
.A2(n_1942),
.B(n_1936),
.Y(n_3980)
);

A2O1A1Ixp33_ASAP7_75t_L g3981 ( 
.A1(n_3735),
.A2(n_945),
.B(n_982),
.C(n_858),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_L g3982 ( 
.A(n_3582),
.B(n_942),
.Y(n_3982)
);

AOI21x1_ASAP7_75t_L g3983 ( 
.A1(n_3708),
.A2(n_1507),
.B(n_1503),
.Y(n_3983)
);

OAI21xp33_ASAP7_75t_L g3984 ( 
.A1(n_3742),
.A2(n_946),
.B(n_944),
.Y(n_3984)
);

NAND3xp33_ASAP7_75t_L g3985 ( 
.A(n_3714),
.B(n_949),
.C(n_947),
.Y(n_3985)
);

BUFx3_ASAP7_75t_L g3986 ( 
.A(n_3607),
.Y(n_3986)
);

HB1xp67_ASAP7_75t_L g3987 ( 
.A(n_3590),
.Y(n_3987)
);

AOI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_3729),
.A2(n_2032),
.B(n_2026),
.Y(n_3988)
);

A2O1A1Ixp33_ASAP7_75t_L g3989 ( 
.A1(n_3746),
.A2(n_1098),
.B(n_1105),
.C(n_982),
.Y(n_3989)
);

AND2x4_ASAP7_75t_L g3990 ( 
.A(n_3570),
.B(n_1942),
.Y(n_3990)
);

AOI21xp5_ASAP7_75t_L g3991 ( 
.A1(n_3661),
.A2(n_2035),
.B(n_2032),
.Y(n_3991)
);

NOR2xp33_ASAP7_75t_SL g3992 ( 
.A(n_3592),
.B(n_952),
.Y(n_3992)
);

AND2x4_ASAP7_75t_L g3993 ( 
.A(n_3570),
.B(n_1942),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3598),
.Y(n_3994)
);

O2A1O1Ixp5_ASAP7_75t_L g3995 ( 
.A1(n_3752),
.A2(n_3758),
.B(n_3638),
.C(n_3625),
.Y(n_3995)
);

AND2x2_ASAP7_75t_L g3996 ( 
.A(n_3623),
.B(n_1508),
.Y(n_3996)
);

NOR2xp67_ASAP7_75t_L g3997 ( 
.A(n_3660),
.B(n_543),
.Y(n_3997)
);

BUFx6f_ASAP7_75t_L g3998 ( 
.A(n_3617),
.Y(n_3998)
);

OAI22xp5_ASAP7_75t_L g3999 ( 
.A1(n_3748),
.A2(n_960),
.B1(n_962),
.B2(n_959),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3632),
.B(n_963),
.Y(n_4000)
);

AND2x4_ASAP7_75t_L g4001 ( 
.A(n_3646),
.B(n_1510),
.Y(n_4001)
);

NOR2x1_ASAP7_75t_L g4002 ( 
.A(n_3750),
.B(n_1512),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3724),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3684),
.Y(n_4004)
);

INVx2_ASAP7_75t_L g4005 ( 
.A(n_3698),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_L g4006 ( 
.A(n_3552),
.B(n_964),
.Y(n_4006)
);

AOI21xp5_ASAP7_75t_L g4007 ( 
.A1(n_3697),
.A2(n_2035),
.B(n_2032),
.Y(n_4007)
);

NOR2xp33_ASAP7_75t_SL g4008 ( 
.A(n_3617),
.B(n_965),
.Y(n_4008)
);

INVx2_ASAP7_75t_L g4009 ( 
.A(n_3698),
.Y(n_4009)
);

INVx2_ASAP7_75t_L g4010 ( 
.A(n_3698),
.Y(n_4010)
);

OAI22xp5_ASAP7_75t_L g4011 ( 
.A1(n_3736),
.A2(n_970),
.B1(n_971),
.B2(n_967),
.Y(n_4011)
);

INVx1_ASAP7_75t_SL g4012 ( 
.A(n_3617),
.Y(n_4012)
);

O2A1O1Ixp33_ASAP7_75t_L g4013 ( 
.A1(n_3630),
.A2(n_1105),
.B(n_1130),
.C(n_1098),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3685),
.Y(n_4014)
);

BUFx3_ASAP7_75t_L g4015 ( 
.A(n_3629),
.Y(n_4015)
);

AND2x2_ASAP7_75t_L g4016 ( 
.A(n_3759),
.B(n_1518),
.Y(n_4016)
);

AO32x1_ASAP7_75t_L g4017 ( 
.A1(n_3651),
.A2(n_1146),
.A3(n_1142),
.B1(n_1130),
.B2(n_1523),
.Y(n_4017)
);

AOI22xp5_ASAP7_75t_L g4018 ( 
.A1(n_3649),
.A2(n_973),
.B1(n_976),
.B2(n_974),
.Y(n_4018)
);

INVx2_ASAP7_75t_L g4019 ( 
.A(n_3564),
.Y(n_4019)
);

AOI21xp5_ASAP7_75t_L g4020 ( 
.A1(n_3699),
.A2(n_2036),
.B(n_2035),
.Y(n_4020)
);

A2O1A1Ixp33_ASAP7_75t_L g4021 ( 
.A1(n_3737),
.A2(n_1146),
.B(n_1142),
.C(n_979),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3644),
.B(n_3642),
.Y(n_4022)
);

NAND2x1p5_ASAP7_75t_L g4023 ( 
.A(n_3821),
.B(n_3660),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3898),
.B(n_3662),
.Y(n_4024)
);

INVx3_ASAP7_75t_L g4025 ( 
.A(n_3890),
.Y(n_4025)
);

AND2x4_ASAP7_75t_L g4026 ( 
.A(n_3954),
.B(n_3629),
.Y(n_4026)
);

OAI22xp5_ASAP7_75t_L g4027 ( 
.A1(n_3775),
.A2(n_3739),
.B1(n_3691),
.B2(n_3541),
.Y(n_4027)
);

AND2x4_ASAP7_75t_L g4028 ( 
.A(n_3954),
.B(n_3629),
.Y(n_4028)
);

OR2x2_ASAP7_75t_L g4029 ( 
.A(n_3770),
.B(n_3681),
.Y(n_4029)
);

O2A1O1Ixp5_ASAP7_75t_L g4030 ( 
.A1(n_3863),
.A2(n_3749),
.B(n_3615),
.C(n_3688),
.Y(n_4030)
);

AOI22x1_ASAP7_75t_L g4031 ( 
.A1(n_3971),
.A2(n_3768),
.B1(n_3595),
.B2(n_3589),
.Y(n_4031)
);

BUFx6f_ASAP7_75t_L g4032 ( 
.A(n_3949),
.Y(n_4032)
);

INVx3_ASAP7_75t_L g4033 ( 
.A(n_3890),
.Y(n_4033)
);

OAI22xp5_ASAP7_75t_L g4034 ( 
.A1(n_3816),
.A2(n_3675),
.B1(n_3626),
.B2(n_3728),
.Y(n_4034)
);

OAI21x1_ASAP7_75t_L g4035 ( 
.A1(n_3832),
.A2(n_3609),
.B(n_3740),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_L g4036 ( 
.A(n_3839),
.B(n_3636),
.Y(n_4036)
);

CKINVDCx5p33_ASAP7_75t_R g4037 ( 
.A(n_3865),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_3987),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3905),
.Y(n_4039)
);

NOR2xp33_ASAP7_75t_L g4040 ( 
.A(n_3780),
.B(n_3636),
.Y(n_4040)
);

OAI21xp5_ASAP7_75t_L g4041 ( 
.A1(n_3783),
.A2(n_3797),
.B(n_3952),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_L g4042 ( 
.A(n_4019),
.B(n_3864),
.Y(n_4042)
);

BUFx3_ASAP7_75t_L g4043 ( 
.A(n_3842),
.Y(n_4043)
);

OAI21x1_ASAP7_75t_L g4044 ( 
.A1(n_3941),
.A2(n_3741),
.B(n_3620),
.Y(n_4044)
);

AOI21xp5_ASAP7_75t_L g4045 ( 
.A1(n_3877),
.A2(n_3653),
.B(n_3702),
.Y(n_4045)
);

OAI21x1_ASAP7_75t_L g4046 ( 
.A1(n_3837),
.A2(n_3643),
.B(n_3700),
.Y(n_4046)
);

AOI21x1_ASAP7_75t_L g4047 ( 
.A1(n_3906),
.A2(n_3723),
.B(n_3650),
.Y(n_4047)
);

OAI21x1_ASAP7_75t_L g4048 ( 
.A1(n_3924),
.A2(n_3710),
.B(n_3706),
.Y(n_4048)
);

AO21x1_ASAP7_75t_L g4049 ( 
.A1(n_3791),
.A2(n_3673),
.B(n_3766),
.Y(n_4049)
);

BUFx3_ASAP7_75t_L g4050 ( 
.A(n_3848),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_L g4051 ( 
.A(n_3777),
.B(n_3636),
.Y(n_4051)
);

AOI22xp5_ASAP7_75t_L g4052 ( 
.A1(n_3802),
.A2(n_980),
.B1(n_983),
.B2(n_981),
.Y(n_4052)
);

OAI21x1_ASAP7_75t_L g4053 ( 
.A1(n_3957),
.A2(n_3983),
.B(n_3988),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_L g4054 ( 
.A(n_3829),
.B(n_3674),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_SL g4055 ( 
.A(n_3923),
.B(n_3723),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_SL g4056 ( 
.A(n_3816),
.B(n_3674),
.Y(n_4056)
);

OAI21xp5_ASAP7_75t_L g4057 ( 
.A1(n_3820),
.A2(n_3712),
.B(n_3703),
.Y(n_4057)
);

HB1xp67_ASAP7_75t_L g4058 ( 
.A(n_3826),
.Y(n_4058)
);

OAI21xp5_ASAP7_75t_L g4059 ( 
.A1(n_3824),
.A2(n_3932),
.B(n_3771),
.Y(n_4059)
);

INVx1_ASAP7_75t_SL g4060 ( 
.A(n_3834),
.Y(n_4060)
);

AOI221xp5_ASAP7_75t_SL g4061 ( 
.A1(n_3806),
.A2(n_1528),
.B1(n_1530),
.B2(n_1526),
.C(n_1524),
.Y(n_4061)
);

NAND3x1_ASAP7_75t_L g4062 ( 
.A(n_3819),
.B(n_1532),
.C(n_1531),
.Y(n_4062)
);

INVx2_ASAP7_75t_L g4063 ( 
.A(n_3789),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_3774),
.B(n_3674),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3827),
.B(n_984),
.Y(n_4065)
);

OR2x6_ASAP7_75t_L g4066 ( 
.A(n_3870),
.B(n_1533),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_SL g4067 ( 
.A(n_3809),
.B(n_3845),
.Y(n_4067)
);

CKINVDCx6p67_ASAP7_75t_R g4068 ( 
.A(n_3849),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_3784),
.B(n_986),
.Y(n_4069)
);

INVxp67_ASAP7_75t_L g4070 ( 
.A(n_3781),
.Y(n_4070)
);

OAI21x1_ASAP7_75t_L g4071 ( 
.A1(n_3778),
.A2(n_3991),
.B(n_3959),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_3978),
.Y(n_4072)
);

AO21x2_ASAP7_75t_L g4073 ( 
.A1(n_3773),
.A2(n_3665),
.B(n_3664),
.Y(n_4073)
);

AND2x4_ASAP7_75t_L g4074 ( 
.A(n_3885),
.B(n_544),
.Y(n_4074)
);

OAI21x1_ASAP7_75t_SL g4075 ( 
.A1(n_3844),
.A2(n_3672),
.B(n_3668),
.Y(n_4075)
);

AOI21xp5_ASAP7_75t_L g4076 ( 
.A1(n_3903),
.A2(n_2036),
.B(n_2035),
.Y(n_4076)
);

CKINVDCx5p33_ASAP7_75t_R g4077 ( 
.A(n_3794),
.Y(n_4077)
);

NOR2xp33_ASAP7_75t_L g4078 ( 
.A(n_3893),
.B(n_987),
.Y(n_4078)
);

AOI21xp5_ASAP7_75t_L g4079 ( 
.A1(n_3882),
.A2(n_2050),
.B(n_2036),
.Y(n_4079)
);

BUFx6f_ASAP7_75t_L g4080 ( 
.A(n_3772),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_3994),
.Y(n_4081)
);

BUFx6f_ASAP7_75t_L g4082 ( 
.A(n_3772),
.Y(n_4082)
);

A2O1A1Ixp33_ASAP7_75t_L g4083 ( 
.A1(n_3779),
.A2(n_1536),
.B(n_1537),
.C(n_1535),
.Y(n_4083)
);

OA22x2_ASAP7_75t_L g4084 ( 
.A1(n_3796),
.A2(n_989),
.B1(n_990),
.B2(n_988),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_3841),
.Y(n_4085)
);

INVx2_ASAP7_75t_L g4086 ( 
.A(n_3867),
.Y(n_4086)
);

CKINVDCx9p33_ASAP7_75t_R g4087 ( 
.A(n_3895),
.Y(n_4087)
);

CKINVDCx20_ASAP7_75t_R g4088 ( 
.A(n_3817),
.Y(n_4088)
);

AOI21xp5_ASAP7_75t_L g4089 ( 
.A1(n_3922),
.A2(n_2050),
.B(n_2036),
.Y(n_4089)
);

NAND2xp33_ASAP7_75t_L g4090 ( 
.A(n_3942),
.B(n_997),
.Y(n_4090)
);

OAI21x1_ASAP7_75t_L g4091 ( 
.A1(n_3795),
.A2(n_1702),
.B(n_1540),
.Y(n_4091)
);

INVx1_ASAP7_75t_SL g4092 ( 
.A(n_3828),
.Y(n_4092)
);

AND2x6_ASAP7_75t_SL g4093 ( 
.A(n_3920),
.B(n_1539),
.Y(n_4093)
);

OAI21x1_ASAP7_75t_L g4094 ( 
.A1(n_3945),
.A2(n_1545),
.B(n_1541),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_3785),
.B(n_992),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_4003),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3830),
.B(n_993),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_3969),
.Y(n_4098)
);

INVx2_ASAP7_75t_L g4099 ( 
.A(n_3874),
.Y(n_4099)
);

INVx2_ASAP7_75t_SL g4100 ( 
.A(n_3921),
.Y(n_4100)
);

OAI22x1_ASAP7_75t_L g4101 ( 
.A1(n_3880),
.A2(n_996),
.B1(n_1002),
.B2(n_995),
.Y(n_4101)
);

INVx5_ASAP7_75t_L g4102 ( 
.A(n_3821),
.Y(n_4102)
);

AOI21xp5_ASAP7_75t_L g4103 ( 
.A1(n_3792),
.A2(n_2053),
.B(n_2050),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_3861),
.B(n_1003),
.Y(n_4104)
);

OAI22xp5_ASAP7_75t_L g4105 ( 
.A1(n_3800),
.A2(n_1007),
.B1(n_1008),
.B2(n_1006),
.Y(n_4105)
);

OAI21x1_ASAP7_75t_L g4106 ( 
.A1(n_3937),
.A2(n_1549),
.B(n_1547),
.Y(n_4106)
);

AOI21xp5_ASAP7_75t_SL g4107 ( 
.A1(n_3866),
.A2(n_2053),
.B(n_2050),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_SL g4108 ( 
.A(n_3896),
.B(n_1552),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_SL g4109 ( 
.A(n_3855),
.B(n_1557),
.Y(n_4109)
);

AOI31xp67_ASAP7_75t_L g4110 ( 
.A1(n_3946),
.A2(n_2248),
.A3(n_2259),
.B(n_2254),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_3814),
.Y(n_4111)
);

OAI21xp5_ASAP7_75t_L g4112 ( 
.A1(n_4021),
.A2(n_3944),
.B(n_3968),
.Y(n_4112)
);

OAI21x1_ASAP7_75t_L g4113 ( 
.A1(n_3799),
.A2(n_1564),
.B(n_1563),
.Y(n_4113)
);

OAI22xp5_ASAP7_75t_L g4114 ( 
.A1(n_3805),
.A2(n_1013),
.B1(n_1016),
.B2(n_1012),
.Y(n_4114)
);

AOI21xp5_ASAP7_75t_L g4115 ( 
.A1(n_3875),
.A2(n_2059),
.B(n_2053),
.Y(n_4115)
);

AOI21xp5_ASAP7_75t_L g4116 ( 
.A1(n_3815),
.A2(n_2059),
.B(n_2053),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_3886),
.Y(n_4117)
);

AND2x2_ASAP7_75t_L g4118 ( 
.A(n_3811),
.B(n_1566),
.Y(n_4118)
);

AOI221xp5_ASAP7_75t_SL g4119 ( 
.A1(n_3822),
.A2(n_1571),
.B1(n_1572),
.B2(n_1568),
.C(n_1567),
.Y(n_4119)
);

AND2x2_ASAP7_75t_L g4120 ( 
.A(n_3852),
.B(n_1573),
.Y(n_4120)
);

OAI21xp5_ASAP7_75t_L g4121 ( 
.A1(n_3880),
.A2(n_1578),
.B(n_1575),
.Y(n_4121)
);

AO31x2_ASAP7_75t_L g4122 ( 
.A1(n_3976),
.A2(n_1579),
.A3(n_1582),
.B(n_1580),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_3892),
.B(n_1021),
.Y(n_4123)
);

OAI21xp5_ASAP7_75t_L g4124 ( 
.A1(n_3840),
.A2(n_1024),
.B(n_1022),
.Y(n_4124)
);

AO31x2_ASAP7_75t_L g4125 ( 
.A1(n_3977),
.A2(n_2248),
.A3(n_2259),
.B(n_2254),
.Y(n_4125)
);

OAI21x1_ASAP7_75t_L g4126 ( 
.A1(n_3869),
.A2(n_2266),
.B(n_2265),
.Y(n_4126)
);

OAI21x1_ASAP7_75t_L g4127 ( 
.A1(n_3966),
.A2(n_2266),
.B(n_2265),
.Y(n_4127)
);

OR2x6_ASAP7_75t_L g4128 ( 
.A(n_3870),
.B(n_2059),
.Y(n_4128)
);

INVx2_ASAP7_75t_L g4129 ( 
.A(n_3907),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3910),
.Y(n_4130)
);

OAI21xp5_ASAP7_75t_L g4131 ( 
.A1(n_3917),
.A2(n_1028),
.B(n_1025),
.Y(n_4131)
);

INVx3_ASAP7_75t_L g4132 ( 
.A(n_3909),
.Y(n_4132)
);

OAI21x1_ASAP7_75t_L g4133 ( 
.A1(n_3908),
.A2(n_2275),
.B(n_2267),
.Y(n_4133)
);

OAI21x1_ASAP7_75t_L g4134 ( 
.A1(n_3884),
.A2(n_2275),
.B(n_2267),
.Y(n_4134)
);

AOI21x1_ASAP7_75t_L g4135 ( 
.A1(n_3793),
.A2(n_2291),
.B(n_2290),
.Y(n_4135)
);

AOI21x1_ASAP7_75t_L g4136 ( 
.A1(n_3939),
.A2(n_2291),
.B(n_2290),
.Y(n_4136)
);

OAI21x1_ASAP7_75t_L g4137 ( 
.A1(n_3889),
.A2(n_2293),
.B(n_2144),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_3894),
.B(n_1030),
.Y(n_4138)
);

INVx2_ASAP7_75t_L g4139 ( 
.A(n_3919),
.Y(n_4139)
);

BUFx6f_ASAP7_75t_L g4140 ( 
.A(n_3772),
.Y(n_4140)
);

AOI22xp5_ASAP7_75t_L g4141 ( 
.A1(n_3818),
.A2(n_1032),
.B1(n_1039),
.B2(n_1033),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_3825),
.B(n_1040),
.Y(n_4142)
);

OAI22xp5_ASAP7_75t_L g4143 ( 
.A1(n_3812),
.A2(n_1044),
.B1(n_1046),
.B2(n_1041),
.Y(n_4143)
);

OAI21x1_ASAP7_75t_L g4144 ( 
.A1(n_3901),
.A2(n_2293),
.B(n_2144),
.Y(n_4144)
);

OAI21xp5_ASAP7_75t_L g4145 ( 
.A1(n_3925),
.A2(n_1050),
.B(n_1049),
.Y(n_4145)
);

OAI22xp5_ASAP7_75t_L g4146 ( 
.A1(n_3860),
.A2(n_3835),
.B1(n_3786),
.B2(n_3810),
.Y(n_4146)
);

AOI21xp5_ASAP7_75t_L g4147 ( 
.A1(n_3856),
.A2(n_3813),
.B(n_3851),
.Y(n_4147)
);

AOI21xp5_ASAP7_75t_L g4148 ( 
.A1(n_3872),
.A2(n_2071),
.B(n_2059),
.Y(n_4148)
);

INVx3_ASAP7_75t_L g4149 ( 
.A(n_3909),
.Y(n_4149)
);

OAI21x1_ASAP7_75t_L g4150 ( 
.A1(n_3902),
.A2(n_2144),
.B(n_2133),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_3926),
.Y(n_4151)
);

NOR2xp33_ASAP7_75t_L g4152 ( 
.A(n_3911),
.B(n_1051),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_3857),
.B(n_1053),
.Y(n_4153)
);

A2O1A1Ixp33_ASAP7_75t_L g4154 ( 
.A1(n_3808),
.A2(n_1072),
.B(n_1091),
.C(n_1060),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_3871),
.B(n_3876),
.Y(n_4155)
);

OAI21x1_ASAP7_75t_SL g4156 ( 
.A1(n_3914),
.A2(n_3951),
.B(n_3927),
.Y(n_4156)
);

OAI21x1_ASAP7_75t_L g4157 ( 
.A1(n_3787),
.A2(n_2151),
.B(n_2133),
.Y(n_4157)
);

INVxp67_ASAP7_75t_L g4158 ( 
.A(n_3913),
.Y(n_4158)
);

NOR2xp33_ASAP7_75t_L g4159 ( 
.A(n_3912),
.B(n_1054),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_3955),
.Y(n_4160)
);

HB1xp67_ASAP7_75t_L g4161 ( 
.A(n_3807),
.Y(n_4161)
);

AO31x2_ASAP7_75t_L g4162 ( 
.A1(n_3928),
.A2(n_863),
.A3(n_1880),
.B(n_548),
.Y(n_4162)
);

AO31x2_ASAP7_75t_L g4163 ( 
.A1(n_4005),
.A2(n_863),
.A3(n_1880),
.B(n_549),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_3953),
.Y(n_4164)
);

OAI21xp5_ASAP7_75t_L g4165 ( 
.A1(n_3788),
.A2(n_1058),
.B(n_1056),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_L g4166 ( 
.A(n_3878),
.B(n_1059),
.Y(n_4166)
);

OAI21xp5_ASAP7_75t_L g4167 ( 
.A1(n_3929),
.A2(n_1063),
.B(n_1062),
.Y(n_4167)
);

AO31x2_ASAP7_75t_L g4168 ( 
.A1(n_4009),
.A2(n_863),
.A3(n_1880),
.B(n_550),
.Y(n_4168)
);

OAI21x1_ASAP7_75t_L g4169 ( 
.A1(n_3935),
.A2(n_2151),
.B(n_2133),
.Y(n_4169)
);

AO31x2_ASAP7_75t_L g4170 ( 
.A1(n_4010),
.A2(n_863),
.A3(n_551),
.B(n_559),
.Y(n_4170)
);

AOI22xp33_ASAP7_75t_L g4171 ( 
.A1(n_3881),
.A2(n_1065),
.B1(n_1066),
.B2(n_1064),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_L g4172 ( 
.A(n_3899),
.B(n_1067),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_3836),
.B(n_1068),
.Y(n_4173)
);

NAND2xp5_ASAP7_75t_L g4174 ( 
.A(n_3883),
.B(n_1073),
.Y(n_4174)
);

AOI21xp5_ASAP7_75t_L g4175 ( 
.A1(n_3804),
.A2(n_2104),
.B(n_2071),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_3996),
.Y(n_4176)
);

INVx3_ASAP7_75t_L g4177 ( 
.A(n_3870),
.Y(n_4177)
);

OAI21x1_ASAP7_75t_L g4178 ( 
.A1(n_4007),
.A2(n_2168),
.B(n_2151),
.Y(n_4178)
);

AND2x4_ASAP7_75t_L g4179 ( 
.A(n_3938),
.B(n_546),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_3891),
.B(n_1074),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_L g4181 ( 
.A(n_4004),
.B(n_1076),
.Y(n_4181)
);

AND2x6_ASAP7_75t_SL g4182 ( 
.A(n_3934),
.B(n_1077),
.Y(n_4182)
);

OA21x2_ASAP7_75t_L g4183 ( 
.A1(n_3995),
.A2(n_1080),
.B(n_1078),
.Y(n_4183)
);

AOI21xp5_ASAP7_75t_L g4184 ( 
.A1(n_4022),
.A2(n_2104),
.B(n_2071),
.Y(n_4184)
);

AND3x4_ASAP7_75t_L g4185 ( 
.A(n_3850),
.B(n_1092),
.C(n_1084),
.Y(n_4185)
);

AOI21xp5_ASAP7_75t_L g4186 ( 
.A1(n_3964),
.A2(n_2104),
.B(n_2071),
.Y(n_4186)
);

NOR2xp67_ASAP7_75t_SL g4187 ( 
.A(n_3985),
.B(n_1093),
.Y(n_4187)
);

OAI21xp5_ASAP7_75t_L g4188 ( 
.A1(n_4006),
.A2(n_1096),
.B(n_1094),
.Y(n_4188)
);

OAI21x1_ASAP7_75t_L g4189 ( 
.A1(n_4020),
.A2(n_2185),
.B(n_2168),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_4001),
.Y(n_4190)
);

AO31x2_ASAP7_75t_L g4191 ( 
.A1(n_3981),
.A2(n_566),
.A3(n_567),
.B(n_561),
.Y(n_4191)
);

OAI21x1_ASAP7_75t_L g4192 ( 
.A1(n_3831),
.A2(n_2185),
.B(n_2168),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_4014),
.B(n_1097),
.Y(n_4193)
);

OAI21x1_ASAP7_75t_L g4194 ( 
.A1(n_3980),
.A2(n_3873),
.B(n_3862),
.Y(n_4194)
);

AO21x2_ASAP7_75t_L g4195 ( 
.A1(n_3823),
.A2(n_2108),
.B(n_2104),
.Y(n_4195)
);

AOI21xp5_ASAP7_75t_L g4196 ( 
.A1(n_3846),
.A2(n_2110),
.B(n_2108),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_3833),
.B(n_1108),
.Y(n_4197)
);

OAI21xp5_ASAP7_75t_L g4198 ( 
.A1(n_3967),
.A2(n_1113),
.B(n_1109),
.Y(n_4198)
);

NAND2xp5_ASAP7_75t_L g4199 ( 
.A(n_4016),
.B(n_1115),
.Y(n_4199)
);

AND2x2_ASAP7_75t_L g4200 ( 
.A(n_3904),
.B(n_4002),
.Y(n_4200)
);

AOI21xp5_ASAP7_75t_L g4201 ( 
.A1(n_3888),
.A2(n_2110),
.B(n_2108),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_L g4202 ( 
.A(n_3918),
.B(n_1116),
.Y(n_4202)
);

INVx2_ASAP7_75t_L g4203 ( 
.A(n_4001),
.Y(n_4203)
);

NOR2xp33_ASAP7_75t_L g4204 ( 
.A(n_3853),
.B(n_3992),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_3854),
.B(n_1118),
.Y(n_4205)
);

NOR2xp33_ASAP7_75t_L g4206 ( 
.A(n_3947),
.B(n_1119),
.Y(n_4206)
);

BUFx6f_ASAP7_75t_L g4207 ( 
.A(n_3887),
.Y(n_4207)
);

NOR2xp33_ASAP7_75t_L g4208 ( 
.A(n_3979),
.B(n_1120),
.Y(n_4208)
);

O2A1O1Ixp5_ASAP7_75t_L g4209 ( 
.A1(n_3943),
.A2(n_3847),
.B(n_3930),
.C(n_3900),
.Y(n_4209)
);

OAI21xp5_ASAP7_75t_L g4210 ( 
.A1(n_3915),
.A2(n_1122),
.B(n_1121),
.Y(n_4210)
);

NAND2xp33_ASAP7_75t_L g4211 ( 
.A(n_3931),
.B(n_1138),
.Y(n_4211)
);

NOR2x1_ASAP7_75t_SL g4212 ( 
.A(n_3821),
.B(n_2108),
.Y(n_4212)
);

AO31x2_ASAP7_75t_L g4213 ( 
.A1(n_3989),
.A2(n_570),
.A3(n_572),
.B(n_568),
.Y(n_4213)
);

INVx4_ASAP7_75t_L g4214 ( 
.A(n_3887),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_3835),
.B(n_1125),
.Y(n_4215)
);

AND2x2_ASAP7_75t_L g4216 ( 
.A(n_3936),
.B(n_573),
.Y(n_4216)
);

OAI21x1_ASAP7_75t_L g4217 ( 
.A1(n_3838),
.A2(n_2185),
.B(n_2233),
.Y(n_4217)
);

INVx3_ASAP7_75t_L g4218 ( 
.A(n_3887),
.Y(n_4218)
);

NAND2x1p5_ASAP7_75t_L g4219 ( 
.A(n_3798),
.B(n_2110),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_3859),
.Y(n_4220)
);

A2O1A1Ixp33_ASAP7_75t_L g4221 ( 
.A1(n_3984),
.A2(n_1161),
.B(n_1131),
.C(n_1128),
.Y(n_4221)
);

BUFx3_ASAP7_75t_L g4222 ( 
.A(n_3986),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_3972),
.Y(n_4223)
);

NAND2xp5_ASAP7_75t_L g4224 ( 
.A(n_4018),
.B(n_1126),
.Y(n_4224)
);

NAND2x1p5_ASAP7_75t_L g4225 ( 
.A(n_3798),
.B(n_2110),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_L g4226 ( 
.A(n_4018),
.B(n_3960),
.Y(n_4226)
);

OAI21x1_ASAP7_75t_L g4227 ( 
.A1(n_3997),
.A2(n_2241),
.B(n_2233),
.Y(n_4227)
);

AOI21xp5_ASAP7_75t_L g4228 ( 
.A1(n_4017),
.A2(n_3997),
.B(n_3974),
.Y(n_4228)
);

OAI21x1_ASAP7_75t_L g4229 ( 
.A1(n_4013),
.A2(n_2241),
.B(n_2233),
.Y(n_4229)
);

OAI21xp5_ASAP7_75t_L g4230 ( 
.A1(n_3958),
.A2(n_1134),
.B(n_1132),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_3950),
.B(n_1140),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_3956),
.B(n_1147),
.Y(n_4232)
);

AOI21xp5_ASAP7_75t_L g4233 ( 
.A1(n_4017),
.A2(n_1926),
.B(n_1922),
.Y(n_4233)
);

AOI21xp5_ASAP7_75t_L g4234 ( 
.A1(n_4017),
.A2(n_1926),
.B(n_1922),
.Y(n_4234)
);

AO31x2_ASAP7_75t_L g4235 ( 
.A1(n_4011),
.A2(n_575),
.A3(n_576),
.B(n_574),
.Y(n_4235)
);

AOI21xp5_ASAP7_75t_SL g4236 ( 
.A1(n_3801),
.A2(n_1154),
.B(n_1148),
.Y(n_4236)
);

NOR2xp67_ASAP7_75t_L g4237 ( 
.A(n_3933),
.B(n_582),
.Y(n_4237)
);

BUFx3_ASAP7_75t_L g4238 ( 
.A(n_4015),
.Y(n_4238)
);

AOI21xp5_ASAP7_75t_L g4239 ( 
.A1(n_3974),
.A2(n_1926),
.B(n_1922),
.Y(n_4239)
);

AOI21xp5_ASAP7_75t_L g4240 ( 
.A1(n_3803),
.A2(n_1926),
.B(n_1922),
.Y(n_4240)
);

OAI21x1_ASAP7_75t_L g4241 ( 
.A1(n_3962),
.A2(n_3879),
.B(n_3803),
.Y(n_4241)
);

O2A1O1Ixp33_ASAP7_75t_L g4242 ( 
.A1(n_3858),
.A2(n_1163),
.B(n_1165),
.C(n_1160),
.Y(n_4242)
);

AO31x2_ASAP7_75t_L g4243 ( 
.A1(n_3948),
.A2(n_3940),
.A3(n_3999),
.B(n_3963),
.Y(n_4243)
);

AO32x2_ASAP7_75t_L g4244 ( 
.A1(n_3776),
.A2(n_1169),
.A3(n_1166),
.B1(n_4),
.B2(n_2),
.Y(n_4244)
);

AOI21xp5_ASAP7_75t_L g4245 ( 
.A1(n_3879),
.A2(n_1926),
.B(n_1922),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_3961),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_L g4247 ( 
.A(n_3965),
.B(n_2),
.Y(n_4247)
);

OAI21xp5_ASAP7_75t_L g4248 ( 
.A1(n_3916),
.A2(n_1767),
.B(n_1703),
.Y(n_4248)
);

NAND2xp5_ASAP7_75t_L g4249 ( 
.A(n_3970),
.B(n_3),
.Y(n_4249)
);

OAI21xp5_ASAP7_75t_L g4250 ( 
.A1(n_3973),
.A2(n_1767),
.B(n_1703),
.Y(n_4250)
);

OR2x2_ASAP7_75t_L g4251 ( 
.A(n_3975),
.B(n_4),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_3982),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_4000),
.B(n_4012),
.Y(n_4253)
);

BUFx3_ASAP7_75t_L g4254 ( 
.A(n_3998),
.Y(n_4254)
);

OAI22xp5_ASAP7_75t_L g4255 ( 
.A1(n_3850),
.A2(n_1959),
.B1(n_1970),
.B2(n_1948),
.Y(n_4255)
);

OAI21x1_ASAP7_75t_L g4256 ( 
.A1(n_3790),
.A2(n_2242),
.B(n_2241),
.Y(n_4256)
);

NAND2xp33_ASAP7_75t_SL g4257 ( 
.A(n_3782),
.B(n_5),
.Y(n_4257)
);

OAI21x1_ASAP7_75t_L g4258 ( 
.A1(n_3843),
.A2(n_2262),
.B(n_2242),
.Y(n_4258)
);

INVxp67_ASAP7_75t_L g4259 ( 
.A(n_3998),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_3998),
.Y(n_4260)
);

AOI21xp5_ASAP7_75t_L g4261 ( 
.A1(n_4008),
.A2(n_1943),
.B(n_1927),
.Y(n_4261)
);

OAI21xp33_ASAP7_75t_L g4262 ( 
.A1(n_3897),
.A2(n_5),
.B(n_6),
.Y(n_4262)
);

INVxp33_ASAP7_75t_SL g4263 ( 
.A(n_4077),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_SL g4264 ( 
.A(n_4146),
.B(n_4112),
.Y(n_4264)
);

INVx3_ASAP7_75t_L g4265 ( 
.A(n_4177),
.Y(n_4265)
);

OR2x2_ASAP7_75t_L g4266 ( 
.A(n_4038),
.B(n_3868),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_4098),
.B(n_3868),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_4155),
.B(n_3990),
.Y(n_4268)
);

O2A1O1Ixp33_ASAP7_75t_L g4269 ( 
.A1(n_4041),
.A2(n_3993),
.B(n_3990),
.C(n_8),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_4039),
.Y(n_4270)
);

CKINVDCx11_ASAP7_75t_R g4271 ( 
.A(n_4088),
.Y(n_4271)
);

BUFx3_ASAP7_75t_L g4272 ( 
.A(n_4043),
.Y(n_4272)
);

BUFx2_ASAP7_75t_L g4273 ( 
.A(n_4050),
.Y(n_4273)
);

OAI21xp5_ASAP7_75t_L g4274 ( 
.A1(n_4209),
.A2(n_3993),
.B(n_3776),
.Y(n_4274)
);

CKINVDCx16_ASAP7_75t_R g4275 ( 
.A(n_4032),
.Y(n_4275)
);

CKINVDCx11_ASAP7_75t_R g4276 ( 
.A(n_4032),
.Y(n_4276)
);

BUFx4_ASAP7_75t_SL g4277 ( 
.A(n_4037),
.Y(n_4277)
);

INVx1_ASAP7_75t_SL g4278 ( 
.A(n_4060),
.Y(n_4278)
);

AND2x4_ASAP7_75t_L g4279 ( 
.A(n_4177),
.B(n_586),
.Y(n_4279)
);

HB1xp67_ASAP7_75t_L g4280 ( 
.A(n_4058),
.Y(n_4280)
);

AND2x2_ASAP7_75t_L g4281 ( 
.A(n_4200),
.B(n_6),
.Y(n_4281)
);

INVxp67_ASAP7_75t_SL g4282 ( 
.A(n_4029),
.Y(n_4282)
);

INVxp67_ASAP7_75t_SL g4283 ( 
.A(n_4194),
.Y(n_4283)
);

INVx2_ASAP7_75t_L g4284 ( 
.A(n_4111),
.Y(n_4284)
);

AND2x4_ASAP7_75t_L g4285 ( 
.A(n_4072),
.B(n_591),
.Y(n_4285)
);

NAND2x1p5_ASAP7_75t_L g4286 ( 
.A(n_4102),
.B(n_1948),
.Y(n_4286)
);

AND2x2_ASAP7_75t_L g4287 ( 
.A(n_4040),
.B(n_7),
.Y(n_4287)
);

AOI21xp5_ASAP7_75t_L g4288 ( 
.A1(n_4147),
.A2(n_1943),
.B(n_1927),
.Y(n_4288)
);

O2A1O1Ixp33_ASAP7_75t_SL g4289 ( 
.A1(n_4262),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_4289)
);

INVx3_ASAP7_75t_SL g4290 ( 
.A(n_4068),
.Y(n_4290)
);

AND2x4_ASAP7_75t_L g4291 ( 
.A(n_4081),
.B(n_4096),
.Y(n_4291)
);

BUFx2_ASAP7_75t_L g4292 ( 
.A(n_4025),
.Y(n_4292)
);

INVx3_ASAP7_75t_L g4293 ( 
.A(n_4026),
.Y(n_4293)
);

BUFx2_ASAP7_75t_L g4294 ( 
.A(n_4025),
.Y(n_4294)
);

INVx2_ASAP7_75t_SL g4295 ( 
.A(n_4032),
.Y(n_4295)
);

AND2x2_ASAP7_75t_L g4296 ( 
.A(n_4070),
.B(n_9),
.Y(n_4296)
);

BUFx6f_ASAP7_75t_L g4297 ( 
.A(n_4080),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4117),
.Y(n_4298)
);

NOR2xp33_ASAP7_75t_L g4299 ( 
.A(n_4093),
.B(n_10),
.Y(n_4299)
);

NAND2xp5_ASAP7_75t_L g4300 ( 
.A(n_4042),
.B(n_13),
.Y(n_4300)
);

BUFx2_ASAP7_75t_L g4301 ( 
.A(n_4033),
.Y(n_4301)
);

AOI21xp5_ASAP7_75t_L g4302 ( 
.A1(n_4107),
.A2(n_1943),
.B(n_1927),
.Y(n_4302)
);

OAI22xp5_ASAP7_75t_L g4303 ( 
.A1(n_4226),
.A2(n_1883),
.B1(n_1890),
.B2(n_1878),
.Y(n_4303)
);

BUFx12f_ASAP7_75t_L g4304 ( 
.A(n_4066),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_L g4305 ( 
.A(n_4161),
.B(n_14),
.Y(n_4305)
);

OAI22x1_ASAP7_75t_L g4306 ( 
.A1(n_4067),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_4306)
);

OR2x6_ASAP7_75t_L g4307 ( 
.A(n_4261),
.B(n_1948),
.Y(n_4307)
);

AND2x4_ASAP7_75t_L g4308 ( 
.A(n_4033),
.B(n_592),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_4118),
.B(n_15),
.Y(n_4309)
);

BUFx12f_ASAP7_75t_L g4310 ( 
.A(n_4066),
.Y(n_4310)
);

INVx2_ASAP7_75t_SL g4311 ( 
.A(n_4222),
.Y(n_4311)
);

OAI21x1_ASAP7_75t_L g4312 ( 
.A1(n_4079),
.A2(n_4045),
.B(n_4148),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4130),
.Y(n_4313)
);

AOI22xp33_ASAP7_75t_L g4314 ( 
.A1(n_4101),
.A2(n_1883),
.B1(n_1890),
.B2(n_1878),
.Y(n_4314)
);

INVx2_ASAP7_75t_L g4315 ( 
.A(n_4063),
.Y(n_4315)
);

INVx5_ASAP7_75t_SL g4316 ( 
.A(n_4087),
.Y(n_4316)
);

NOR2xp33_ASAP7_75t_L g4317 ( 
.A(n_4152),
.B(n_16),
.Y(n_4317)
);

AOI22xp33_ASAP7_75t_L g4318 ( 
.A1(n_4257),
.A2(n_1883),
.B1(n_1890),
.B2(n_1878),
.Y(n_4318)
);

BUFx6f_ASAP7_75t_L g4319 ( 
.A(n_4080),
.Y(n_4319)
);

AND2x4_ASAP7_75t_L g4320 ( 
.A(n_4132),
.B(n_595),
.Y(n_4320)
);

CKINVDCx20_ASAP7_75t_R g4321 ( 
.A(n_4092),
.Y(n_4321)
);

AOI22xp33_ASAP7_75t_L g4322 ( 
.A1(n_4215),
.A2(n_1883),
.B1(n_1890),
.B2(n_1878),
.Y(n_4322)
);

AOI21xp5_ASAP7_75t_L g4323 ( 
.A1(n_4175),
.A2(n_1943),
.B(n_1927),
.Y(n_4323)
);

AOI21xp5_ASAP7_75t_L g4324 ( 
.A1(n_4059),
.A2(n_1943),
.B(n_1927),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_4024),
.B(n_17),
.Y(n_4325)
);

OAI22xp5_ASAP7_75t_L g4326 ( 
.A1(n_4141),
.A2(n_1906),
.B1(n_1959),
.B2(n_1948),
.Y(n_4326)
);

AOI22xp33_ASAP7_75t_SL g4327 ( 
.A1(n_4205),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_4327)
);

NOR2x1_ASAP7_75t_L g4328 ( 
.A(n_4054),
.B(n_1959),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4151),
.Y(n_4329)
);

BUFx2_ASAP7_75t_L g4330 ( 
.A(n_4132),
.Y(n_4330)
);

BUFx10_ASAP7_75t_L g4331 ( 
.A(n_4206),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4160),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_L g4333 ( 
.A(n_4246),
.B(n_4252),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_4085),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4086),
.Y(n_4335)
);

BUFx3_ASAP7_75t_L g4336 ( 
.A(n_4238),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4099),
.Y(n_4337)
);

OAI22xp5_ASAP7_75t_L g4338 ( 
.A1(n_4078),
.A2(n_4224),
.B1(n_4158),
.B2(n_4062),
.Y(n_4338)
);

AOI21xp5_ASAP7_75t_L g4339 ( 
.A1(n_4196),
.A2(n_1970),
.B(n_1959),
.Y(n_4339)
);

AND2x4_ASAP7_75t_L g4340 ( 
.A(n_4149),
.B(n_596),
.Y(n_4340)
);

AND2x4_ASAP7_75t_L g4341 ( 
.A(n_4149),
.B(n_4026),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_4036),
.B(n_18),
.Y(n_4342)
);

OAI22xp5_ASAP7_75t_L g4343 ( 
.A1(n_4159),
.A2(n_1906),
.B1(n_1970),
.B2(n_27),
.Y(n_4343)
);

BUFx2_ASAP7_75t_L g4344 ( 
.A(n_4028),
.Y(n_4344)
);

AND2x2_ASAP7_75t_L g4345 ( 
.A(n_4176),
.B(n_21),
.Y(n_4345)
);

NAND2xp5_ASAP7_75t_L g4346 ( 
.A(n_4164),
.B(n_21),
.Y(n_4346)
);

NAND2xp5_ASAP7_75t_L g4347 ( 
.A(n_4064),
.B(n_26),
.Y(n_4347)
);

INVxp67_ASAP7_75t_L g4348 ( 
.A(n_4253),
.Y(n_4348)
);

AOI22xp33_ASAP7_75t_L g4349 ( 
.A1(n_4084),
.A2(n_1906),
.B1(n_1767),
.B2(n_1703),
.Y(n_4349)
);

AND2x2_ASAP7_75t_L g4350 ( 
.A(n_4203),
.B(n_27),
.Y(n_4350)
);

AOI21xp5_ASAP7_75t_L g4351 ( 
.A1(n_4057),
.A2(n_1970),
.B(n_2242),
.Y(n_4351)
);

AND2x2_ASAP7_75t_L g4352 ( 
.A(n_4190),
.B(n_28),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_4129),
.B(n_29),
.Y(n_4353)
);

INVx2_ASAP7_75t_L g4354 ( 
.A(n_4139),
.Y(n_4354)
);

AOI21xp5_ASAP7_75t_L g4355 ( 
.A1(n_4116),
.A2(n_2268),
.B(n_2262),
.Y(n_4355)
);

INVxp67_ASAP7_75t_SL g4356 ( 
.A(n_4220),
.Y(n_4356)
);

INVx2_ASAP7_75t_L g4357 ( 
.A(n_4051),
.Y(n_4357)
);

OAI21x1_ASAP7_75t_L g4358 ( 
.A1(n_4115),
.A2(n_4135),
.B(n_4053),
.Y(n_4358)
);

AND2x4_ASAP7_75t_L g4359 ( 
.A(n_4028),
.B(n_597),
.Y(n_4359)
);

AND2x2_ASAP7_75t_L g4360 ( 
.A(n_4120),
.B(n_30),
.Y(n_4360)
);

BUFx3_ASAP7_75t_L g4361 ( 
.A(n_4254),
.Y(n_4361)
);

OR2x2_ASAP7_75t_L g4362 ( 
.A(n_4100),
.B(n_31),
.Y(n_4362)
);

BUFx4f_ASAP7_75t_SL g4363 ( 
.A(n_4080),
.Y(n_4363)
);

AOI22xp5_ASAP7_75t_L g4364 ( 
.A1(n_4055),
.A2(n_1906),
.B1(n_1767),
.B2(n_1703),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_L g4365 ( 
.A(n_4069),
.B(n_32),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4244),
.Y(n_4366)
);

INVx1_ASAP7_75t_SL g4367 ( 
.A(n_4204),
.Y(n_4367)
);

AND2x2_ASAP7_75t_L g4368 ( 
.A(n_4260),
.B(n_33),
.Y(n_4368)
);

AO21x2_ASAP7_75t_L g4369 ( 
.A1(n_4103),
.A2(n_33),
.B(n_34),
.Y(n_4369)
);

INVx8_ASAP7_75t_L g4370 ( 
.A(n_4102),
.Y(n_4370)
);

NOR2xp33_ASAP7_75t_L g4371 ( 
.A(n_4182),
.B(n_34),
.Y(n_4371)
);

NOR2x1_ASAP7_75t_SL g4372 ( 
.A(n_4102),
.B(n_1600),
.Y(n_4372)
);

OR2x2_ASAP7_75t_L g4373 ( 
.A(n_4056),
.B(n_35),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_SL g4374 ( 
.A(n_4237),
.B(n_1600),
.Y(n_4374)
);

A2O1A1Ixp33_ASAP7_75t_SL g4375 ( 
.A1(n_4187),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_4375)
);

INVx5_ASAP7_75t_L g4376 ( 
.A(n_4128),
.Y(n_4376)
);

CKINVDCx6p67_ASAP7_75t_R g4377 ( 
.A(n_4082),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4244),
.Y(n_4378)
);

AND2x2_ASAP7_75t_L g4379 ( 
.A(n_4074),
.B(n_36),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_L g4380 ( 
.A(n_4095),
.B(n_37),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_4244),
.Y(n_4381)
);

INVx1_ASAP7_75t_SL g4382 ( 
.A(n_4082),
.Y(n_4382)
);

AOI21xp5_ASAP7_75t_L g4383 ( 
.A1(n_4030),
.A2(n_2268),
.B(n_2262),
.Y(n_4383)
);

AOI21xp33_ASAP7_75t_L g4384 ( 
.A1(n_4124),
.A2(n_38),
.B(n_40),
.Y(n_4384)
);

CKINVDCx6p67_ASAP7_75t_R g4385 ( 
.A(n_4082),
.Y(n_4385)
);

AOI21xp5_ASAP7_75t_L g4386 ( 
.A1(n_4076),
.A2(n_2285),
.B(n_2268),
.Y(n_4386)
);

BUFx2_ASAP7_75t_SL g4387 ( 
.A(n_4214),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_L g4388 ( 
.A(n_4197),
.B(n_38),
.Y(n_4388)
);

BUFx12f_ASAP7_75t_L g4389 ( 
.A(n_4074),
.Y(n_4389)
);

INVx5_ASAP7_75t_L g4390 ( 
.A(n_4128),
.Y(n_4390)
);

INVx2_ASAP7_75t_L g4391 ( 
.A(n_4218),
.Y(n_4391)
);

NAND2x1p5_ASAP7_75t_L g4392 ( 
.A(n_4241),
.B(n_4214),
.Y(n_4392)
);

A2O1A1Ixp33_ASAP7_75t_L g4393 ( 
.A1(n_4242),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_4393)
);

NOR2xp33_ASAP7_75t_L g4394 ( 
.A(n_4104),
.B(n_41),
.Y(n_4394)
);

BUFx6f_ASAP7_75t_L g4395 ( 
.A(n_4140),
.Y(n_4395)
);

INVx3_ASAP7_75t_L g4396 ( 
.A(n_4140),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4170),
.Y(n_4397)
);

INVx3_ASAP7_75t_L g4398 ( 
.A(n_4140),
.Y(n_4398)
);

AOI22xp5_ASAP7_75t_L g4399 ( 
.A1(n_4208),
.A2(n_1767),
.B1(n_1703),
.B2(n_1638),
.Y(n_4399)
);

AOI22xp33_ASAP7_75t_L g4400 ( 
.A1(n_4165),
.A2(n_1638),
.B1(n_1701),
.B2(n_1656),
.Y(n_4400)
);

AOI21xp5_ASAP7_75t_L g4401 ( 
.A1(n_4089),
.A2(n_2288),
.B(n_2285),
.Y(n_4401)
);

A2O1A1Ixp33_ASAP7_75t_L g4402 ( 
.A1(n_4210),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_4402)
);

CKINVDCx6p67_ASAP7_75t_R g4403 ( 
.A(n_4207),
.Y(n_4403)
);

AND2x2_ASAP7_75t_L g4404 ( 
.A(n_4259),
.B(n_43),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_L g4405 ( 
.A(n_4172),
.B(n_44),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_4170),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_SL g4407 ( 
.A(n_4027),
.B(n_1627),
.Y(n_4407)
);

BUFx3_ASAP7_75t_L g4408 ( 
.A(n_4207),
.Y(n_4408)
);

A2O1A1Ixp33_ASAP7_75t_L g4409 ( 
.A1(n_4154),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_4409)
);

NAND2xp5_ASAP7_75t_L g4410 ( 
.A(n_4123),
.B(n_47),
.Y(n_4410)
);

BUFx6f_ASAP7_75t_SL g4411 ( 
.A(n_4207),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_L g4412 ( 
.A(n_4138),
.B(n_48),
.Y(n_4412)
);

NOR2xp33_ASAP7_75t_L g4413 ( 
.A(n_4065),
.B(n_50),
.Y(n_4413)
);

INVx8_ASAP7_75t_L g4414 ( 
.A(n_4218),
.Y(n_4414)
);

INVx2_ASAP7_75t_L g4415 ( 
.A(n_4170),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4163),
.Y(n_4416)
);

OAI22xp5_ASAP7_75t_L g4417 ( 
.A1(n_4052),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_4417)
);

AO21x1_ASAP7_75t_L g4418 ( 
.A1(n_4143),
.A2(n_53),
.B(n_54),
.Y(n_4418)
);

OR2x6_ASAP7_75t_SL g4419 ( 
.A(n_4251),
.B(n_4247),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4113),
.Y(n_4420)
);

AOI21xp5_ASAP7_75t_L g4421 ( 
.A1(n_4183),
.A2(n_2288),
.B(n_2285),
.Y(n_4421)
);

O2A1O1Ixp5_ASAP7_75t_SL g4422 ( 
.A1(n_4108),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_4422)
);

AND2x2_ASAP7_75t_L g4423 ( 
.A(n_4216),
.B(n_4243),
.Y(n_4423)
);

NAND2xp5_ASAP7_75t_L g4424 ( 
.A(n_4153),
.B(n_55),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4106),
.Y(n_4425)
);

AOI22xp33_ASAP7_75t_L g4426 ( 
.A1(n_4223),
.A2(n_1701),
.B1(n_1656),
.B2(n_1664),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_4122),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_4122),
.Y(n_4428)
);

NAND2x1_ASAP7_75t_L g4429 ( 
.A(n_4156),
.B(n_4075),
.Y(n_4429)
);

INVx3_ASAP7_75t_L g4430 ( 
.A(n_4023),
.Y(n_4430)
);

AOI22xp33_ASAP7_75t_L g4431 ( 
.A1(n_4185),
.A2(n_1701),
.B1(n_1656),
.B2(n_1664),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_L g4432 ( 
.A(n_4166),
.B(n_56),
.Y(n_4432)
);

INVx3_ASAP7_75t_L g4433 ( 
.A(n_4219),
.Y(n_4433)
);

OAI22xp5_ASAP7_75t_L g4434 ( 
.A1(n_4171),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_4434)
);

BUFx3_ASAP7_75t_L g4435 ( 
.A(n_4225),
.Y(n_4435)
);

INVx3_ASAP7_75t_L g4436 ( 
.A(n_4243),
.Y(n_4436)
);

AO31x2_ASAP7_75t_L g4437 ( 
.A1(n_4049),
.A2(n_61),
.A3(n_59),
.B(n_60),
.Y(n_4437)
);

AOI22xp33_ASAP7_75t_L g4438 ( 
.A1(n_4249),
.A2(n_1701),
.B1(n_1656),
.B2(n_1664),
.Y(n_4438)
);

CKINVDCx5p33_ASAP7_75t_R g4439 ( 
.A(n_4202),
.Y(n_4439)
);

CKINVDCx5p33_ASAP7_75t_R g4440 ( 
.A(n_4097),
.Y(n_4440)
);

INVx1_ASAP7_75t_SL g4441 ( 
.A(n_4109),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_L g4442 ( 
.A(n_4173),
.B(n_60),
.Y(n_4442)
);

AOI22xp33_ASAP7_75t_L g4443 ( 
.A1(n_4105),
.A2(n_1701),
.B1(n_1664),
.B2(n_1627),
.Y(n_4443)
);

AND2x4_ASAP7_75t_L g4444 ( 
.A(n_4243),
.B(n_601),
.Y(n_4444)
);

AND2x2_ASAP7_75t_L g4445 ( 
.A(n_4235),
.B(n_61),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_4163),
.Y(n_4446)
);

INVx2_ASAP7_75t_L g4447 ( 
.A(n_4163),
.Y(n_4447)
);

INVx3_ASAP7_75t_L g4448 ( 
.A(n_4179),
.Y(n_4448)
);

INVx1_ASAP7_75t_SL g4449 ( 
.A(n_4181),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_L g4450 ( 
.A(n_4174),
.B(n_62),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4168),
.Y(n_4451)
);

AOI21xp5_ASAP7_75t_L g4452 ( 
.A1(n_4183),
.A2(n_2296),
.B(n_2288),
.Y(n_4452)
);

NAND2x1p5_ASAP7_75t_L g4453 ( 
.A(n_4031),
.B(n_1627),
.Y(n_4453)
);

BUFx12f_ASAP7_75t_L g4454 ( 
.A(n_4179),
.Y(n_4454)
);

BUFx4f_ASAP7_75t_SL g4455 ( 
.A(n_4090),
.Y(n_4455)
);

INVxp67_ASAP7_75t_L g4456 ( 
.A(n_4199),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4122),
.Y(n_4457)
);

CKINVDCx11_ASAP7_75t_R g4458 ( 
.A(n_4114),
.Y(n_4458)
);

AOI21xp5_ASAP7_75t_L g4459 ( 
.A1(n_4186),
.A2(n_4184),
.B(n_4034),
.Y(n_4459)
);

AND2x2_ASAP7_75t_L g4460 ( 
.A(n_4235),
.B(n_62),
.Y(n_4460)
);

AOI22xp33_ASAP7_75t_L g4461 ( 
.A1(n_4188),
.A2(n_1627),
.B1(n_1762),
.B2(n_66),
.Y(n_4461)
);

OAI21x1_ASAP7_75t_L g4462 ( 
.A1(n_4035),
.A2(n_2296),
.B(n_607),
.Y(n_4462)
);

CKINVDCx5p33_ASAP7_75t_R g4463 ( 
.A(n_4193),
.Y(n_4463)
);

INVx2_ASAP7_75t_L g4464 ( 
.A(n_4168),
.Y(n_4464)
);

CKINVDCx20_ASAP7_75t_R g4465 ( 
.A(n_4142),
.Y(n_4465)
);

INVx2_ASAP7_75t_L g4466 ( 
.A(n_4168),
.Y(n_4466)
);

BUFx10_ASAP7_75t_L g4467 ( 
.A(n_4211),
.Y(n_4467)
);

OAI22xp5_ASAP7_75t_SL g4468 ( 
.A1(n_4131),
.A2(n_67),
.B1(n_63),
.B2(n_64),
.Y(n_4468)
);

INVx1_ASAP7_75t_L g4469 ( 
.A(n_4125),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_SL g4470 ( 
.A(n_4180),
.B(n_1762),
.Y(n_4470)
);

OR2x6_ASAP7_75t_L g4471 ( 
.A(n_4239),
.B(n_604),
.Y(n_4471)
);

AOI22xp5_ASAP7_75t_L g4472 ( 
.A1(n_4061),
.A2(n_68),
.B1(n_64),
.B2(n_67),
.Y(n_4472)
);

NAND2xp5_ASAP7_75t_L g4473 ( 
.A(n_4231),
.B(n_68),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_L g4474 ( 
.A(n_4232),
.B(n_70),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4125),
.Y(n_4475)
);

INVxp67_ASAP7_75t_SL g4476 ( 
.A(n_4201),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_4125),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4094),
.Y(n_4478)
);

OAI22xp5_ASAP7_75t_L g4479 ( 
.A1(n_4236),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_4479)
);

AOI21xp5_ASAP7_75t_L g4480 ( 
.A1(n_4046),
.A2(n_2296),
.B(n_2214),
.Y(n_4480)
);

OAI22xp5_ASAP7_75t_L g4481 ( 
.A1(n_4230),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_4235),
.Y(n_4482)
);

INVx2_ASAP7_75t_L g4483 ( 
.A(n_4195),
.Y(n_4483)
);

BUFx6f_ASAP7_75t_L g4484 ( 
.A(n_4256),
.Y(n_4484)
);

NAND2xp5_ASAP7_75t_L g4485 ( 
.A(n_4145),
.B(n_75),
.Y(n_4485)
);

AOI21xp5_ASAP7_75t_L g4486 ( 
.A1(n_4071),
.A2(n_4250),
.B(n_4073),
.Y(n_4486)
);

AND2x2_ASAP7_75t_L g4487 ( 
.A(n_4213),
.B(n_75),
.Y(n_4487)
);

NAND2xp5_ASAP7_75t_L g4488 ( 
.A(n_4167),
.B(n_76),
.Y(n_4488)
);

AOI21xp5_ASAP7_75t_L g4489 ( 
.A1(n_4228),
.A2(n_2214),
.B(n_2210),
.Y(n_4489)
);

OAI21x1_ASAP7_75t_L g4490 ( 
.A1(n_4048),
.A2(n_609),
.B(n_608),
.Y(n_4490)
);

AND2x2_ASAP7_75t_L g4491 ( 
.A(n_4213),
.B(n_77),
.Y(n_4491)
);

AO21x1_ASAP7_75t_L g4492 ( 
.A1(n_4121),
.A2(n_78),
.B(n_79),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_L g4493 ( 
.A(n_4083),
.B(n_78),
.Y(n_4493)
);

AO21x2_ASAP7_75t_L g4494 ( 
.A1(n_4047),
.A2(n_83),
.B(n_85),
.Y(n_4494)
);

OAI22xp5_ASAP7_75t_L g4495 ( 
.A1(n_4221),
.A2(n_87),
.B1(n_83),
.B2(n_86),
.Y(n_4495)
);

INVx3_ASAP7_75t_L g4496 ( 
.A(n_4213),
.Y(n_4496)
);

INVx5_ASAP7_75t_L g4497 ( 
.A(n_4212),
.Y(n_4497)
);

INVx2_ASAP7_75t_SL g4498 ( 
.A(n_4191),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4191),
.Y(n_4499)
);

AOI22xp5_ASAP7_75t_L g4500 ( 
.A1(n_4119),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_4500)
);

NAND2xp5_ASAP7_75t_L g4501 ( 
.A(n_4162),
.B(n_89),
.Y(n_4501)
);

INVx2_ASAP7_75t_SL g4502 ( 
.A(n_4191),
.Y(n_4502)
);

AND2x2_ASAP7_75t_L g4503 ( 
.A(n_4217),
.B(n_89),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_L g4504 ( 
.A(n_4282),
.B(n_4162),
.Y(n_4504)
);

INVx5_ASAP7_75t_L g4505 ( 
.A(n_4370),
.Y(n_4505)
);

AOI22xp33_ASAP7_75t_L g4506 ( 
.A1(n_4264),
.A2(n_4198),
.B1(n_4248),
.B2(n_4255),
.Y(n_4506)
);

AOI22xp33_ASAP7_75t_L g4507 ( 
.A1(n_4468),
.A2(n_4091),
.B1(n_4227),
.B2(n_4229),
.Y(n_4507)
);

OAI22xp33_ASAP7_75t_L g4508 ( 
.A1(n_4472),
.A2(n_4240),
.B1(n_4245),
.B2(n_4136),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_4280),
.B(n_4162),
.Y(n_4509)
);

OAI22xp5_ASAP7_75t_L g4510 ( 
.A1(n_4402),
.A2(n_4234),
.B1(n_4233),
.B2(n_4212),
.Y(n_4510)
);

AOI22xp5_ASAP7_75t_L g4511 ( 
.A1(n_4481),
.A2(n_4044),
.B1(n_4258),
.B2(n_4127),
.Y(n_4511)
);

BUFx12f_ASAP7_75t_L g4512 ( 
.A(n_4276),
.Y(n_4512)
);

AOI22xp33_ASAP7_75t_L g4513 ( 
.A1(n_4458),
.A2(n_4134),
.B1(n_4133),
.B2(n_4137),
.Y(n_4513)
);

OAI22xp33_ASAP7_75t_L g4514 ( 
.A1(n_4500),
.A2(n_4110),
.B1(n_92),
.B2(n_90),
.Y(n_4514)
);

INVx1_ASAP7_75t_SL g4515 ( 
.A(n_4367),
.Y(n_4515)
);

INVx4_ASAP7_75t_L g4516 ( 
.A(n_4370),
.Y(n_4516)
);

INVx4_ASAP7_75t_L g4517 ( 
.A(n_4414),
.Y(n_4517)
);

BUFx3_ASAP7_75t_L g4518 ( 
.A(n_4336),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_4270),
.Y(n_4519)
);

AOI22xp33_ASAP7_75t_L g4520 ( 
.A1(n_4317),
.A2(n_4144),
.B1(n_4189),
.B2(n_4178),
.Y(n_4520)
);

BUFx2_ASAP7_75t_SL g4521 ( 
.A(n_4411),
.Y(n_4521)
);

INVx1_ASAP7_75t_L g4522 ( 
.A(n_4298),
.Y(n_4522)
);

AOI22xp33_ASAP7_75t_SL g4523 ( 
.A1(n_4445),
.A2(n_4460),
.B1(n_4338),
.B2(n_4485),
.Y(n_4523)
);

AOI22xp33_ASAP7_75t_L g4524 ( 
.A1(n_4384),
.A2(n_4157),
.B1(n_4150),
.B2(n_4126),
.Y(n_4524)
);

AOI22xp5_ASAP7_75t_L g4525 ( 
.A1(n_4479),
.A2(n_4418),
.B1(n_4495),
.B2(n_4492),
.Y(n_4525)
);

INVx3_ASAP7_75t_L g4526 ( 
.A(n_4291),
.Y(n_4526)
);

AOI22xp33_ASAP7_75t_SL g4527 ( 
.A1(n_4488),
.A2(n_4192),
.B1(n_4169),
.B2(n_93),
.Y(n_4527)
);

BUFx10_ASAP7_75t_L g4528 ( 
.A(n_4463),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4298),
.Y(n_4529)
);

CKINVDCx6p67_ASAP7_75t_R g4530 ( 
.A(n_4290),
.Y(n_4530)
);

INVx6_ASAP7_75t_L g4531 ( 
.A(n_4275),
.Y(n_4531)
);

OR2x2_ASAP7_75t_L g4532 ( 
.A(n_4278),
.B(n_91),
.Y(n_4532)
);

AOI22xp33_ASAP7_75t_L g4533 ( 
.A1(n_4371),
.A2(n_95),
.B1(n_92),
.B2(n_94),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4313),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4313),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4291),
.Y(n_4536)
);

INVx2_ASAP7_75t_SL g4537 ( 
.A(n_4272),
.Y(n_4537)
);

CKINVDCx11_ASAP7_75t_R g4538 ( 
.A(n_4271),
.Y(n_4538)
);

INVx6_ASAP7_75t_L g4539 ( 
.A(n_4467),
.Y(n_4539)
);

CKINVDCx11_ASAP7_75t_R g4540 ( 
.A(n_4321),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_4284),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4329),
.Y(n_4542)
);

BUFx12f_ASAP7_75t_L g4543 ( 
.A(n_4467),
.Y(n_4543)
);

CKINVDCx20_ASAP7_75t_R g4544 ( 
.A(n_4455),
.Y(n_4544)
);

BUFx12f_ASAP7_75t_L g4545 ( 
.A(n_4331),
.Y(n_4545)
);

AOI22xp33_ASAP7_75t_L g4546 ( 
.A1(n_4299),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_4546)
);

INVxp67_ASAP7_75t_SL g4547 ( 
.A(n_4356),
.Y(n_4547)
);

AOI22xp33_ASAP7_75t_L g4548 ( 
.A1(n_4394),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_4548)
);

CKINVDCx6p67_ASAP7_75t_R g4549 ( 
.A(n_4304),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_4273),
.B(n_101),
.Y(n_4550)
);

INVx2_ASAP7_75t_SL g4551 ( 
.A(n_4311),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_L g4552 ( 
.A(n_4348),
.B(n_101),
.Y(n_4552)
);

AOI22xp33_ASAP7_75t_L g4553 ( 
.A1(n_4423),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_4332),
.Y(n_4554)
);

OAI22xp5_ASAP7_75t_L g4555 ( 
.A1(n_4393),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_4555)
);

AND2x4_ASAP7_75t_L g4556 ( 
.A(n_4292),
.B(n_105),
.Y(n_4556)
);

INVx4_ASAP7_75t_L g4557 ( 
.A(n_4414),
.Y(n_4557)
);

NAND2x1p5_ASAP7_75t_L g4558 ( 
.A(n_4376),
.B(n_1674),
.Y(n_4558)
);

AOI22xp33_ASAP7_75t_L g4559 ( 
.A1(n_4327),
.A2(n_4417),
.B1(n_4444),
.B2(n_4434),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_4334),
.Y(n_4560)
);

INVx2_ASAP7_75t_L g4561 ( 
.A(n_4335),
.Y(n_4561)
);

NAND2xp5_ASAP7_75t_L g4562 ( 
.A(n_4357),
.B(n_107),
.Y(n_4562)
);

INVx3_ASAP7_75t_L g4563 ( 
.A(n_4265),
.Y(n_4563)
);

AOI22xp33_ASAP7_75t_L g4564 ( 
.A1(n_4444),
.A2(n_110),
.B1(n_107),
.B2(n_109),
.Y(n_4564)
);

INVx6_ASAP7_75t_L g4565 ( 
.A(n_4310),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_L g4566 ( 
.A(n_4333),
.B(n_109),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_4337),
.Y(n_4567)
);

CKINVDCx11_ASAP7_75t_R g4568 ( 
.A(n_4331),
.Y(n_4568)
);

INVx6_ASAP7_75t_L g4569 ( 
.A(n_4297),
.Y(n_4569)
);

BUFx3_ASAP7_75t_L g4570 ( 
.A(n_4263),
.Y(n_4570)
);

CKINVDCx5p33_ASAP7_75t_R g4571 ( 
.A(n_4277),
.Y(n_4571)
);

INVx2_ASAP7_75t_L g4572 ( 
.A(n_4315),
.Y(n_4572)
);

OAI21xp5_ASAP7_75t_L g4573 ( 
.A1(n_4269),
.A2(n_110),
.B(n_111),
.Y(n_4573)
);

OAI22xp33_ASAP7_75t_L g4574 ( 
.A1(n_4471),
.A2(n_116),
.B1(n_112),
.B2(n_115),
.Y(n_4574)
);

INVx2_ASAP7_75t_L g4575 ( 
.A(n_4354),
.Y(n_4575)
);

AOI22xp33_ASAP7_75t_L g4576 ( 
.A1(n_4470),
.A2(n_117),
.B1(n_112),
.B2(n_116),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_4482),
.Y(n_4577)
);

INVx2_ASAP7_75t_SL g4578 ( 
.A(n_4361),
.Y(n_4578)
);

HB1xp67_ASAP7_75t_L g4579 ( 
.A(n_4294),
.Y(n_4579)
);

CKINVDCx11_ASAP7_75t_R g4580 ( 
.A(n_4419),
.Y(n_4580)
);

AOI22xp33_ASAP7_75t_L g4581 ( 
.A1(n_4407),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_4581)
);

CKINVDCx5p33_ASAP7_75t_R g4582 ( 
.A(n_4440),
.Y(n_4582)
);

OAI22xp5_ASAP7_75t_L g4583 ( 
.A1(n_4461),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_4583)
);

INVx4_ASAP7_75t_SL g4584 ( 
.A(n_4411),
.Y(n_4584)
);

BUFx3_ASAP7_75t_L g4585 ( 
.A(n_4295),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_4406),
.Y(n_4586)
);

AOI22xp5_ASAP7_75t_L g4587 ( 
.A1(n_4449),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4406),
.Y(n_4588)
);

BUFx2_ASAP7_75t_SL g4589 ( 
.A(n_4465),
.Y(n_4589)
);

BUFx2_ASAP7_75t_L g4590 ( 
.A(n_4344),
.Y(n_4590)
);

INVxp67_ASAP7_75t_SL g4591 ( 
.A(n_4436),
.Y(n_4591)
);

NAND2xp5_ASAP7_75t_L g4592 ( 
.A(n_4268),
.B(n_123),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_4366),
.Y(n_4593)
);

BUFx6f_ASAP7_75t_L g4594 ( 
.A(n_4297),
.Y(n_4594)
);

OAI22xp5_ASAP7_75t_L g4595 ( 
.A1(n_4493),
.A2(n_4316),
.B1(n_4409),
.B2(n_4441),
.Y(n_4595)
);

AOI22xp5_ASAP7_75t_L g4596 ( 
.A1(n_4454),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4378),
.Y(n_4597)
);

OAI22xp5_ASAP7_75t_L g4598 ( 
.A1(n_4316),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_4598)
);

AOI22xp5_ASAP7_75t_L g4599 ( 
.A1(n_4343),
.A2(n_4413),
.B1(n_4439),
.B2(n_4448),
.Y(n_4599)
);

BUFx6f_ASAP7_75t_L g4600 ( 
.A(n_4297),
.Y(n_4600)
);

BUFx12f_ASAP7_75t_L g4601 ( 
.A(n_4362),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_4266),
.Y(n_4602)
);

BUFx8_ASAP7_75t_L g4603 ( 
.A(n_4281),
.Y(n_4603)
);

INVx5_ASAP7_75t_L g4604 ( 
.A(n_4471),
.Y(n_4604)
);

INVx6_ASAP7_75t_L g4605 ( 
.A(n_4319),
.Y(n_4605)
);

CKINVDCx20_ASAP7_75t_R g4606 ( 
.A(n_4363),
.Y(n_4606)
);

CKINVDCx5p33_ASAP7_75t_R g4607 ( 
.A(n_4408),
.Y(n_4607)
);

OAI22xp33_ASAP7_75t_SL g4608 ( 
.A1(n_4381),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_4608)
);

AOI22xp33_ASAP7_75t_L g4609 ( 
.A1(n_4487),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4397),
.Y(n_4610)
);

INVx2_ASAP7_75t_L g4611 ( 
.A(n_4301),
.Y(n_4611)
);

INVx3_ASAP7_75t_L g4612 ( 
.A(n_4265),
.Y(n_4612)
);

NOR2xp33_ASAP7_75t_L g4613 ( 
.A(n_4456),
.B(n_132),
.Y(n_4613)
);

INVx2_ASAP7_75t_L g4614 ( 
.A(n_4330),
.Y(n_4614)
);

INVx3_ASAP7_75t_L g4615 ( 
.A(n_4293),
.Y(n_4615)
);

INVx2_ASAP7_75t_L g4616 ( 
.A(n_4391),
.Y(n_4616)
);

INVx6_ASAP7_75t_L g4617 ( 
.A(n_4319),
.Y(n_4617)
);

BUFx12f_ASAP7_75t_L g4618 ( 
.A(n_4287),
.Y(n_4618)
);

INVx2_ASAP7_75t_L g4619 ( 
.A(n_4436),
.Y(n_4619)
);

AOI22xp33_ASAP7_75t_L g4620 ( 
.A1(n_4491),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_4620)
);

OAI22xp33_ASAP7_75t_L g4621 ( 
.A1(n_4373),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4283),
.Y(n_4622)
);

AOI22xp33_ASAP7_75t_SL g4623 ( 
.A1(n_4448),
.A2(n_139),
.B1(n_135),
.B2(n_138),
.Y(n_4623)
);

INVx1_ASAP7_75t_L g4624 ( 
.A(n_4427),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4428),
.Y(n_4625)
);

CKINVDCx11_ASAP7_75t_R g4626 ( 
.A(n_4389),
.Y(n_4626)
);

CKINVDCx11_ASAP7_75t_R g4627 ( 
.A(n_4377),
.Y(n_4627)
);

AND2x2_ASAP7_75t_L g4628 ( 
.A(n_4293),
.B(n_4341),
.Y(n_4628)
);

INVx6_ASAP7_75t_L g4629 ( 
.A(n_4319),
.Y(n_4629)
);

BUFx10_ASAP7_75t_L g4630 ( 
.A(n_4279),
.Y(n_4630)
);

INVx3_ASAP7_75t_L g4631 ( 
.A(n_4392),
.Y(n_4631)
);

INVx5_ASAP7_75t_L g4632 ( 
.A(n_4307),
.Y(n_4632)
);

INVx2_ASAP7_75t_L g4633 ( 
.A(n_4415),
.Y(n_4633)
);

INVx6_ASAP7_75t_L g4634 ( 
.A(n_4395),
.Y(n_4634)
);

OAI22xp5_ASAP7_75t_L g4635 ( 
.A1(n_4431),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_4635)
);

AOI22xp33_ASAP7_75t_L g4636 ( 
.A1(n_4306),
.A2(n_143),
.B1(n_140),
.B2(n_142),
.Y(n_4636)
);

BUFx8_ASAP7_75t_L g4637 ( 
.A(n_4360),
.Y(n_4637)
);

BUFx12f_ASAP7_75t_L g4638 ( 
.A(n_4309),
.Y(n_4638)
);

INVx2_ASAP7_75t_L g4639 ( 
.A(n_4267),
.Y(n_4639)
);

INVx2_ASAP7_75t_L g4640 ( 
.A(n_4483),
.Y(n_4640)
);

OAI21xp5_ASAP7_75t_L g4641 ( 
.A1(n_4429),
.A2(n_4324),
.B(n_4459),
.Y(n_4641)
);

AOI22xp33_ASAP7_75t_L g4642 ( 
.A1(n_4285),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4457),
.Y(n_4643)
);

AOI22xp5_ASAP7_75t_L g4644 ( 
.A1(n_4374),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_4644)
);

NAND2x1p5_ASAP7_75t_L g4645 ( 
.A(n_4376),
.B(n_1674),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4416),
.Y(n_4646)
);

BUFx2_ASAP7_75t_L g4647 ( 
.A(n_4341),
.Y(n_4647)
);

INVx2_ASAP7_75t_L g4648 ( 
.A(n_4396),
.Y(n_4648)
);

AOI22xp33_ASAP7_75t_SL g4649 ( 
.A1(n_4501),
.A2(n_149),
.B1(n_145),
.B2(n_148),
.Y(n_4649)
);

INVx2_ASAP7_75t_L g4650 ( 
.A(n_4396),
.Y(n_4650)
);

AOI22xp33_ASAP7_75t_SL g4651 ( 
.A1(n_4285),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_4416),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4446),
.Y(n_4653)
);

BUFx2_ASAP7_75t_L g4654 ( 
.A(n_4398),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_4398),
.Y(n_4655)
);

BUFx6f_ASAP7_75t_L g4656 ( 
.A(n_4395),
.Y(n_4656)
);

CKINVDCx11_ASAP7_75t_R g4657 ( 
.A(n_4385),
.Y(n_4657)
);

INVx2_ASAP7_75t_L g4658 ( 
.A(n_4446),
.Y(n_4658)
);

AOI22xp33_ASAP7_75t_L g4659 ( 
.A1(n_4326),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_4659)
);

INVx1_ASAP7_75t_L g4660 ( 
.A(n_4451),
.Y(n_4660)
);

BUFx2_ASAP7_75t_SL g4661 ( 
.A(n_4395),
.Y(n_4661)
);

OAI22xp5_ASAP7_75t_L g4662 ( 
.A1(n_4349),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_4662)
);

BUFx6f_ASAP7_75t_L g4663 ( 
.A(n_4403),
.Y(n_4663)
);

BUFx12f_ASAP7_75t_L g4664 ( 
.A(n_4359),
.Y(n_4664)
);

OAI22xp33_ASAP7_75t_L g4665 ( 
.A1(n_4274),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_4665)
);

AOI22xp33_ASAP7_75t_L g4666 ( 
.A1(n_4314),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_4666)
);

AOI22xp33_ASAP7_75t_SL g4667 ( 
.A1(n_4369),
.A2(n_163),
.B1(n_157),
.B2(n_159),
.Y(n_4667)
);

BUFx12f_ASAP7_75t_SL g4668 ( 
.A(n_4379),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4451),
.Y(n_4669)
);

CKINVDCx11_ASAP7_75t_R g4670 ( 
.A(n_4382),
.Y(n_4670)
);

CKINVDCx11_ASAP7_75t_R g4671 ( 
.A(n_4359),
.Y(n_4671)
);

OAI21xp5_ASAP7_75t_SL g4672 ( 
.A1(n_4405),
.A2(n_163),
.B(n_164),
.Y(n_4672)
);

BUFx6f_ASAP7_75t_L g4673 ( 
.A(n_4435),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_4499),
.Y(n_4674)
);

BUFx4_ASAP7_75t_SL g4675 ( 
.A(n_4307),
.Y(n_4675)
);

BUFx12f_ASAP7_75t_L g4676 ( 
.A(n_4296),
.Y(n_4676)
);

AOI22xp33_ASAP7_75t_SL g4677 ( 
.A1(n_4494),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4437),
.Y(n_4678)
);

AOI22xp33_ASAP7_75t_L g4679 ( 
.A1(n_4503),
.A2(n_168),
.B1(n_165),
.B2(n_167),
.Y(n_4679)
);

CKINVDCx10_ASAP7_75t_R g4680 ( 
.A(n_4387),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_4437),
.Y(n_4681)
);

BUFx2_ASAP7_75t_L g4682 ( 
.A(n_4430),
.Y(n_4682)
);

AOI22xp33_ASAP7_75t_SL g4683 ( 
.A1(n_4388),
.A2(n_4412),
.B1(n_4424),
.B2(n_4410),
.Y(n_4683)
);

INVx2_ASAP7_75t_L g4684 ( 
.A(n_4447),
.Y(n_4684)
);

BUFx3_ASAP7_75t_L g4685 ( 
.A(n_4430),
.Y(n_4685)
);

BUFx6f_ASAP7_75t_L g4686 ( 
.A(n_4279),
.Y(n_4686)
);

INVx2_ASAP7_75t_SL g4687 ( 
.A(n_4376),
.Y(n_4687)
);

CKINVDCx20_ASAP7_75t_R g4688 ( 
.A(n_4342),
.Y(n_4688)
);

OAI22xp5_ASAP7_75t_L g4689 ( 
.A1(n_4318),
.A2(n_170),
.B1(n_167),
.B2(n_169),
.Y(n_4689)
);

INVx2_ASAP7_75t_L g4690 ( 
.A(n_4464),
.Y(n_4690)
);

INVx1_ASAP7_75t_L g4691 ( 
.A(n_4437),
.Y(n_4691)
);

AOI22xp33_ASAP7_75t_L g4692 ( 
.A1(n_4473),
.A2(n_173),
.B1(n_169),
.B2(n_172),
.Y(n_4692)
);

CKINVDCx11_ASAP7_75t_R g4693 ( 
.A(n_4308),
.Y(n_4693)
);

NAND2xp5_ASAP7_75t_L g4694 ( 
.A(n_4639),
.B(n_4476),
.Y(n_4694)
);

AND2x2_ASAP7_75t_L g4695 ( 
.A(n_4647),
.B(n_4496),
.Y(n_4695)
);

AND2x4_ASAP7_75t_L g4696 ( 
.A(n_4631),
.B(n_4390),
.Y(n_4696)
);

AND2x2_ASAP7_75t_L g4697 ( 
.A(n_4526),
.B(n_4496),
.Y(n_4697)
);

AOI21xp5_ASAP7_75t_L g4698 ( 
.A1(n_4573),
.A2(n_4289),
.B(n_4375),
.Y(n_4698)
);

AND2x2_ASAP7_75t_L g4699 ( 
.A(n_4526),
.B(n_4498),
.Y(n_4699)
);

CKINVDCx9p33_ASAP7_75t_R g4700 ( 
.A(n_4538),
.Y(n_4700)
);

NOR2xp33_ASAP7_75t_L g4701 ( 
.A(n_4539),
.B(n_4474),
.Y(n_4701)
);

OA21x2_ASAP7_75t_L g4702 ( 
.A1(n_4641),
.A2(n_4489),
.B(n_4323),
.Y(n_4702)
);

AND2x4_ASAP7_75t_L g4703 ( 
.A(n_4631),
.B(n_4390),
.Y(n_4703)
);

INVx3_ASAP7_75t_L g4704 ( 
.A(n_4685),
.Y(n_4704)
);

INVxp67_ASAP7_75t_L g4705 ( 
.A(n_4579),
.Y(n_4705)
);

OAI22xp5_ASAP7_75t_L g4706 ( 
.A1(n_4559),
.A2(n_4390),
.B1(n_4347),
.B2(n_4300),
.Y(n_4706)
);

O2A1O1Ixp33_ASAP7_75t_L g4707 ( 
.A1(n_4672),
.A2(n_4442),
.B(n_4450),
.C(n_4432),
.Y(n_4707)
);

AND2x2_ASAP7_75t_L g4708 ( 
.A(n_4590),
.B(n_4628),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_L g4709 ( 
.A(n_4602),
.B(n_4305),
.Y(n_4709)
);

OR2x2_ASAP7_75t_L g4710 ( 
.A(n_4611),
.B(n_4469),
.Y(n_4710)
);

INVx2_ASAP7_75t_L g4711 ( 
.A(n_4536),
.Y(n_4711)
);

O2A1O1Ixp33_ASAP7_75t_L g4712 ( 
.A1(n_4555),
.A2(n_4380),
.B(n_4365),
.C(n_4325),
.Y(n_4712)
);

BUFx6f_ASAP7_75t_L g4713 ( 
.A(n_4568),
.Y(n_4713)
);

AND2x2_ASAP7_75t_L g4714 ( 
.A(n_4614),
.B(n_4502),
.Y(n_4714)
);

CKINVDCx5p33_ASAP7_75t_R g4715 ( 
.A(n_4540),
.Y(n_4715)
);

O2A1O1Ixp33_ASAP7_75t_L g4716 ( 
.A1(n_4595),
.A2(n_4346),
.B(n_4353),
.C(n_4352),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_L g4717 ( 
.A(n_4547),
.B(n_4345),
.Y(n_4717)
);

AND2x2_ASAP7_75t_L g4718 ( 
.A(n_4682),
.B(n_4466),
.Y(n_4718)
);

AND2x2_ASAP7_75t_L g4719 ( 
.A(n_4615),
.B(n_4368),
.Y(n_4719)
);

CKINVDCx20_ASAP7_75t_R g4720 ( 
.A(n_4544),
.Y(n_4720)
);

NAND2xp5_ASAP7_75t_L g4721 ( 
.A(n_4561),
.B(n_4328),
.Y(n_4721)
);

O2A1O1Ixp5_ASAP7_75t_L g4722 ( 
.A1(n_4665),
.A2(n_4486),
.B(n_4350),
.C(n_4351),
.Y(n_4722)
);

O2A1O1Ixp5_ASAP7_75t_L g4723 ( 
.A1(n_4574),
.A2(n_4303),
.B(n_4404),
.C(n_4288),
.Y(n_4723)
);

INVx2_ASAP7_75t_L g4724 ( 
.A(n_4519),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_4560),
.B(n_4475),
.Y(n_4725)
);

CKINVDCx5p33_ASAP7_75t_R g4726 ( 
.A(n_4571),
.Y(n_4726)
);

AND2x2_ASAP7_75t_L g4727 ( 
.A(n_4615),
.B(n_4477),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_L g4728 ( 
.A(n_4567),
.B(n_4420),
.Y(n_4728)
);

AOI21xp5_ASAP7_75t_SL g4729 ( 
.A1(n_4525),
.A2(n_4372),
.B(n_4302),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4522),
.Y(n_4730)
);

INVx1_ASAP7_75t_L g4731 ( 
.A(n_4529),
.Y(n_4731)
);

OA21x2_ASAP7_75t_L g4732 ( 
.A1(n_4591),
.A2(n_4619),
.B(n_4678),
.Y(n_4732)
);

OAI22xp5_ASAP7_75t_L g4733 ( 
.A1(n_4523),
.A2(n_4433),
.B1(n_4286),
.B2(n_4399),
.Y(n_4733)
);

HB1xp67_ASAP7_75t_L g4734 ( 
.A(n_4622),
.Y(n_4734)
);

AND2x2_ASAP7_75t_L g4735 ( 
.A(n_4531),
.B(n_4497),
.Y(n_4735)
);

AND2x2_ASAP7_75t_L g4736 ( 
.A(n_4531),
.B(n_4497),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4534),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4535),
.Y(n_4738)
);

OA21x2_ASAP7_75t_L g4739 ( 
.A1(n_4681),
.A2(n_4312),
.B(n_4462),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_L g4740 ( 
.A(n_4572),
.B(n_4425),
.Y(n_4740)
);

OR2x2_ASAP7_75t_L g4741 ( 
.A(n_4509),
.B(n_4478),
.Y(n_4741)
);

AND2x2_ASAP7_75t_L g4742 ( 
.A(n_4654),
.B(n_4497),
.Y(n_4742)
);

AND2x2_ASAP7_75t_L g4743 ( 
.A(n_4563),
.B(n_4484),
.Y(n_4743)
);

OA21x2_ASAP7_75t_L g4744 ( 
.A1(n_4691),
.A2(n_4480),
.B(n_4358),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4575),
.B(n_4484),
.Y(n_4745)
);

AOI21x1_ASAP7_75t_SL g4746 ( 
.A1(n_4504),
.A2(n_4320),
.B(n_4308),
.Y(n_4746)
);

OAI22xp5_ASAP7_75t_L g4747 ( 
.A1(n_4553),
.A2(n_4433),
.B1(n_4339),
.B2(n_4340),
.Y(n_4747)
);

NAND2xp5_ASAP7_75t_L g4748 ( 
.A(n_4541),
.B(n_4484),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4542),
.Y(n_4749)
);

AOI211xp5_ASAP7_75t_L g4750 ( 
.A1(n_4598),
.A2(n_4340),
.B(n_4320),
.C(n_4490),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4554),
.B(n_4422),
.Y(n_4751)
);

NOR2x1_ASAP7_75t_SL g4752 ( 
.A(n_4512),
.B(n_4604),
.Y(n_4752)
);

AND2x2_ASAP7_75t_L g4753 ( 
.A(n_4563),
.B(n_4372),
.Y(n_4753)
);

AND2x2_ASAP7_75t_L g4754 ( 
.A(n_4612),
.B(n_4453),
.Y(n_4754)
);

OAI22xp5_ASAP7_75t_L g4755 ( 
.A1(n_4609),
.A2(n_4322),
.B1(n_4400),
.B2(n_4438),
.Y(n_4755)
);

O2A1O1Ixp33_ASAP7_75t_L g4756 ( 
.A1(n_4608),
.A2(n_4421),
.B(n_4452),
.C(n_4383),
.Y(n_4756)
);

AND2x2_ASAP7_75t_L g4757 ( 
.A(n_4612),
.B(n_173),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_4586),
.Y(n_4758)
);

OAI22xp5_ASAP7_75t_L g4759 ( 
.A1(n_4620),
.A2(n_4364),
.B1(n_4426),
.B2(n_4443),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4588),
.Y(n_4760)
);

NAND2xp5_ASAP7_75t_L g4761 ( 
.A(n_4616),
.B(n_175),
.Y(n_4761)
);

A2O1A1Ixp33_ASAP7_75t_L g4762 ( 
.A1(n_4596),
.A2(n_178),
.B(n_175),
.C(n_176),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_L g4763 ( 
.A(n_4515),
.B(n_4683),
.Y(n_4763)
);

OAI22xp5_ASAP7_75t_L g4764 ( 
.A1(n_4564),
.A2(n_4355),
.B1(n_4386),
.B2(n_4401),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_L g4765 ( 
.A(n_4648),
.B(n_4650),
.Y(n_4765)
);

A2O1A1Ixp33_ASAP7_75t_L g4766 ( 
.A1(n_4587),
.A2(n_180),
.B(n_178),
.C(n_179),
.Y(n_4766)
);

O2A1O1Ixp33_ASAP7_75t_L g4767 ( 
.A1(n_4621),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_4767)
);

AND2x2_ASAP7_75t_L g4768 ( 
.A(n_4537),
.B(n_4578),
.Y(n_4768)
);

OR2x2_ASAP7_75t_L g4769 ( 
.A(n_4593),
.B(n_181),
.Y(n_4769)
);

NAND2xp5_ASAP7_75t_L g4770 ( 
.A(n_4655),
.B(n_4597),
.Y(n_4770)
);

AND2x2_ASAP7_75t_L g4771 ( 
.A(n_4585),
.B(n_182),
.Y(n_4771)
);

NAND2xp5_ASAP7_75t_L g4772 ( 
.A(n_4592),
.B(n_183),
.Y(n_4772)
);

O2A1O1Ixp33_ASAP7_75t_L g4773 ( 
.A1(n_4583),
.A2(n_189),
.B(n_186),
.C(n_187),
.Y(n_4773)
);

AND2x2_ASAP7_75t_L g4774 ( 
.A(n_4518),
.B(n_189),
.Y(n_4774)
);

OR2x2_ASAP7_75t_L g4775 ( 
.A(n_4640),
.B(n_190),
.Y(n_4775)
);

BUFx3_ASAP7_75t_L g4776 ( 
.A(n_4570),
.Y(n_4776)
);

INVxp67_ASAP7_75t_L g4777 ( 
.A(n_4613),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4646),
.Y(n_4778)
);

AOI21x1_ASAP7_75t_L g4779 ( 
.A1(n_4566),
.A2(n_4562),
.B(n_4552),
.Y(n_4779)
);

NOR2xp67_ASAP7_75t_L g4780 ( 
.A(n_4505),
.B(n_190),
.Y(n_4780)
);

AND2x4_ASAP7_75t_L g4781 ( 
.A(n_4687),
.B(n_4505),
.Y(n_4781)
);

OR2x2_ASAP7_75t_L g4782 ( 
.A(n_4577),
.B(n_191),
.Y(n_4782)
);

AOI21x1_ASAP7_75t_SL g4783 ( 
.A1(n_4556),
.A2(n_192),
.B(n_193),
.Y(n_4783)
);

AND2x2_ASAP7_75t_L g4784 ( 
.A(n_4551),
.B(n_192),
.Y(n_4784)
);

OAI22xp5_ASAP7_75t_L g4785 ( 
.A1(n_4667),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_L g4786 ( 
.A(n_4674),
.B(n_194),
.Y(n_4786)
);

HB1xp67_ASAP7_75t_L g4787 ( 
.A(n_4658),
.Y(n_4787)
);

OA22x2_ASAP7_75t_L g4788 ( 
.A1(n_4599),
.A2(n_200),
.B1(n_195),
.B2(n_196),
.Y(n_4788)
);

AOI21xp5_ASAP7_75t_SL g4789 ( 
.A1(n_4558),
.A2(n_196),
.B(n_200),
.Y(n_4789)
);

NAND2xp5_ASAP7_75t_L g4790 ( 
.A(n_4610),
.B(n_201),
.Y(n_4790)
);

OAI22xp5_ASAP7_75t_L g4791 ( 
.A1(n_4604),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_4791)
);

O2A1O1Ixp5_ASAP7_75t_L g4792 ( 
.A1(n_4508),
.A2(n_4514),
.B(n_4556),
.C(n_4510),
.Y(n_4792)
);

AOI21x1_ASAP7_75t_SL g4793 ( 
.A1(n_4550),
.A2(n_203),
.B(n_204),
.Y(n_4793)
);

AND2x2_ASAP7_75t_L g4794 ( 
.A(n_4580),
.B(n_205),
.Y(n_4794)
);

INVx2_ASAP7_75t_L g4795 ( 
.A(n_4652),
.Y(n_4795)
);

AND2x4_ASAP7_75t_L g4796 ( 
.A(n_4505),
.B(n_207),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4653),
.Y(n_4797)
);

AOI21x1_ASAP7_75t_SL g4798 ( 
.A1(n_4584),
.A2(n_208),
.B(n_209),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4660),
.Y(n_4799)
);

A2O1A1Ixp33_ASAP7_75t_L g4800 ( 
.A1(n_4548),
.A2(n_4546),
.B(n_4533),
.C(n_4649),
.Y(n_4800)
);

O2A1O1Ixp33_ASAP7_75t_L g4801 ( 
.A1(n_4689),
.A2(n_210),
.B(n_208),
.C(n_209),
.Y(n_4801)
);

OAI31xp33_ASAP7_75t_L g4802 ( 
.A1(n_4636),
.A2(n_214),
.A3(n_212),
.B(n_213),
.Y(n_4802)
);

OR2x2_ASAP7_75t_L g4803 ( 
.A(n_4669),
.B(n_212),
.Y(n_4803)
);

INVx3_ASAP7_75t_L g4804 ( 
.A(n_4673),
.Y(n_4804)
);

OA21x2_ASAP7_75t_L g4805 ( 
.A1(n_4624),
.A2(n_4643),
.B(n_4625),
.Y(n_4805)
);

NAND2xp5_ASAP7_75t_L g4806 ( 
.A(n_4532),
.B(n_213),
.Y(n_4806)
);

NOR2xp67_ASAP7_75t_L g4807 ( 
.A(n_4516),
.B(n_215),
.Y(n_4807)
);

HB1xp67_ASAP7_75t_L g4808 ( 
.A(n_4633),
.Y(n_4808)
);

AOI21x1_ASAP7_75t_SL g4809 ( 
.A1(n_4584),
.A2(n_215),
.B(n_216),
.Y(n_4809)
);

AOI21xp5_ASAP7_75t_SL g4810 ( 
.A1(n_4645),
.A2(n_216),
.B(n_217),
.Y(n_4810)
);

INVx2_ASAP7_75t_L g4811 ( 
.A(n_4684),
.Y(n_4811)
);

HB1xp67_ASAP7_75t_L g4812 ( 
.A(n_4690),
.Y(n_4812)
);

BUFx2_ASAP7_75t_L g4813 ( 
.A(n_4545),
.Y(n_4813)
);

AOI21xp5_ASAP7_75t_SL g4814 ( 
.A1(n_4516),
.A2(n_217),
.B(n_218),
.Y(n_4814)
);

CKINVDCx11_ASAP7_75t_R g4815 ( 
.A(n_4606),
.Y(n_4815)
);

AND2x4_ASAP7_75t_L g4816 ( 
.A(n_4632),
.B(n_218),
.Y(n_4816)
);

O2A1O1Ixp5_ASAP7_75t_L g4817 ( 
.A1(n_4635),
.A2(n_221),
.B(n_219),
.C(n_220),
.Y(n_4817)
);

O2A1O1Ixp33_ASAP7_75t_L g4818 ( 
.A1(n_4692),
.A2(n_223),
.B(n_219),
.C(n_220),
.Y(n_4818)
);

OAI22xp5_ASAP7_75t_L g4819 ( 
.A1(n_4677),
.A2(n_4651),
.B1(n_4679),
.B2(n_4506),
.Y(n_4819)
);

AOI21x1_ASAP7_75t_SL g4820 ( 
.A1(n_4680),
.A2(n_223),
.B(n_224),
.Y(n_4820)
);

OR2x2_ASAP7_75t_L g4821 ( 
.A(n_4589),
.B(n_225),
.Y(n_4821)
);

OR2x2_ASAP7_75t_L g4822 ( 
.A(n_4673),
.B(n_226),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_4673),
.Y(n_4823)
);

CKINVDCx12_ASAP7_75t_R g4824 ( 
.A(n_4530),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4569),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4569),
.Y(n_4826)
);

OAI22xp5_ASAP7_75t_L g4827 ( 
.A1(n_4642),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_4827)
);

AND2x2_ASAP7_75t_L g4828 ( 
.A(n_4607),
.B(n_4670),
.Y(n_4828)
);

O2A1O1Ixp33_ASAP7_75t_L g4829 ( 
.A1(n_4662),
.A2(n_230),
.B(n_227),
.C(n_229),
.Y(n_4829)
);

O2A1O1Ixp5_ASAP7_75t_L g4830 ( 
.A1(n_4517),
.A2(n_232),
.B(n_230),
.C(n_231),
.Y(n_4830)
);

AOI21x1_ASAP7_75t_SL g4831 ( 
.A1(n_4521),
.A2(n_4675),
.B(n_4657),
.Y(n_4831)
);

OR2x2_ASAP7_75t_L g4832 ( 
.A(n_4661),
.B(n_233),
.Y(n_4832)
);

A2O1A1Ixp33_ASAP7_75t_L g4833 ( 
.A1(n_4604),
.A2(n_236),
.B(n_234),
.C(n_235),
.Y(n_4833)
);

AND2x2_ASAP7_75t_L g4834 ( 
.A(n_4539),
.B(n_234),
.Y(n_4834)
);

AOI21xp5_ASAP7_75t_SL g4835 ( 
.A1(n_4517),
.A2(n_236),
.B(n_237),
.Y(n_4835)
);

NAND2xp5_ASAP7_75t_L g4836 ( 
.A(n_4688),
.B(n_4527),
.Y(n_4836)
);

AOI21xp5_ASAP7_75t_SL g4837 ( 
.A1(n_4557),
.A2(n_237),
.B(n_238),
.Y(n_4837)
);

NAND2xp5_ASAP7_75t_L g4838 ( 
.A(n_4594),
.B(n_239),
.Y(n_4838)
);

AND2x2_ASAP7_75t_L g4839 ( 
.A(n_4521),
.B(n_240),
.Y(n_4839)
);

NAND2xp5_ASAP7_75t_SL g4840 ( 
.A(n_4528),
.B(n_1674),
.Y(n_4840)
);

AND2x2_ASAP7_75t_L g4841 ( 
.A(n_4708),
.B(n_4549),
.Y(n_4841)
);

OR2x2_ASAP7_75t_L g4842 ( 
.A(n_4741),
.B(n_4686),
.Y(n_4842)
);

NAND2xp5_ASAP7_75t_L g4843 ( 
.A(n_4694),
.B(n_4594),
.Y(n_4843)
);

AND2x2_ASAP7_75t_L g4844 ( 
.A(n_4735),
.B(n_4528),
.Y(n_4844)
);

NOR2xp33_ASAP7_75t_R g4845 ( 
.A(n_4715),
.B(n_4582),
.Y(n_4845)
);

INVx8_ASAP7_75t_L g4846 ( 
.A(n_4796),
.Y(n_4846)
);

AND2x2_ASAP7_75t_L g4847 ( 
.A(n_4736),
.B(n_4565),
.Y(n_4847)
);

CKINVDCx5p33_ASAP7_75t_R g4848 ( 
.A(n_4815),
.Y(n_4848)
);

AOI211xp5_ASAP7_75t_L g4849 ( 
.A1(n_4819),
.A2(n_4644),
.B(n_4686),
.C(n_4623),
.Y(n_4849)
);

NAND2x1p5_ASAP7_75t_L g4850 ( 
.A(n_4704),
.B(n_4632),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_L g4851 ( 
.A(n_4705),
.B(n_4594),
.Y(n_4851)
);

AOI22xp33_ASAP7_75t_L g4852 ( 
.A1(n_4819),
.A2(n_4601),
.B1(n_4659),
.B2(n_4676),
.Y(n_4852)
);

AND2x2_ASAP7_75t_L g4853 ( 
.A(n_4704),
.B(n_4565),
.Y(n_4853)
);

OAI21x1_ASAP7_75t_L g4854 ( 
.A1(n_4805),
.A2(n_4513),
.B(n_4511),
.Y(n_4854)
);

AOI22xp33_ASAP7_75t_SL g4855 ( 
.A1(n_4706),
.A2(n_4752),
.B1(n_4836),
.B2(n_4794),
.Y(n_4855)
);

NAND3xp33_ASAP7_75t_SL g4856 ( 
.A(n_4792),
.B(n_4576),
.C(n_4581),
.Y(n_4856)
);

INVx2_ASAP7_75t_L g4857 ( 
.A(n_4695),
.Y(n_4857)
);

HB1xp67_ASAP7_75t_L g4858 ( 
.A(n_4734),
.Y(n_4858)
);

AO31x2_ASAP7_75t_L g4859 ( 
.A1(n_4751),
.A2(n_4760),
.A3(n_4778),
.B(n_4758),
.Y(n_4859)
);

INVx2_ASAP7_75t_L g4860 ( 
.A(n_4795),
.Y(n_4860)
);

OR2x6_ASAP7_75t_L g4861 ( 
.A(n_4729),
.B(n_4543),
.Y(n_4861)
);

CKINVDCx5p33_ASAP7_75t_R g4862 ( 
.A(n_4720),
.Y(n_4862)
);

NOR2xp33_ASAP7_75t_R g4863 ( 
.A(n_4824),
.B(n_4627),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4797),
.Y(n_4864)
);

NOR3xp33_ASAP7_75t_SL g4865 ( 
.A(n_4833),
.B(n_4626),
.C(n_4557),
.Y(n_4865)
);

NAND2xp5_ASAP7_75t_L g4866 ( 
.A(n_4709),
.B(n_4600),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4799),
.Y(n_4867)
);

NAND2xp33_ASAP7_75t_R g4868 ( 
.A(n_4726),
.B(n_241),
.Y(n_4868)
);

CKINVDCx5p33_ASAP7_75t_R g4869 ( 
.A(n_4700),
.Y(n_4869)
);

BUFx2_ASAP7_75t_L g4870 ( 
.A(n_4781),
.Y(n_4870)
);

CKINVDCx5p33_ASAP7_75t_R g4871 ( 
.A(n_4776),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_L g4872 ( 
.A(n_4749),
.B(n_4600),
.Y(n_4872)
);

AND4x1_ASAP7_75t_L g4873 ( 
.A(n_4814),
.B(n_4666),
.C(n_4507),
.D(n_4520),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_4730),
.Y(n_4874)
);

OR2x2_ASAP7_75t_L g4875 ( 
.A(n_4717),
.B(n_4711),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4731),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4737),
.Y(n_4877)
);

INVx2_ASAP7_75t_L g4878 ( 
.A(n_4732),
.Y(n_4878)
);

NOR2xp33_ASAP7_75t_R g4879 ( 
.A(n_4713),
.B(n_4671),
.Y(n_4879)
);

INVx2_ASAP7_75t_L g4880 ( 
.A(n_4732),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_4738),
.Y(n_4881)
);

INVx2_ASAP7_75t_L g4882 ( 
.A(n_4805),
.Y(n_4882)
);

AND2x2_ASAP7_75t_L g4883 ( 
.A(n_4719),
.B(n_4663),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4728),
.Y(n_4884)
);

NAND2xp33_ASAP7_75t_R g4885 ( 
.A(n_4816),
.B(n_241),
.Y(n_4885)
);

CKINVDCx5p33_ASAP7_75t_R g4886 ( 
.A(n_4713),
.Y(n_4886)
);

CKINVDCx16_ASAP7_75t_R g4887 ( 
.A(n_4713),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4724),
.Y(n_4888)
);

NOR2x1_ASAP7_75t_L g4889 ( 
.A(n_4781),
.B(n_4663),
.Y(n_4889)
);

NOR2xp33_ASAP7_75t_R g4890 ( 
.A(n_4828),
.B(n_4693),
.Y(n_4890)
);

HB1xp67_ASAP7_75t_L g4891 ( 
.A(n_4787),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4725),
.Y(n_4892)
);

OAI21xp5_ASAP7_75t_SL g4893 ( 
.A1(n_4800),
.A2(n_4686),
.B(n_4663),
.Y(n_4893)
);

NAND4xp25_ASAP7_75t_L g4894 ( 
.A(n_4767),
.B(n_4524),
.C(n_247),
.D(n_242),
.Y(n_4894)
);

AND2x2_ASAP7_75t_L g4895 ( 
.A(n_4742),
.B(n_4632),
.Y(n_4895)
);

INVx2_ASAP7_75t_L g4896 ( 
.A(n_4811),
.Y(n_4896)
);

AND2x2_ASAP7_75t_L g4897 ( 
.A(n_4823),
.B(n_4618),
.Y(n_4897)
);

OAI21x1_ASAP7_75t_L g4898 ( 
.A1(n_4740),
.A2(n_4617),
.B(n_4605),
.Y(n_4898)
);

NOR3xp33_ASAP7_75t_SL g4899 ( 
.A(n_4791),
.B(n_4637),
.C(n_4603),
.Y(n_4899)
);

CKINVDCx5p33_ASAP7_75t_R g4900 ( 
.A(n_4813),
.Y(n_4900)
);

AND2x2_ASAP7_75t_L g4901 ( 
.A(n_4753),
.B(n_4638),
.Y(n_4901)
);

AND2x2_ASAP7_75t_L g4902 ( 
.A(n_4768),
.B(n_4630),
.Y(n_4902)
);

AND2x2_ASAP7_75t_L g4903 ( 
.A(n_4743),
.B(n_4630),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4770),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4808),
.Y(n_4905)
);

O2A1O1Ixp33_ASAP7_75t_SL g4906 ( 
.A1(n_4763),
.A2(n_4668),
.B(n_4603),
.C(n_4637),
.Y(n_4906)
);

OR2x2_ASAP7_75t_L g4907 ( 
.A(n_4710),
.B(n_4600),
.Y(n_4907)
);

BUFx2_ASAP7_75t_L g4908 ( 
.A(n_4696),
.Y(n_4908)
);

BUFx3_ASAP7_75t_L g4909 ( 
.A(n_4804),
.Y(n_4909)
);

CKINVDCx20_ASAP7_75t_R g4910 ( 
.A(n_4821),
.Y(n_4910)
);

CKINVDCx14_ASAP7_75t_R g4911 ( 
.A(n_4839),
.Y(n_4911)
);

BUFx2_ASAP7_75t_L g4912 ( 
.A(n_4696),
.Y(n_4912)
);

AO31x2_ASAP7_75t_L g4913 ( 
.A1(n_4786),
.A2(n_4617),
.A3(n_4629),
.B(n_4605),
.Y(n_4913)
);

CKINVDCx16_ASAP7_75t_R g4914 ( 
.A(n_4816),
.Y(n_4914)
);

AND2x2_ASAP7_75t_L g4915 ( 
.A(n_4825),
.B(n_4826),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4812),
.Y(n_4916)
);

AND2x2_ASAP7_75t_L g4917 ( 
.A(n_4804),
.B(n_4703),
.Y(n_4917)
);

AND2x4_ASAP7_75t_L g4918 ( 
.A(n_4703),
.B(n_4656),
.Y(n_4918)
);

AOI22xp33_ASAP7_75t_L g4919 ( 
.A1(n_4698),
.A2(n_4664),
.B1(n_4634),
.B2(n_4629),
.Y(n_4919)
);

BUFx3_ASAP7_75t_L g4920 ( 
.A(n_4774),
.Y(n_4920)
);

BUFx8_ASAP7_75t_L g4921 ( 
.A(n_4796),
.Y(n_4921)
);

OAI22xp5_ASAP7_75t_L g4922 ( 
.A1(n_4750),
.A2(n_4634),
.B1(n_4656),
.B2(n_247),
.Y(n_4922)
);

INVx4_ASAP7_75t_L g4923 ( 
.A(n_4832),
.Y(n_4923)
);

HB1xp67_ASAP7_75t_L g4924 ( 
.A(n_4721),
.Y(n_4924)
);

OR2x2_ASAP7_75t_L g4925 ( 
.A(n_4765),
.B(n_4656),
.Y(n_4925)
);

NAND2xp5_ASAP7_75t_SL g4926 ( 
.A(n_4779),
.B(n_1674),
.Y(n_4926)
);

INVx2_ASAP7_75t_L g4927 ( 
.A(n_4727),
.Y(n_4927)
);

BUFx12f_ASAP7_75t_L g4928 ( 
.A(n_4822),
.Y(n_4928)
);

INVxp67_ASAP7_75t_L g4929 ( 
.A(n_4772),
.Y(n_4929)
);

BUFx2_ASAP7_75t_L g4930 ( 
.A(n_4718),
.Y(n_4930)
);

INVx2_ASAP7_75t_L g4931 ( 
.A(n_4699),
.Y(n_4931)
);

OR2x2_ASAP7_75t_L g4932 ( 
.A(n_4745),
.B(n_242),
.Y(n_4932)
);

NAND2xp33_ASAP7_75t_R g4933 ( 
.A(n_4834),
.B(n_243),
.Y(n_4933)
);

NAND2xp5_ASAP7_75t_L g4934 ( 
.A(n_4775),
.B(n_248),
.Y(n_4934)
);

NAND2xp5_ASAP7_75t_L g4935 ( 
.A(n_4748),
.B(n_248),
.Y(n_4935)
);

CKINVDCx16_ASAP7_75t_R g4936 ( 
.A(n_4701),
.Y(n_4936)
);

INVx1_ASAP7_75t_L g4937 ( 
.A(n_4803),
.Y(n_4937)
);

HB1xp67_ASAP7_75t_L g4938 ( 
.A(n_4782),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4790),
.Y(n_4939)
);

OAI21xp5_ASAP7_75t_L g4940 ( 
.A1(n_4722),
.A2(n_249),
.B(n_250),
.Y(n_4940)
);

HB1xp67_ASAP7_75t_L g4941 ( 
.A(n_4769),
.Y(n_4941)
);

INVx2_ASAP7_75t_L g4942 ( 
.A(n_4697),
.Y(n_4942)
);

NOR2xp33_ASAP7_75t_R g4943 ( 
.A(n_4806),
.B(n_249),
.Y(n_4943)
);

INVx1_ASAP7_75t_L g4944 ( 
.A(n_4761),
.Y(n_4944)
);

CKINVDCx5p33_ASAP7_75t_R g4945 ( 
.A(n_4771),
.Y(n_4945)
);

NAND2xp33_ASAP7_75t_R g4946 ( 
.A(n_4757),
.B(n_251),
.Y(n_4946)
);

CKINVDCx5p33_ASAP7_75t_R g4947 ( 
.A(n_4784),
.Y(n_4947)
);

CKINVDCx20_ASAP7_75t_R g4948 ( 
.A(n_4777),
.Y(n_4948)
);

AND2x4_ASAP7_75t_L g4949 ( 
.A(n_4754),
.B(n_254),
.Y(n_4949)
);

AOI21xp33_ASAP7_75t_L g4950 ( 
.A1(n_4712),
.A2(n_255),
.B(n_257),
.Y(n_4950)
);

OR2x2_ASAP7_75t_L g4951 ( 
.A(n_4714),
.B(n_258),
.Y(n_4951)
);

HB1xp67_ASAP7_75t_L g4952 ( 
.A(n_4780),
.Y(n_4952)
);

NAND2xp5_ASAP7_75t_L g4953 ( 
.A(n_4707),
.B(n_4716),
.Y(n_4953)
);

CKINVDCx5p33_ASAP7_75t_R g4954 ( 
.A(n_4838),
.Y(n_4954)
);

AND2x4_ASAP7_75t_L g4955 ( 
.A(n_4780),
.B(n_4807),
.Y(n_4955)
);

NAND2xp5_ASAP7_75t_L g4956 ( 
.A(n_4756),
.B(n_258),
.Y(n_4956)
);

INVx1_ASAP7_75t_SL g4957 ( 
.A(n_4840),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_4739),
.Y(n_4958)
);

OAI22xp5_ASAP7_75t_L g4959 ( 
.A1(n_4750),
.A2(n_262),
.B1(n_259),
.B2(n_261),
.Y(n_4959)
);

BUFx6f_ASAP7_75t_L g4960 ( 
.A(n_4739),
.Y(n_4960)
);

INVx2_ASAP7_75t_L g4961 ( 
.A(n_4744),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4744),
.Y(n_4962)
);

NOR2x1p5_ASAP7_75t_L g4963 ( 
.A(n_4831),
.B(n_263),
.Y(n_4963)
);

OR2x6_ASAP7_75t_L g4964 ( 
.A(n_4835),
.B(n_265),
.Y(n_4964)
);

AND2x2_ASAP7_75t_L g4965 ( 
.A(n_4702),
.B(n_265),
.Y(n_4965)
);

INVx1_ASAP7_75t_SL g4966 ( 
.A(n_4788),
.Y(n_4966)
);

AND2x4_ASAP7_75t_L g4967 ( 
.A(n_4807),
.B(n_266),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4702),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4723),
.Y(n_4969)
);

CKINVDCx5p33_ASAP7_75t_R g4970 ( 
.A(n_4837),
.Y(n_4970)
);

INVx1_ASAP7_75t_L g4971 ( 
.A(n_4830),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4764),
.Y(n_4972)
);

O2A1O1Ixp33_ASAP7_75t_SL g4973 ( 
.A1(n_4762),
.A2(n_269),
.B(n_267),
.C(n_268),
.Y(n_4973)
);

AOI22xp33_ASAP7_75t_L g4974 ( 
.A1(n_4802),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_4974)
);

INVx2_ASAP7_75t_L g4975 ( 
.A(n_4733),
.Y(n_4975)
);

INVx1_ASAP7_75t_L g4976 ( 
.A(n_4747),
.Y(n_4976)
);

AND2x4_ASAP7_75t_L g4977 ( 
.A(n_4746),
.B(n_271),
.Y(n_4977)
);

NAND2xp33_ASAP7_75t_R g4978 ( 
.A(n_4820),
.B(n_273),
.Y(n_4978)
);

AND2x2_ASAP7_75t_L g4979 ( 
.A(n_4747),
.B(n_273),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4864),
.Y(n_4980)
);

OA21x2_ASAP7_75t_L g4981 ( 
.A1(n_4962),
.A2(n_4817),
.B(n_4766),
.Y(n_4981)
);

INVx2_ASAP7_75t_L g4982 ( 
.A(n_4878),
.Y(n_4982)
);

INVx1_ASAP7_75t_L g4983 ( 
.A(n_4867),
.Y(n_4983)
);

BUFx2_ASAP7_75t_L g4984 ( 
.A(n_4889),
.Y(n_4984)
);

INVx2_ASAP7_75t_L g4985 ( 
.A(n_4880),
.Y(n_4985)
);

OR2x2_ASAP7_75t_L g4986 ( 
.A(n_4859),
.B(n_4785),
.Y(n_4986)
);

HB1xp67_ASAP7_75t_L g4987 ( 
.A(n_4882),
.Y(n_4987)
);

OAI211xp5_ASAP7_75t_SL g4988 ( 
.A1(n_4953),
.A2(n_4802),
.B(n_4773),
.C(n_4801),
.Y(n_4988)
);

AO21x2_ASAP7_75t_L g4989 ( 
.A1(n_4968),
.A2(n_4965),
.B(n_4958),
.Y(n_4989)
);

INVx1_ASAP7_75t_L g4990 ( 
.A(n_4874),
.Y(n_4990)
);

NAND3xp33_ASAP7_75t_L g4991 ( 
.A(n_4873),
.B(n_4829),
.C(n_4818),
.Y(n_4991)
);

AO21x2_ASAP7_75t_L g4992 ( 
.A1(n_4961),
.A2(n_4810),
.B(n_4789),
.Y(n_4992)
);

INVx3_ASAP7_75t_L g4993 ( 
.A(n_4960),
.Y(n_4993)
);

INVxp67_ASAP7_75t_SL g4994 ( 
.A(n_4952),
.Y(n_4994)
);

INVx3_ASAP7_75t_L g4995 ( 
.A(n_4960),
.Y(n_4995)
);

AND2x2_ASAP7_75t_L g4996 ( 
.A(n_4908),
.B(n_4827),
.Y(n_4996)
);

INVx1_ASAP7_75t_SL g4997 ( 
.A(n_4879),
.Y(n_4997)
);

INVx2_ASAP7_75t_L g4998 ( 
.A(n_4960),
.Y(n_4998)
);

CKINVDCx5p33_ASAP7_75t_R g4999 ( 
.A(n_4868),
.Y(n_4999)
);

AND2x2_ASAP7_75t_L g5000 ( 
.A(n_4912),
.B(n_4827),
.Y(n_5000)
);

BUFx3_ASAP7_75t_L g5001 ( 
.A(n_4921),
.Y(n_5001)
);

BUFx2_ASAP7_75t_L g5002 ( 
.A(n_4889),
.Y(n_5002)
);

OR2x6_ASAP7_75t_L g5003 ( 
.A(n_4861),
.B(n_4755),
.Y(n_5003)
);

NAND2xp5_ASAP7_75t_L g5004 ( 
.A(n_4969),
.B(n_4972),
.Y(n_5004)
);

BUFx2_ASAP7_75t_L g5005 ( 
.A(n_4870),
.Y(n_5005)
);

INVxp67_ASAP7_75t_SL g5006 ( 
.A(n_4955),
.Y(n_5006)
);

OAI211xp5_ASAP7_75t_L g5007 ( 
.A1(n_4893),
.A2(n_4849),
.B(n_4940),
.C(n_4894),
.Y(n_5007)
);

OAI21xp5_ASAP7_75t_L g5008 ( 
.A1(n_4893),
.A2(n_4755),
.B(n_4759),
.Y(n_5008)
);

AND2x2_ASAP7_75t_L g5009 ( 
.A(n_4917),
.B(n_4759),
.Y(n_5009)
);

OAI221xp5_ASAP7_75t_L g5010 ( 
.A1(n_4855),
.A2(n_4793),
.B1(n_4798),
.B2(n_4809),
.C(n_4783),
.Y(n_5010)
);

AOI21xp5_ASAP7_75t_L g5011 ( 
.A1(n_4959),
.A2(n_274),
.B(n_275),
.Y(n_5011)
);

INVx2_ASAP7_75t_L g5012 ( 
.A(n_4860),
.Y(n_5012)
);

BUFx2_ASAP7_75t_SL g5013 ( 
.A(n_4955),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4876),
.Y(n_5014)
);

OA21x2_ASAP7_75t_L g5015 ( 
.A1(n_4854),
.A2(n_275),
.B(n_277),
.Y(n_5015)
);

AO21x2_ASAP7_75t_L g5016 ( 
.A1(n_4926),
.A2(n_278),
.B(n_279),
.Y(n_5016)
);

AO21x2_ASAP7_75t_L g5017 ( 
.A1(n_4956),
.A2(n_279),
.B(n_280),
.Y(n_5017)
);

INVx3_ASAP7_75t_L g5018 ( 
.A(n_4850),
.Y(n_5018)
);

AND2x2_ASAP7_75t_L g5019 ( 
.A(n_4895),
.B(n_281),
.Y(n_5019)
);

INVx1_ASAP7_75t_L g5020 ( 
.A(n_4877),
.Y(n_5020)
);

AOI22xp33_ASAP7_75t_L g5021 ( 
.A1(n_4856),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_5021)
);

INVx1_ASAP7_75t_L g5022 ( 
.A(n_4881),
.Y(n_5022)
);

AO21x2_ASAP7_75t_L g5023 ( 
.A1(n_4950),
.A2(n_282),
.B(n_284),
.Y(n_5023)
);

OR2x2_ASAP7_75t_L g5024 ( 
.A(n_4875),
.B(n_285),
.Y(n_5024)
);

HB1xp67_ASAP7_75t_L g5025 ( 
.A(n_4858),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_4904),
.Y(n_5026)
);

AND2x2_ASAP7_75t_L g5027 ( 
.A(n_4924),
.B(n_286),
.Y(n_5027)
);

NAND2xp5_ASAP7_75t_L g5028 ( 
.A(n_4976),
.B(n_286),
.Y(n_5028)
);

OA21x2_ASAP7_75t_L g5029 ( 
.A1(n_4898),
.A2(n_287),
.B(n_288),
.Y(n_5029)
);

AND2x2_ASAP7_75t_L g5030 ( 
.A(n_4942),
.B(n_4918),
.Y(n_5030)
);

INVx2_ASAP7_75t_L g5031 ( 
.A(n_4927),
.Y(n_5031)
);

INVx1_ASAP7_75t_L g5032 ( 
.A(n_4888),
.Y(n_5032)
);

AND2x2_ASAP7_75t_L g5033 ( 
.A(n_4918),
.B(n_289),
.Y(n_5033)
);

AO21x2_ASAP7_75t_L g5034 ( 
.A1(n_4943),
.A2(n_290),
.B(n_291),
.Y(n_5034)
);

OR2x2_ASAP7_75t_L g5035 ( 
.A(n_4859),
.B(n_292),
.Y(n_5035)
);

OA21x2_ASAP7_75t_L g5036 ( 
.A1(n_4971),
.A2(n_292),
.B(n_295),
.Y(n_5036)
);

AOI21x1_ASAP7_75t_L g5037 ( 
.A1(n_4861),
.A2(n_295),
.B(n_296),
.Y(n_5037)
);

AOI21xp33_ASAP7_75t_L g5038 ( 
.A1(n_4978),
.A2(n_4922),
.B(n_4964),
.Y(n_5038)
);

OR2x2_ASAP7_75t_L g5039 ( 
.A(n_4859),
.B(n_296),
.Y(n_5039)
);

OR2x6_ASAP7_75t_L g5040 ( 
.A(n_4861),
.B(n_297),
.Y(n_5040)
);

INVx2_ASAP7_75t_L g5041 ( 
.A(n_4913),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_4938),
.Y(n_5042)
);

BUFx2_ASAP7_75t_L g5043 ( 
.A(n_4890),
.Y(n_5043)
);

INVx5_ASAP7_75t_L g5044 ( 
.A(n_4964),
.Y(n_5044)
);

OAI321xp33_ASAP7_75t_L g5045 ( 
.A1(n_4894),
.A2(n_298),
.A3(n_299),
.B1(n_300),
.B2(n_301),
.C(n_302),
.Y(n_5045)
);

AO21x2_ASAP7_75t_L g5046 ( 
.A1(n_4873),
.A2(n_299),
.B(n_303),
.Y(n_5046)
);

AO21x2_ASAP7_75t_L g5047 ( 
.A1(n_4935),
.A2(n_305),
.B(n_306),
.Y(n_5047)
);

INVxp67_ASAP7_75t_L g5048 ( 
.A(n_4885),
.Y(n_5048)
);

AND2x2_ASAP7_75t_L g5049 ( 
.A(n_4913),
.B(n_305),
.Y(n_5049)
);

INVx2_ASAP7_75t_L g5050 ( 
.A(n_4913),
.Y(n_5050)
);

OAI22xp33_ASAP7_75t_L g5051 ( 
.A1(n_4964),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_5051)
);

AO21x2_ASAP7_75t_L g5052 ( 
.A1(n_4934),
.A2(n_307),
.B(n_309),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4941),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_4937),
.Y(n_5054)
);

OR2x6_ASAP7_75t_L g5055 ( 
.A(n_4977),
.B(n_309),
.Y(n_5055)
);

BUFx6f_ASAP7_75t_L g5056 ( 
.A(n_4886),
.Y(n_5056)
);

OAI21xp5_ASAP7_75t_L g5057 ( 
.A1(n_4865),
.A2(n_312),
.B(n_313),
.Y(n_5057)
);

INVx2_ASAP7_75t_L g5058 ( 
.A(n_4896),
.Y(n_5058)
);

AND2x2_ASAP7_75t_L g5059 ( 
.A(n_4847),
.B(n_312),
.Y(n_5059)
);

OA21x2_ASAP7_75t_L g5060 ( 
.A1(n_4975),
.A2(n_313),
.B(n_316),
.Y(n_5060)
);

BUFx3_ASAP7_75t_L g5061 ( 
.A(n_4921),
.Y(n_5061)
);

INVx2_ASAP7_75t_L g5062 ( 
.A(n_4905),
.Y(n_5062)
);

BUFx3_ASAP7_75t_L g5063 ( 
.A(n_4846),
.Y(n_5063)
);

NAND2xp5_ASAP7_75t_L g5064 ( 
.A(n_4939),
.B(n_317),
.Y(n_5064)
);

AO21x2_ASAP7_75t_L g5065 ( 
.A1(n_4979),
.A2(n_317),
.B(n_318),
.Y(n_5065)
);

AND2x2_ASAP7_75t_L g5066 ( 
.A(n_4930),
.B(n_318),
.Y(n_5066)
);

INVx2_ASAP7_75t_L g5067 ( 
.A(n_4916),
.Y(n_5067)
);

INVx1_ASAP7_75t_L g5068 ( 
.A(n_4891),
.Y(n_5068)
);

NAND2xp5_ASAP7_75t_L g5069 ( 
.A(n_4944),
.B(n_321),
.Y(n_5069)
);

INVxp67_ASAP7_75t_SL g5070 ( 
.A(n_4946),
.Y(n_5070)
);

AND2x2_ASAP7_75t_L g5071 ( 
.A(n_4844),
.B(n_4857),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_4929),
.B(n_321),
.Y(n_5072)
);

INVxp67_ASAP7_75t_SL g5073 ( 
.A(n_4910),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_4884),
.Y(n_5074)
);

OA21x2_ASAP7_75t_L g5075 ( 
.A1(n_4919),
.A2(n_322),
.B(n_323),
.Y(n_5075)
);

AO21x2_ASAP7_75t_L g5076 ( 
.A1(n_4863),
.A2(n_323),
.B(n_324),
.Y(n_5076)
);

INVx1_ASAP7_75t_SL g5077 ( 
.A(n_4887),
.Y(n_5077)
);

OA21x2_ASAP7_75t_L g5078 ( 
.A1(n_4966),
.A2(n_325),
.B(n_326),
.Y(n_5078)
);

AND2x2_ASAP7_75t_L g5079 ( 
.A(n_4853),
.B(n_327),
.Y(n_5079)
);

AO21x1_ASAP7_75t_SL g5080 ( 
.A1(n_4852),
.A2(n_328),
.B(n_330),
.Y(n_5080)
);

OR2x2_ASAP7_75t_L g5081 ( 
.A(n_4842),
.B(n_333),
.Y(n_5081)
);

BUFx3_ASAP7_75t_L g5082 ( 
.A(n_4846),
.Y(n_5082)
);

INVx2_ASAP7_75t_L g5083 ( 
.A(n_4907),
.Y(n_5083)
);

OA21x2_ASAP7_75t_L g5084 ( 
.A1(n_4892),
.A2(n_334),
.B(n_335),
.Y(n_5084)
);

AND2x2_ASAP7_75t_L g5085 ( 
.A(n_4903),
.B(n_335),
.Y(n_5085)
);

OR2x2_ASAP7_75t_L g5086 ( 
.A(n_5004),
.B(n_4951),
.Y(n_5086)
);

AND2x2_ASAP7_75t_L g5087 ( 
.A(n_5013),
.B(n_4911),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_5025),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_5025),
.Y(n_5089)
);

AOI22xp33_ASAP7_75t_SL g5090 ( 
.A1(n_5070),
.A2(n_4970),
.B1(n_4936),
.B2(n_4948),
.Y(n_5090)
);

HB1xp67_ASAP7_75t_L g5091 ( 
.A(n_4987),
.Y(n_5091)
);

HB1xp67_ASAP7_75t_L g5092 ( 
.A(n_4987),
.Y(n_5092)
);

AND2x2_ASAP7_75t_L g5093 ( 
.A(n_5009),
.B(n_4909),
.Y(n_5093)
);

INVx1_ASAP7_75t_L g5094 ( 
.A(n_4980),
.Y(n_5094)
);

HB1xp67_ASAP7_75t_L g5095 ( 
.A(n_5035),
.Y(n_5095)
);

AND2x2_ASAP7_75t_L g5096 ( 
.A(n_5006),
.B(n_4914),
.Y(n_5096)
);

OR2x2_ASAP7_75t_L g5097 ( 
.A(n_5042),
.B(n_4932),
.Y(n_5097)
);

AND2x2_ASAP7_75t_L g5098 ( 
.A(n_5009),
.B(n_4923),
.Y(n_5098)
);

AND2x2_ASAP7_75t_L g5099 ( 
.A(n_5030),
.B(n_4923),
.Y(n_5099)
);

HB1xp67_ASAP7_75t_L g5100 ( 
.A(n_5035),
.Y(n_5100)
);

AND2x2_ASAP7_75t_L g5101 ( 
.A(n_5030),
.B(n_4901),
.Y(n_5101)
);

HB1xp67_ASAP7_75t_L g5102 ( 
.A(n_5039),
.Y(n_5102)
);

INVx2_ASAP7_75t_L g5103 ( 
.A(n_5005),
.Y(n_5103)
);

NAND2xp5_ASAP7_75t_L g5104 ( 
.A(n_5049),
.B(n_4957),
.Y(n_5104)
);

AND2x2_ASAP7_75t_L g5105 ( 
.A(n_5063),
.B(n_4883),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_4983),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_4990),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_5014),
.Y(n_5108)
);

INVx1_ASAP7_75t_L g5109 ( 
.A(n_5020),
.Y(n_5109)
);

BUFx2_ASAP7_75t_L g5110 ( 
.A(n_4984),
.Y(n_5110)
);

NAND2x1_ASAP7_75t_L g5111 ( 
.A(n_5002),
.B(n_4841),
.Y(n_5111)
);

AND2x2_ASAP7_75t_L g5112 ( 
.A(n_5018),
.B(n_4931),
.Y(n_5112)
);

INVx2_ASAP7_75t_L g5113 ( 
.A(n_4993),
.Y(n_5113)
);

INVx1_ASAP7_75t_L g5114 ( 
.A(n_5022),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_5039),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_4994),
.Y(n_5116)
);

INVx2_ASAP7_75t_L g5117 ( 
.A(n_4993),
.Y(n_5117)
);

AND2x2_ASAP7_75t_L g5118 ( 
.A(n_5063),
.B(n_4915),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_5062),
.Y(n_5119)
);

INVx1_ASAP7_75t_L g5120 ( 
.A(n_5062),
.Y(n_5120)
);

AND2x2_ASAP7_75t_L g5121 ( 
.A(n_5082),
.B(n_4902),
.Y(n_5121)
);

INVx2_ASAP7_75t_L g5122 ( 
.A(n_4993),
.Y(n_5122)
);

INVx1_ASAP7_75t_L g5123 ( 
.A(n_5067),
.Y(n_5123)
);

NAND2x1p5_ASAP7_75t_L g5124 ( 
.A(n_5044),
.B(n_4977),
.Y(n_5124)
);

INVx2_ASAP7_75t_L g5125 ( 
.A(n_4995),
.Y(n_5125)
);

AND2x4_ASAP7_75t_SL g5126 ( 
.A(n_5040),
.B(n_4899),
.Y(n_5126)
);

NAND2xp5_ASAP7_75t_L g5127 ( 
.A(n_5049),
.B(n_4967),
.Y(n_5127)
);

NOR2x1_ASAP7_75t_L g5128 ( 
.A(n_5046),
.B(n_4963),
.Y(n_5128)
);

OR2x2_ASAP7_75t_L g5129 ( 
.A(n_5053),
.B(n_4866),
.Y(n_5129)
);

INVx1_ASAP7_75t_L g5130 ( 
.A(n_5067),
.Y(n_5130)
);

NAND2xp5_ASAP7_75t_L g5131 ( 
.A(n_5017),
.B(n_5046),
.Y(n_5131)
);

OR2x2_ASAP7_75t_L g5132 ( 
.A(n_5083),
.B(n_4925),
.Y(n_5132)
);

AND2x2_ASAP7_75t_L g5133 ( 
.A(n_5082),
.B(n_4869),
.Y(n_5133)
);

INVx2_ASAP7_75t_L g5134 ( 
.A(n_4995),
.Y(n_5134)
);

NAND2xp5_ASAP7_75t_L g5135 ( 
.A(n_5017),
.B(n_4967),
.Y(n_5135)
);

INVx2_ASAP7_75t_L g5136 ( 
.A(n_4995),
.Y(n_5136)
);

NAND2xp5_ASAP7_75t_L g5137 ( 
.A(n_5008),
.B(n_4949),
.Y(n_5137)
);

INVxp67_ASAP7_75t_L g5138 ( 
.A(n_5078),
.Y(n_5138)
);

INVx3_ASAP7_75t_L g5139 ( 
.A(n_5044),
.Y(n_5139)
);

OR2x2_ASAP7_75t_L g5140 ( 
.A(n_5083),
.B(n_4843),
.Y(n_5140)
);

CKINVDCx20_ASAP7_75t_R g5141 ( 
.A(n_4999),
.Y(n_5141)
);

BUFx4f_ASAP7_75t_L g5142 ( 
.A(n_5056),
.Y(n_5142)
);

INVx4_ASAP7_75t_L g5143 ( 
.A(n_5001),
.Y(n_5143)
);

AND2x2_ASAP7_75t_L g5144 ( 
.A(n_4996),
.B(n_4897),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_5032),
.Y(n_5145)
);

OR2x2_ASAP7_75t_L g5146 ( 
.A(n_5068),
.B(n_4872),
.Y(n_5146)
);

AND2x4_ASAP7_75t_L g5147 ( 
.A(n_5018),
.B(n_4920),
.Y(n_5147)
);

INVx2_ASAP7_75t_SL g5148 ( 
.A(n_5044),
.Y(n_5148)
);

OR2x2_ASAP7_75t_L g5149 ( 
.A(n_4996),
.B(n_4851),
.Y(n_5149)
);

AOI22xp33_ASAP7_75t_L g5150 ( 
.A1(n_4991),
.A2(n_4974),
.B1(n_4928),
.B2(n_4954),
.Y(n_5150)
);

AND2x2_ASAP7_75t_L g5151 ( 
.A(n_5000),
.B(n_4900),
.Y(n_5151)
);

INVx5_ASAP7_75t_L g5152 ( 
.A(n_5040),
.Y(n_5152)
);

AOI22xp5_ASAP7_75t_L g5153 ( 
.A1(n_5007),
.A2(n_4849),
.B1(n_4933),
.B2(n_4973),
.Y(n_5153)
);

NAND2xp5_ASAP7_75t_L g5154 ( 
.A(n_5078),
.B(n_4949),
.Y(n_5154)
);

OR2x2_ASAP7_75t_L g5155 ( 
.A(n_5000),
.B(n_5024),
.Y(n_5155)
);

INVx2_ASAP7_75t_L g5156 ( 
.A(n_5044),
.Y(n_5156)
);

INVx2_ASAP7_75t_L g5157 ( 
.A(n_4998),
.Y(n_5157)
);

INVx2_ASAP7_75t_L g5158 ( 
.A(n_4998),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_5054),
.Y(n_5159)
);

INVx2_ASAP7_75t_L g5160 ( 
.A(n_5029),
.Y(n_5160)
);

AND2x2_ASAP7_75t_L g5161 ( 
.A(n_5071),
.B(n_5077),
.Y(n_5161)
);

OAI222xp33_ASAP7_75t_L g5162 ( 
.A1(n_5048),
.A2(n_4947),
.B1(n_4945),
.B2(n_4871),
.C1(n_4848),
.C2(n_4862),
.Y(n_5162)
);

OAI31xp33_ASAP7_75t_SL g5163 ( 
.A1(n_5128),
.A2(n_5038),
.A3(n_5090),
.B(n_4988),
.Y(n_5163)
);

BUFx2_ASAP7_75t_L g5164 ( 
.A(n_5141),
.Y(n_5164)
);

NOR2x2_ASAP7_75t_L g5165 ( 
.A(n_5103),
.B(n_5003),
.Y(n_5165)
);

INVx1_ASAP7_75t_L g5166 ( 
.A(n_5091),
.Y(n_5166)
);

AND2x2_ASAP7_75t_L g5167 ( 
.A(n_5087),
.B(n_5043),
.Y(n_5167)
);

CKINVDCx16_ASAP7_75t_R g5168 ( 
.A(n_5141),
.Y(n_5168)
);

OR2x2_ASAP7_75t_L g5169 ( 
.A(n_5155),
.B(n_4986),
.Y(n_5169)
);

NAND2xp5_ASAP7_75t_L g5170 ( 
.A(n_5153),
.B(n_5096),
.Y(n_5170)
);

OAI31xp33_ASAP7_75t_L g5171 ( 
.A1(n_5131),
.A2(n_5010),
.A3(n_5051),
.B(n_5021),
.Y(n_5171)
);

OAI22xp5_ASAP7_75t_L g5172 ( 
.A1(n_5090),
.A2(n_4999),
.B1(n_5003),
.B2(n_5124),
.Y(n_5172)
);

BUFx2_ASAP7_75t_L g5173 ( 
.A(n_5124),
.Y(n_5173)
);

OR2x6_ASAP7_75t_L g5174 ( 
.A(n_5148),
.B(n_5040),
.Y(n_5174)
);

OA21x2_ASAP7_75t_L g5175 ( 
.A1(n_5138),
.A2(n_5050),
.B(n_5041),
.Y(n_5175)
);

AO21x1_ASAP7_75t_L g5176 ( 
.A1(n_5095),
.A2(n_4986),
.B(n_5051),
.Y(n_5176)
);

OAI221xp5_ASAP7_75t_L g5177 ( 
.A1(n_5150),
.A2(n_5021),
.B1(n_5057),
.B2(n_5003),
.C(n_5040),
.Y(n_5177)
);

AND2x2_ASAP7_75t_L g5178 ( 
.A(n_5096),
.B(n_5071),
.Y(n_5178)
);

AOI221xp5_ASAP7_75t_L g5179 ( 
.A1(n_5095),
.A2(n_5045),
.B1(n_5011),
.B2(n_5034),
.C(n_5076),
.Y(n_5179)
);

AND2x4_ASAP7_75t_L g5180 ( 
.A(n_5152),
.B(n_5001),
.Y(n_5180)
);

INVxp67_ASAP7_75t_L g5181 ( 
.A(n_5151),
.Y(n_5181)
);

NAND4xp25_ASAP7_75t_L g5182 ( 
.A(n_5150),
.B(n_5115),
.C(n_5143),
.D(n_5138),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_5091),
.Y(n_5183)
);

INVx1_ASAP7_75t_L g5184 ( 
.A(n_5092),
.Y(n_5184)
);

AND2x4_ASAP7_75t_SL g5185 ( 
.A(n_5143),
.B(n_5056),
.Y(n_5185)
);

INVx2_ASAP7_75t_L g5186 ( 
.A(n_5139),
.Y(n_5186)
);

INVx2_ASAP7_75t_L g5187 ( 
.A(n_5139),
.Y(n_5187)
);

OR2x2_ASAP7_75t_L g5188 ( 
.A(n_5149),
.B(n_4981),
.Y(n_5188)
);

OAI22xp5_ASAP7_75t_L g5189 ( 
.A1(n_5152),
.A2(n_5003),
.B1(n_5055),
.B2(n_4981),
.Y(n_5189)
);

NOR4xp25_ASAP7_75t_SL g5190 ( 
.A(n_5110),
.B(n_4906),
.C(n_5073),
.D(n_5076),
.Y(n_5190)
);

AND2x4_ASAP7_75t_SL g5191 ( 
.A(n_5143),
.B(n_5056),
.Y(n_5191)
);

NAND3xp33_ASAP7_75t_L g5192 ( 
.A(n_5100),
.B(n_5078),
.C(n_5036),
.Y(n_5192)
);

AOI22xp33_ASAP7_75t_L g5193 ( 
.A1(n_5152),
.A2(n_4981),
.B1(n_4992),
.B2(n_5015),
.Y(n_5193)
);

NAND4xp25_ASAP7_75t_L g5194 ( 
.A(n_5135),
.B(n_5028),
.C(n_5072),
.D(n_5061),
.Y(n_5194)
);

OAI221xp5_ASAP7_75t_L g5195 ( 
.A1(n_5111),
.A2(n_5055),
.B1(n_4997),
.B2(n_5018),
.C(n_5061),
.Y(n_5195)
);

AOI22xp33_ASAP7_75t_L g5196 ( 
.A1(n_5152),
.A2(n_4992),
.B1(n_5015),
.B2(n_4989),
.Y(n_5196)
);

AOI22xp33_ASAP7_75t_SL g5197 ( 
.A1(n_5100),
.A2(n_5034),
.B1(n_5036),
.B2(n_5055),
.Y(n_5197)
);

BUFx2_ASAP7_75t_L g5198 ( 
.A(n_5139),
.Y(n_5198)
);

AO21x2_ASAP7_75t_L g5199 ( 
.A1(n_5102),
.A2(n_5050),
.B(n_5041),
.Y(n_5199)
);

AOI21xp5_ASAP7_75t_L g5200 ( 
.A1(n_5162),
.A2(n_5055),
.B(n_5036),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_5092),
.Y(n_5201)
);

OAI22xp5_ASAP7_75t_L g5202 ( 
.A1(n_5154),
.A2(n_5075),
.B1(n_5015),
.B2(n_5084),
.Y(n_5202)
);

OA21x2_ASAP7_75t_L g5203 ( 
.A1(n_5160),
.A2(n_4985),
.B(n_4982),
.Y(n_5203)
);

AOI22xp33_ASAP7_75t_L g5204 ( 
.A1(n_5126),
.A2(n_4989),
.B1(n_5080),
.B2(n_5075),
.Y(n_5204)
);

OR2x2_ASAP7_75t_L g5205 ( 
.A(n_5116),
.B(n_5026),
.Y(n_5205)
);

INVxp67_ASAP7_75t_SL g5206 ( 
.A(n_5098),
.Y(n_5206)
);

INVx2_ASAP7_75t_L g5207 ( 
.A(n_5148),
.Y(n_5207)
);

BUFx2_ASAP7_75t_L g5208 ( 
.A(n_5147),
.Y(n_5208)
);

AOI211xp5_ASAP7_75t_L g5209 ( 
.A1(n_5162),
.A2(n_5027),
.B(n_5064),
.C(n_5069),
.Y(n_5209)
);

INVx1_ASAP7_75t_L g5210 ( 
.A(n_5088),
.Y(n_5210)
);

AND2x2_ASAP7_75t_L g5211 ( 
.A(n_5144),
.B(n_5019),
.Y(n_5211)
);

INVx2_ASAP7_75t_L g5212 ( 
.A(n_5161),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_5176),
.Y(n_5213)
);

INVx2_ASAP7_75t_L g5214 ( 
.A(n_5164),
.Y(n_5214)
);

AND2x2_ASAP7_75t_L g5215 ( 
.A(n_5167),
.B(n_5099),
.Y(n_5215)
);

AND2x2_ASAP7_75t_L g5216 ( 
.A(n_5178),
.B(n_5103),
.Y(n_5216)
);

BUFx2_ASAP7_75t_L g5217 ( 
.A(n_5168),
.Y(n_5217)
);

OR2x2_ASAP7_75t_L g5218 ( 
.A(n_5192),
.B(n_5169),
.Y(n_5218)
);

AND2x2_ASAP7_75t_L g5219 ( 
.A(n_5208),
.B(n_5147),
.Y(n_5219)
);

AND2x4_ASAP7_75t_L g5220 ( 
.A(n_5198),
.B(n_5156),
.Y(n_5220)
);

INVx3_ASAP7_75t_L g5221 ( 
.A(n_5180),
.Y(n_5221)
);

AND2x2_ASAP7_75t_L g5222 ( 
.A(n_5180),
.B(n_5211),
.Y(n_5222)
);

INVx1_ASAP7_75t_L g5223 ( 
.A(n_5166),
.Y(n_5223)
);

INVx2_ASAP7_75t_SL g5224 ( 
.A(n_5185),
.Y(n_5224)
);

NOR3xp33_ASAP7_75t_L g5225 ( 
.A(n_5182),
.B(n_5156),
.C(n_5102),
.Y(n_5225)
);

NAND2xp5_ASAP7_75t_L g5226 ( 
.A(n_5171),
.B(n_5127),
.Y(n_5226)
);

INVx1_ASAP7_75t_L g5227 ( 
.A(n_5183),
.Y(n_5227)
);

NAND2xp5_ASAP7_75t_L g5228 ( 
.A(n_5171),
.B(n_5137),
.Y(n_5228)
);

INVx2_ASAP7_75t_L g5229 ( 
.A(n_5174),
.Y(n_5229)
);

INVx4_ASAP7_75t_L g5230 ( 
.A(n_5191),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_5184),
.Y(n_5231)
);

AND2x2_ASAP7_75t_L g5232 ( 
.A(n_5174),
.B(n_5147),
.Y(n_5232)
);

HB1xp67_ASAP7_75t_L g5233 ( 
.A(n_5174),
.Y(n_5233)
);

INVx4_ASAP7_75t_L g5234 ( 
.A(n_5173),
.Y(n_5234)
);

AND2x4_ASAP7_75t_L g5235 ( 
.A(n_5192),
.B(n_5113),
.Y(n_5235)
);

INVx2_ASAP7_75t_L g5236 ( 
.A(n_5203),
.Y(n_5236)
);

INVx1_ASAP7_75t_L g5237 ( 
.A(n_5201),
.Y(n_5237)
);

AND2x2_ASAP7_75t_L g5238 ( 
.A(n_5206),
.B(n_5126),
.Y(n_5238)
);

AND2x4_ASAP7_75t_L g5239 ( 
.A(n_5186),
.B(n_5113),
.Y(n_5239)
);

AND2x2_ASAP7_75t_L g5240 ( 
.A(n_5212),
.B(n_5093),
.Y(n_5240)
);

NAND2xp5_ASAP7_75t_L g5241 ( 
.A(n_5179),
.B(n_5104),
.Y(n_5241)
);

INVx2_ASAP7_75t_L g5242 ( 
.A(n_5203),
.Y(n_5242)
);

OR2x2_ASAP7_75t_L g5243 ( 
.A(n_5194),
.B(n_5089),
.Y(n_5243)
);

INVx1_ASAP7_75t_L g5244 ( 
.A(n_5199),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_5199),
.Y(n_5245)
);

BUFx2_ASAP7_75t_L g5246 ( 
.A(n_5165),
.Y(n_5246)
);

INVx2_ASAP7_75t_L g5247 ( 
.A(n_5187),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_5244),
.Y(n_5248)
);

NOR2x1_ASAP7_75t_L g5249 ( 
.A(n_5213),
.B(n_5182),
.Y(n_5249)
);

NAND2xp5_ASAP7_75t_L g5250 ( 
.A(n_5213),
.B(n_5163),
.Y(n_5250)
);

INVx2_ASAP7_75t_L g5251 ( 
.A(n_5217),
.Y(n_5251)
);

AND2x2_ASAP7_75t_L g5252 ( 
.A(n_5217),
.B(n_5142),
.Y(n_5252)
);

OR2x2_ASAP7_75t_L g5253 ( 
.A(n_5214),
.B(n_5194),
.Y(n_5253)
);

NAND2xp5_ASAP7_75t_SL g5254 ( 
.A(n_5228),
.B(n_5197),
.Y(n_5254)
);

INVx1_ASAP7_75t_L g5255 ( 
.A(n_5244),
.Y(n_5255)
);

INVx4_ASAP7_75t_L g5256 ( 
.A(n_5230),
.Y(n_5256)
);

AND2x2_ASAP7_75t_L g5257 ( 
.A(n_5215),
.B(n_5142),
.Y(n_5257)
);

OR2x2_ASAP7_75t_L g5258 ( 
.A(n_5214),
.B(n_5243),
.Y(n_5258)
);

INVx2_ASAP7_75t_L g5259 ( 
.A(n_5221),
.Y(n_5259)
);

INVx1_ASAP7_75t_L g5260 ( 
.A(n_5245),
.Y(n_5260)
);

AND2x2_ASAP7_75t_L g5261 ( 
.A(n_5215),
.B(n_5101),
.Y(n_5261)
);

INVx1_ASAP7_75t_L g5262 ( 
.A(n_5245),
.Y(n_5262)
);

NAND2xp5_ASAP7_75t_L g5263 ( 
.A(n_5235),
.B(n_5210),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_5235),
.Y(n_5264)
);

OR2x2_ASAP7_75t_L g5265 ( 
.A(n_5243),
.B(n_5170),
.Y(n_5265)
);

INVx1_ASAP7_75t_L g5266 ( 
.A(n_5235),
.Y(n_5266)
);

INVx1_ASAP7_75t_L g5267 ( 
.A(n_5235),
.Y(n_5267)
);

NOR2xp33_ASAP7_75t_L g5268 ( 
.A(n_5230),
.B(n_5181),
.Y(n_5268)
);

INVx1_ASAP7_75t_L g5269 ( 
.A(n_5236),
.Y(n_5269)
);

OR2x2_ASAP7_75t_L g5270 ( 
.A(n_5233),
.B(n_5188),
.Y(n_5270)
);

AND2x2_ASAP7_75t_L g5271 ( 
.A(n_5219),
.B(n_5133),
.Y(n_5271)
);

INVx1_ASAP7_75t_L g5272 ( 
.A(n_5236),
.Y(n_5272)
);

AND2x2_ASAP7_75t_L g5273 ( 
.A(n_5219),
.B(n_5105),
.Y(n_5273)
);

OR2x2_ASAP7_75t_L g5274 ( 
.A(n_5251),
.B(n_5218),
.Y(n_5274)
);

OR2x2_ASAP7_75t_L g5275 ( 
.A(n_5251),
.B(n_5218),
.Y(n_5275)
);

NOR2x1p5_ASAP7_75t_SL g5276 ( 
.A(n_5259),
.B(n_5242),
.Y(n_5276)
);

OR2x6_ASAP7_75t_L g5277 ( 
.A(n_5252),
.B(n_5224),
.Y(n_5277)
);

NAND4xp25_ASAP7_75t_L g5278 ( 
.A(n_5250),
.B(n_5226),
.C(n_5241),
.D(n_5246),
.Y(n_5278)
);

OR2x2_ASAP7_75t_L g5279 ( 
.A(n_5258),
.B(n_5229),
.Y(n_5279)
);

OR2x2_ASAP7_75t_L g5280 ( 
.A(n_5270),
.B(n_5229),
.Y(n_5280)
);

OR2x2_ASAP7_75t_L g5281 ( 
.A(n_5253),
.B(n_5246),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_5264),
.Y(n_5282)
);

OR2x2_ASAP7_75t_L g5283 ( 
.A(n_5265),
.B(n_5216),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_5266),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_5267),
.Y(n_5285)
);

OR2x2_ASAP7_75t_L g5286 ( 
.A(n_5259),
.B(n_5216),
.Y(n_5286)
);

OR2x2_ASAP7_75t_L g5287 ( 
.A(n_5263),
.B(n_5207),
.Y(n_5287)
);

NAND2x1p5_ASAP7_75t_L g5288 ( 
.A(n_5256),
.B(n_5230),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_5269),
.Y(n_5289)
);

INVx1_ASAP7_75t_L g5290 ( 
.A(n_5272),
.Y(n_5290)
);

INVx1_ASAP7_75t_L g5291 ( 
.A(n_5263),
.Y(n_5291)
);

AOI22xp5_ASAP7_75t_L g5292 ( 
.A1(n_5278),
.A2(n_5250),
.B1(n_5254),
.B2(n_5249),
.Y(n_5292)
);

INVx1_ASAP7_75t_SL g5293 ( 
.A(n_5283),
.Y(n_5293)
);

NAND2xp5_ASAP7_75t_L g5294 ( 
.A(n_5281),
.B(n_5273),
.Y(n_5294)
);

NAND2xp5_ASAP7_75t_L g5295 ( 
.A(n_5286),
.B(n_5261),
.Y(n_5295)
);

NAND2xp5_ASAP7_75t_L g5296 ( 
.A(n_5274),
.B(n_5234),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_5276),
.Y(n_5297)
);

OAI22xp33_ASAP7_75t_L g5298 ( 
.A1(n_5275),
.A2(n_5189),
.B1(n_5177),
.B2(n_5200),
.Y(n_5298)
);

OR2x2_ASAP7_75t_L g5299 ( 
.A(n_5280),
.B(n_5247),
.Y(n_5299)
);

INVx3_ASAP7_75t_L g5300 ( 
.A(n_5288),
.Y(n_5300)
);

AND2x4_ASAP7_75t_L g5301 ( 
.A(n_5277),
.B(n_5271),
.Y(n_5301)
);

INVx1_ASAP7_75t_L g5302 ( 
.A(n_5279),
.Y(n_5302)
);

OAI21xp5_ASAP7_75t_L g5303 ( 
.A1(n_5287),
.A2(n_5254),
.B(n_5172),
.Y(n_5303)
);

INVx1_ASAP7_75t_L g5304 ( 
.A(n_5299),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_5294),
.Y(n_5305)
);

INVx1_ASAP7_75t_L g5306 ( 
.A(n_5296),
.Y(n_5306)
);

INVx2_ASAP7_75t_L g5307 ( 
.A(n_5301),
.Y(n_5307)
);

INVx1_ASAP7_75t_SL g5308 ( 
.A(n_5293),
.Y(n_5308)
);

AND3x1_ASAP7_75t_L g5309 ( 
.A(n_5292),
.B(n_5268),
.C(n_5190),
.Y(n_5309)
);

AOI22xp33_ASAP7_75t_L g5310 ( 
.A1(n_5303),
.A2(n_5225),
.B1(n_5224),
.B2(n_5238),
.Y(n_5310)
);

NOR2x1_ASAP7_75t_L g5311 ( 
.A(n_5297),
.B(n_5256),
.Y(n_5311)
);

INVx1_ASAP7_75t_L g5312 ( 
.A(n_5295),
.Y(n_5312)
);

NOR2xp33_ASAP7_75t_L g5313 ( 
.A(n_5300),
.B(n_5230),
.Y(n_5313)
);

AND2x2_ASAP7_75t_L g5314 ( 
.A(n_5302),
.B(n_5257),
.Y(n_5314)
);

INVx1_ASAP7_75t_L g5315 ( 
.A(n_5298),
.Y(n_5315)
);

NAND2xp5_ASAP7_75t_L g5316 ( 
.A(n_5301),
.B(n_5221),
.Y(n_5316)
);

NAND2xp5_ASAP7_75t_L g5317 ( 
.A(n_5301),
.B(n_5221),
.Y(n_5317)
);

OAI22xp5_ASAP7_75t_L g5318 ( 
.A1(n_5310),
.A2(n_5190),
.B1(n_5204),
.B2(n_5193),
.Y(n_5318)
);

OAI221xp5_ASAP7_75t_SL g5319 ( 
.A1(n_5309),
.A2(n_5196),
.B1(n_5232),
.B2(n_5209),
.C(n_5238),
.Y(n_5319)
);

INVx2_ASAP7_75t_L g5320 ( 
.A(n_5307),
.Y(n_5320)
);

O2A1O1Ixp33_ASAP7_75t_L g5321 ( 
.A1(n_5315),
.A2(n_5291),
.B(n_5290),
.C(n_5289),
.Y(n_5321)
);

OR2x2_ASAP7_75t_L g5322 ( 
.A(n_5308),
.B(n_5282),
.Y(n_5322)
);

AOI221x1_ASAP7_75t_SL g5323 ( 
.A1(n_5316),
.A2(n_5268),
.B1(n_5285),
.B2(n_5284),
.C(n_5223),
.Y(n_5323)
);

INVx1_ASAP7_75t_L g5324 ( 
.A(n_5314),
.Y(n_5324)
);

AND2x2_ASAP7_75t_L g5325 ( 
.A(n_5313),
.B(n_5222),
.Y(n_5325)
);

OAI22xp33_ASAP7_75t_L g5326 ( 
.A1(n_5317),
.A2(n_5195),
.B1(n_5202),
.B2(n_5234),
.Y(n_5326)
);

NAND4xp25_ASAP7_75t_SL g5327 ( 
.A(n_5305),
.B(n_5209),
.C(n_5222),
.D(n_5232),
.Y(n_5327)
);

INVx1_ASAP7_75t_L g5328 ( 
.A(n_5304),
.Y(n_5328)
);

OAI221xp5_ASAP7_75t_SL g5329 ( 
.A1(n_5326),
.A2(n_5309),
.B1(n_5247),
.B2(n_5312),
.C(n_5306),
.Y(n_5329)
);

NAND2xp5_ASAP7_75t_L g5330 ( 
.A(n_5325),
.B(n_5256),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_5322),
.Y(n_5331)
);

AND2x2_ASAP7_75t_L g5332 ( 
.A(n_5320),
.B(n_5240),
.Y(n_5332)
);

AND2x2_ASAP7_75t_L g5333 ( 
.A(n_5324),
.B(n_5240),
.Y(n_5333)
);

OAI221xp5_ASAP7_75t_L g5334 ( 
.A1(n_5319),
.A2(n_5234),
.B1(n_5311),
.B2(n_5231),
.C(n_5227),
.Y(n_5334)
);

INVx1_ASAP7_75t_L g5335 ( 
.A(n_5328),
.Y(n_5335)
);

NAND2xp5_ASAP7_75t_L g5336 ( 
.A(n_5323),
.B(n_5234),
.Y(n_5336)
);

OAI22xp5_ASAP7_75t_L g5337 ( 
.A1(n_5318),
.A2(n_5205),
.B1(n_5220),
.B2(n_5223),
.Y(n_5337)
);

NAND2xp5_ASAP7_75t_L g5338 ( 
.A(n_5321),
.B(n_5227),
.Y(n_5338)
);

OR2x2_ASAP7_75t_L g5339 ( 
.A(n_5330),
.B(n_5327),
.Y(n_5339)
);

NOR2x1_ASAP7_75t_L g5340 ( 
.A(n_5331),
.B(n_5248),
.Y(n_5340)
);

BUFx2_ASAP7_75t_L g5341 ( 
.A(n_5332),
.Y(n_5341)
);

INVx2_ASAP7_75t_L g5342 ( 
.A(n_5333),
.Y(n_5342)
);

INVx1_ASAP7_75t_L g5343 ( 
.A(n_5338),
.Y(n_5343)
);

INVx2_ASAP7_75t_L g5344 ( 
.A(n_5335),
.Y(n_5344)
);

NAND2xp5_ASAP7_75t_L g5345 ( 
.A(n_5337),
.B(n_5231),
.Y(n_5345)
);

HB1xp67_ASAP7_75t_L g5346 ( 
.A(n_5334),
.Y(n_5346)
);

AOI222xp33_ASAP7_75t_L g5347 ( 
.A1(n_5336),
.A2(n_5237),
.B1(n_5260),
.B2(n_5255),
.C1(n_5262),
.C2(n_5220),
.Y(n_5347)
);

AND2x2_ASAP7_75t_L g5348 ( 
.A(n_5341),
.B(n_5220),
.Y(n_5348)
);

INVx1_ASAP7_75t_L g5349 ( 
.A(n_5345),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_5340),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_5342),
.Y(n_5351)
);

NOR2xp33_ASAP7_75t_L g5352 ( 
.A(n_5339),
.B(n_5329),
.Y(n_5352)
);

NAND4xp25_ASAP7_75t_L g5353 ( 
.A(n_5347),
.B(n_5343),
.C(n_5344),
.D(n_5237),
.Y(n_5353)
);

NOR3xp33_ASAP7_75t_L g5354 ( 
.A(n_5346),
.B(n_5220),
.C(n_5242),
.Y(n_5354)
);

AOI22xp5_ASAP7_75t_L g5355 ( 
.A1(n_5342),
.A2(n_5239),
.B1(n_5158),
.B2(n_5157),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_5341),
.Y(n_5356)
);

NAND3xp33_ASAP7_75t_SL g5357 ( 
.A(n_5341),
.B(n_4845),
.C(n_5160),
.Y(n_5357)
);

AOI22xp5_ASAP7_75t_L g5358 ( 
.A1(n_5342),
.A2(n_5239),
.B1(n_5158),
.B2(n_5157),
.Y(n_5358)
);

NOR3xp33_ASAP7_75t_L g5359 ( 
.A(n_5341),
.B(n_5239),
.C(n_5122),
.Y(n_5359)
);

OAI31xp33_ASAP7_75t_L g5360 ( 
.A1(n_5341),
.A2(n_5239),
.A3(n_5027),
.B(n_5033),
.Y(n_5360)
);

OA22x2_ASAP7_75t_L g5361 ( 
.A1(n_5346),
.A2(n_5122),
.B1(n_5125),
.B2(n_5117),
.Y(n_5361)
);

NOR2x1_ASAP7_75t_L g5362 ( 
.A(n_5340),
.B(n_5056),
.Y(n_5362)
);

NAND2xp5_ASAP7_75t_L g5363 ( 
.A(n_5341),
.B(n_5159),
.Y(n_5363)
);

NAND2xp5_ASAP7_75t_SL g5364 ( 
.A(n_5341),
.B(n_5117),
.Y(n_5364)
);

NAND2xp5_ASAP7_75t_SL g5365 ( 
.A(n_5341),
.B(n_5125),
.Y(n_5365)
);

OAI21xp5_ASAP7_75t_SL g5366 ( 
.A1(n_5348),
.A2(n_5136),
.B(n_5134),
.Y(n_5366)
);

BUFx12f_ASAP7_75t_L g5367 ( 
.A(n_5356),
.Y(n_5367)
);

NAND5xp2_ASAP7_75t_L g5368 ( 
.A(n_5352),
.B(n_5037),
.C(n_5019),
.D(n_5033),
.E(n_5079),
.Y(n_5368)
);

INVx1_ASAP7_75t_L g5369 ( 
.A(n_5362),
.Y(n_5369)
);

NOR2xp33_ASAP7_75t_L g5370 ( 
.A(n_5357),
.B(n_5134),
.Y(n_5370)
);

INVx1_ASAP7_75t_L g5371 ( 
.A(n_5361),
.Y(n_5371)
);

NAND4xp25_ASAP7_75t_L g5372 ( 
.A(n_5354),
.B(n_5079),
.C(n_5136),
.D(n_5059),
.Y(n_5372)
);

AND2x2_ASAP7_75t_L g5373 ( 
.A(n_5360),
.B(n_5121),
.Y(n_5373)
);

NOR3xp33_ASAP7_75t_L g5374 ( 
.A(n_5353),
.B(n_5059),
.C(n_5097),
.Y(n_5374)
);

XNOR2x1_ASAP7_75t_L g5375 ( 
.A(n_5351),
.B(n_5086),
.Y(n_5375)
);

INVx1_ASAP7_75t_L g5376 ( 
.A(n_5359),
.Y(n_5376)
);

NOR2xp33_ASAP7_75t_L g5377 ( 
.A(n_5365),
.B(n_5175),
.Y(n_5377)
);

NAND2xp5_ASAP7_75t_L g5378 ( 
.A(n_5355),
.B(n_5094),
.Y(n_5378)
);

AOI321xp33_ASAP7_75t_L g5379 ( 
.A1(n_5364),
.A2(n_5066),
.A3(n_5106),
.B1(n_5107),
.B2(n_5108),
.C(n_5109),
.Y(n_5379)
);

OAI221xp5_ASAP7_75t_L g5380 ( 
.A1(n_5358),
.A2(n_5175),
.B1(n_5114),
.B2(n_5145),
.C(n_5119),
.Y(n_5380)
);

INVx1_ASAP7_75t_L g5381 ( 
.A(n_5350),
.Y(n_5381)
);

NAND2xp5_ASAP7_75t_SL g5382 ( 
.A(n_5363),
.B(n_5349),
.Y(n_5382)
);

NOR3xp33_ASAP7_75t_L g5383 ( 
.A(n_5356),
.B(n_5081),
.C(n_5085),
.Y(n_5383)
);

NOR3xp33_ASAP7_75t_L g5384 ( 
.A(n_5356),
.B(n_5085),
.C(n_5066),
.Y(n_5384)
);

OAI322xp33_ASAP7_75t_L g5385 ( 
.A1(n_5364),
.A2(n_5120),
.A3(n_5130),
.B1(n_5123),
.B2(n_4982),
.C1(n_4985),
.C2(n_5146),
.Y(n_5385)
);

AOI211xp5_ASAP7_75t_L g5386 ( 
.A1(n_5348),
.A2(n_5118),
.B(n_5132),
.C(n_5112),
.Y(n_5386)
);

NAND2xp5_ASAP7_75t_SL g5387 ( 
.A(n_5348),
.B(n_5112),
.Y(n_5387)
);

NOR3xp33_ASAP7_75t_L g5388 ( 
.A(n_5356),
.B(n_5129),
.C(n_5140),
.Y(n_5388)
);

INVx1_ASAP7_75t_L g5389 ( 
.A(n_5348),
.Y(n_5389)
);

NOR2xp33_ASAP7_75t_L g5390 ( 
.A(n_5348),
.B(n_5052),
.Y(n_5390)
);

NAND2xp33_ASAP7_75t_L g5391 ( 
.A(n_5362),
.B(n_4846),
.Y(n_5391)
);

NOR3xp33_ASAP7_75t_L g5392 ( 
.A(n_5389),
.B(n_5074),
.C(n_5058),
.Y(n_5392)
);

A2O1A1Ixp33_ASAP7_75t_L g5393 ( 
.A1(n_5377),
.A2(n_5012),
.B(n_5058),
.C(n_5031),
.Y(n_5393)
);

AOI221xp5_ASAP7_75t_L g5394 ( 
.A1(n_5366),
.A2(n_5052),
.B1(n_5065),
.B2(n_5047),
.C(n_5023),
.Y(n_5394)
);

NAND2xp5_ASAP7_75t_L g5395 ( 
.A(n_5384),
.B(n_5047),
.Y(n_5395)
);

NAND4xp25_ASAP7_75t_L g5396 ( 
.A(n_5370),
.B(n_5012),
.C(n_5031),
.D(n_339),
.Y(n_5396)
);

NAND4xp25_ASAP7_75t_L g5397 ( 
.A(n_5373),
.B(n_339),
.C(n_336),
.D(n_337),
.Y(n_5397)
);

NOR3xp33_ASAP7_75t_L g5398 ( 
.A(n_5382),
.B(n_336),
.C(n_337),
.Y(n_5398)
);

NAND2xp5_ASAP7_75t_L g5399 ( 
.A(n_5383),
.B(n_5065),
.Y(n_5399)
);

BUFx2_ASAP7_75t_L g5400 ( 
.A(n_5367),
.Y(n_5400)
);

AOI211xp5_ASAP7_75t_L g5401 ( 
.A1(n_5391),
.A2(n_343),
.B(n_340),
.C(n_342),
.Y(n_5401)
);

AND2x2_ASAP7_75t_L g5402 ( 
.A(n_5374),
.B(n_5029),
.Y(n_5402)
);

OAI211xp5_ASAP7_75t_L g5403 ( 
.A1(n_5371),
.A2(n_5084),
.B(n_5060),
.C(n_5029),
.Y(n_5403)
);

AND2x2_ASAP7_75t_L g5404 ( 
.A(n_5388),
.B(n_5075),
.Y(n_5404)
);

OAI221xp5_ASAP7_75t_L g5405 ( 
.A1(n_5381),
.A2(n_5084),
.B1(n_5060),
.B2(n_5023),
.C(n_5016),
.Y(n_5405)
);

NOR2x1_ASAP7_75t_L g5406 ( 
.A(n_5369),
.B(n_5060),
.Y(n_5406)
);

NOR4xp25_ASAP7_75t_L g5407 ( 
.A(n_5376),
.B(n_340),
.C(n_342),
.D(n_343),
.Y(n_5407)
);

NAND3xp33_ASAP7_75t_SL g5408 ( 
.A(n_5390),
.B(n_345),
.C(n_347),
.Y(n_5408)
);

AOI21xp5_ASAP7_75t_L g5409 ( 
.A1(n_5375),
.A2(n_5016),
.B(n_345),
.Y(n_5409)
);

INVx1_ASAP7_75t_L g5410 ( 
.A(n_5387),
.Y(n_5410)
);

OAI221xp5_ASAP7_75t_L g5411 ( 
.A1(n_5379),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.C(n_353),
.Y(n_5411)
);

NOR4xp25_ASAP7_75t_L g5412 ( 
.A(n_5378),
.B(n_348),
.C(n_353),
.D(n_354),
.Y(n_5412)
);

NOR3xp33_ASAP7_75t_L g5413 ( 
.A(n_5372),
.B(n_5380),
.C(n_5386),
.Y(n_5413)
);

NOR2x1p5_ASAP7_75t_L g5414 ( 
.A(n_5368),
.B(n_355),
.Y(n_5414)
);

NAND3xp33_ASAP7_75t_L g5415 ( 
.A(n_5385),
.B(n_355),
.C(n_359),
.Y(n_5415)
);

AND3x2_ASAP7_75t_L g5416 ( 
.A(n_5369),
.B(n_359),
.C(n_360),
.Y(n_5416)
);

NOR2x1_ASAP7_75t_L g5417 ( 
.A(n_5369),
.B(n_361),
.Y(n_5417)
);

OR2x2_ASAP7_75t_L g5418 ( 
.A(n_5372),
.B(n_363),
.Y(n_5418)
);

INVxp67_ASAP7_75t_SL g5419 ( 
.A(n_5389),
.Y(n_5419)
);

OAI211xp5_ASAP7_75t_L g5420 ( 
.A1(n_5371),
.A2(n_363),
.B(n_365),
.C(n_366),
.Y(n_5420)
);

NAND3xp33_ASAP7_75t_L g5421 ( 
.A(n_5401),
.B(n_365),
.C(n_366),
.Y(n_5421)
);

NOR2x1_ASAP7_75t_L g5422 ( 
.A(n_5417),
.B(n_5408),
.Y(n_5422)
);

AOI211xp5_ASAP7_75t_L g5423 ( 
.A1(n_5420),
.A2(n_367),
.B(n_368),
.C(n_369),
.Y(n_5423)
);

NOR4xp25_ASAP7_75t_L g5424 ( 
.A(n_5397),
.B(n_5410),
.C(n_5415),
.D(n_5418),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_5400),
.Y(n_5425)
);

NOR4xp25_ASAP7_75t_L g5426 ( 
.A(n_5411),
.B(n_5419),
.C(n_5396),
.D(n_5399),
.Y(n_5426)
);

NAND2xp33_ASAP7_75t_SL g5427 ( 
.A(n_5414),
.B(n_368),
.Y(n_5427)
);

NAND4xp25_ASAP7_75t_L g5428 ( 
.A(n_5413),
.B(n_369),
.C(n_371),
.D(n_372),
.Y(n_5428)
);

INVx1_ASAP7_75t_L g5429 ( 
.A(n_5416),
.Y(n_5429)
);

NAND3xp33_ASAP7_75t_SL g5430 ( 
.A(n_5412),
.B(n_371),
.C(n_372),
.Y(n_5430)
);

NOR3xp33_ASAP7_75t_SL g5431 ( 
.A(n_5395),
.B(n_373),
.C(n_374),
.Y(n_5431)
);

XNOR2x2_ASAP7_75t_L g5432 ( 
.A(n_5406),
.B(n_374),
.Y(n_5432)
);

OAI21xp5_ASAP7_75t_SL g5433 ( 
.A1(n_5409),
.A2(n_375),
.B(n_376),
.Y(n_5433)
);

OAI221xp5_ASAP7_75t_SL g5434 ( 
.A1(n_5404),
.A2(n_375),
.B1(n_377),
.B2(n_378),
.C(n_379),
.Y(n_5434)
);

AOI211xp5_ASAP7_75t_L g5435 ( 
.A1(n_5407),
.A2(n_377),
.B(n_379),
.C(n_380),
.Y(n_5435)
);

AND2x2_ASAP7_75t_L g5436 ( 
.A(n_5402),
.B(n_380),
.Y(n_5436)
);

NAND4xp25_ASAP7_75t_L g5437 ( 
.A(n_5398),
.B(n_381),
.C(n_382),
.D(n_383),
.Y(n_5437)
);

AND2x2_ASAP7_75t_L g5438 ( 
.A(n_5392),
.B(n_382),
.Y(n_5438)
);

AND2x2_ASAP7_75t_L g5439 ( 
.A(n_5394),
.B(n_383),
.Y(n_5439)
);

NOR4xp25_ASAP7_75t_L g5440 ( 
.A(n_5393),
.B(n_384),
.C(n_385),
.D(n_386),
.Y(n_5440)
);

NOR2xp67_ASAP7_75t_L g5441 ( 
.A(n_5403),
.B(n_387),
.Y(n_5441)
);

AOI221xp5_ASAP7_75t_L g5442 ( 
.A1(n_5405),
.A2(n_387),
.B1(n_389),
.B2(n_392),
.C(n_393),
.Y(n_5442)
);

AND2x2_ASAP7_75t_L g5443 ( 
.A(n_5400),
.B(n_392),
.Y(n_5443)
);

NAND4xp25_ASAP7_75t_L g5444 ( 
.A(n_5413),
.B(n_393),
.C(n_394),
.D(n_395),
.Y(n_5444)
);

INVx1_ASAP7_75t_L g5445 ( 
.A(n_5400),
.Y(n_5445)
);

AOI311xp33_ASAP7_75t_L g5446 ( 
.A1(n_5425),
.A2(n_394),
.A3(n_396),
.B(n_397),
.C(n_399),
.Y(n_5446)
);

CKINVDCx5p33_ASAP7_75t_R g5447 ( 
.A(n_5445),
.Y(n_5447)
);

XNOR2x1_ASAP7_75t_L g5448 ( 
.A(n_5432),
.B(n_399),
.Y(n_5448)
);

INVx1_ASAP7_75t_L g5449 ( 
.A(n_5443),
.Y(n_5449)
);

NOR2xp33_ASAP7_75t_L g5450 ( 
.A(n_5428),
.B(n_400),
.Y(n_5450)
);

NOR3x1_ASAP7_75t_L g5451 ( 
.A(n_5444),
.B(n_400),
.C(n_401),
.Y(n_5451)
);

INVx1_ASAP7_75t_L g5452 ( 
.A(n_5436),
.Y(n_5452)
);

NAND2xp5_ASAP7_75t_L g5453 ( 
.A(n_5435),
.B(n_402),
.Y(n_5453)
);

NOR2xp33_ASAP7_75t_R g5454 ( 
.A(n_5427),
.B(n_404),
.Y(n_5454)
);

AOI21xp5_ASAP7_75t_L g5455 ( 
.A1(n_5422),
.A2(n_406),
.B(n_409),
.Y(n_5455)
);

OAI322xp33_ASAP7_75t_L g5456 ( 
.A1(n_5429),
.A2(n_406),
.A3(n_409),
.B1(n_410),
.B2(n_411),
.C1(n_412),
.C2(n_413),
.Y(n_5456)
);

NAND2xp5_ASAP7_75t_L g5457 ( 
.A(n_5440),
.B(n_411),
.Y(n_5457)
);

OR5x1_ASAP7_75t_L g5458 ( 
.A(n_5430),
.B(n_412),
.C(n_413),
.D(n_414),
.E(n_415),
.Y(n_5458)
);

AND2x2_ASAP7_75t_L g5459 ( 
.A(n_5431),
.B(n_414),
.Y(n_5459)
);

A2O1A1Ixp33_ASAP7_75t_L g5460 ( 
.A1(n_5441),
.A2(n_416),
.B(n_417),
.C(n_418),
.Y(n_5460)
);

AOI221x1_ASAP7_75t_L g5461 ( 
.A1(n_5437),
.A2(n_416),
.B1(n_418),
.B2(n_419),
.C(n_421),
.Y(n_5461)
);

INVx1_ASAP7_75t_SL g5462 ( 
.A(n_5438),
.Y(n_5462)
);

INVxp67_ASAP7_75t_SL g5463 ( 
.A(n_5423),
.Y(n_5463)
);

XOR2x2_ASAP7_75t_L g5464 ( 
.A(n_5448),
.B(n_5421),
.Y(n_5464)
);

AND2x2_ASAP7_75t_L g5465 ( 
.A(n_5459),
.B(n_5424),
.Y(n_5465)
);

NAND4xp75_ASAP7_75t_L g5466 ( 
.A(n_5451),
.B(n_5439),
.C(n_5442),
.D(n_5426),
.Y(n_5466)
);

INVx1_ASAP7_75t_L g5467 ( 
.A(n_5457),
.Y(n_5467)
);

AOI22xp5_ASAP7_75t_L g5468 ( 
.A1(n_5447),
.A2(n_5433),
.B1(n_5434),
.B2(n_422),
.Y(n_5468)
);

NAND3xp33_ASAP7_75t_L g5469 ( 
.A(n_5460),
.B(n_419),
.C(n_421),
.Y(n_5469)
);

NAND2x1p5_ASAP7_75t_L g5470 ( 
.A(n_5452),
.B(n_5449),
.Y(n_5470)
);

XNOR2xp5_ASAP7_75t_L g5471 ( 
.A(n_5458),
.B(n_422),
.Y(n_5471)
);

INVx1_ASAP7_75t_L g5472 ( 
.A(n_5453),
.Y(n_5472)
);

NOR2x1_ASAP7_75t_L g5473 ( 
.A(n_5456),
.B(n_423),
.Y(n_5473)
);

NAND4xp75_ASAP7_75t_L g5474 ( 
.A(n_5461),
.B(n_423),
.C(n_424),
.D(n_425),
.Y(n_5474)
);

NOR2x1_ASAP7_75t_L g5475 ( 
.A(n_5455),
.B(n_425),
.Y(n_5475)
);

INVx1_ASAP7_75t_L g5476 ( 
.A(n_5450),
.Y(n_5476)
);

INVx2_ASAP7_75t_L g5477 ( 
.A(n_5462),
.Y(n_5477)
);

OAI211xp5_ASAP7_75t_L g5478 ( 
.A1(n_5454),
.A2(n_426),
.B(n_427),
.C(n_428),
.Y(n_5478)
);

NAND4xp25_ASAP7_75t_SL g5479 ( 
.A(n_5468),
.B(n_5446),
.C(n_5463),
.D(n_430),
.Y(n_5479)
);

NAND3xp33_ASAP7_75t_SL g5480 ( 
.A(n_5470),
.B(n_427),
.C(n_429),
.Y(n_5480)
);

NOR3xp33_ASAP7_75t_L g5481 ( 
.A(n_5477),
.B(n_429),
.C(n_430),
.Y(n_5481)
);

OR2x2_ASAP7_75t_L g5482 ( 
.A(n_5469),
.B(n_431),
.Y(n_5482)
);

NAND5xp2_ASAP7_75t_L g5483 ( 
.A(n_5465),
.B(n_431),
.C(n_432),
.D(n_433),
.E(n_435),
.Y(n_5483)
);

INVx2_ASAP7_75t_L g5484 ( 
.A(n_5474),
.Y(n_5484)
);

OAI221xp5_ASAP7_75t_L g5485 ( 
.A1(n_5471),
.A2(n_433),
.B1(n_436),
.B2(n_437),
.C(n_438),
.Y(n_5485)
);

AND2x2_ASAP7_75t_L g5486 ( 
.A(n_5473),
.B(n_436),
.Y(n_5486)
);

NOR4xp25_ASAP7_75t_L g5487 ( 
.A(n_5467),
.B(n_437),
.C(n_438),
.D(n_439),
.Y(n_5487)
);

INVx1_ASAP7_75t_L g5488 ( 
.A(n_5478),
.Y(n_5488)
);

NOR3xp33_ASAP7_75t_SL g5489 ( 
.A(n_5466),
.B(n_439),
.C(n_440),
.Y(n_5489)
);

INVx1_ASAP7_75t_L g5490 ( 
.A(n_5475),
.Y(n_5490)
);

NOR4xp25_ASAP7_75t_L g5491 ( 
.A(n_5476),
.B(n_441),
.C(n_442),
.D(n_443),
.Y(n_5491)
);

NAND4xp25_ASAP7_75t_SL g5492 ( 
.A(n_5472),
.B(n_443),
.C(n_444),
.D(n_445),
.Y(n_5492)
);

INVx1_ASAP7_75t_SL g5493 ( 
.A(n_5482),
.Y(n_5493)
);

INVx1_ASAP7_75t_SL g5494 ( 
.A(n_5486),
.Y(n_5494)
);

OR2x2_ASAP7_75t_L g5495 ( 
.A(n_5487),
.B(n_5464),
.Y(n_5495)
);

NAND2xp5_ASAP7_75t_L g5496 ( 
.A(n_5481),
.B(n_444),
.Y(n_5496)
);

INVx1_ASAP7_75t_L g5497 ( 
.A(n_5489),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_5485),
.Y(n_5498)
);

BUFx2_ASAP7_75t_L g5499 ( 
.A(n_5490),
.Y(n_5499)
);

AND2x2_ASAP7_75t_SL g5500 ( 
.A(n_5484),
.B(n_445),
.Y(n_5500)
);

BUFx12f_ASAP7_75t_L g5501 ( 
.A(n_5488),
.Y(n_5501)
);

CKINVDCx20_ASAP7_75t_R g5502 ( 
.A(n_5480),
.Y(n_5502)
);

OAI221xp5_ASAP7_75t_L g5503 ( 
.A1(n_5499),
.A2(n_5491),
.B1(n_5479),
.B2(n_5483),
.C(n_5492),
.Y(n_5503)
);

OAI221xp5_ASAP7_75t_L g5504 ( 
.A1(n_5496),
.A2(n_446),
.B1(n_447),
.B2(n_448),
.C(n_449),
.Y(n_5504)
);

AOI322xp5_ASAP7_75t_L g5505 ( 
.A1(n_5494),
.A2(n_449),
.A3(n_452),
.B1(n_453),
.B2(n_456),
.C1(n_458),
.C2(n_459),
.Y(n_5505)
);

AOI322xp5_ASAP7_75t_L g5506 ( 
.A1(n_5497),
.A2(n_452),
.A3(n_453),
.B1(n_459),
.B2(n_460),
.C1(n_461),
.C2(n_463),
.Y(n_5506)
);

AOI322xp5_ASAP7_75t_L g5507 ( 
.A1(n_5493),
.A2(n_460),
.A3(n_464),
.B1(n_466),
.B2(n_468),
.C1(n_469),
.C2(n_471),
.Y(n_5507)
);

OAI22xp5_ASAP7_75t_L g5508 ( 
.A1(n_5502),
.A2(n_464),
.B1(n_466),
.B2(n_468),
.Y(n_5508)
);

NAND3xp33_ASAP7_75t_SL g5509 ( 
.A(n_5495),
.B(n_471),
.C(n_473),
.Y(n_5509)
);

INVxp67_ASAP7_75t_L g5510 ( 
.A(n_5509),
.Y(n_5510)
);

INVx1_ASAP7_75t_L g5511 ( 
.A(n_5503),
.Y(n_5511)
);

OAI22x1_ASAP7_75t_L g5512 ( 
.A1(n_5504),
.A2(n_5498),
.B1(n_5500),
.B2(n_5501),
.Y(n_5512)
);

NOR3xp33_ASAP7_75t_SL g5513 ( 
.A(n_5511),
.B(n_5508),
.C(n_5505),
.Y(n_5513)
);

OAI22xp33_ASAP7_75t_L g5514 ( 
.A1(n_5510),
.A2(n_5507),
.B1(n_5506),
.B2(n_476),
.Y(n_5514)
);

INVx2_ASAP7_75t_L g5515 ( 
.A(n_5513),
.Y(n_5515)
);

OAI22xp5_ASAP7_75t_L g5516 ( 
.A1(n_5514),
.A2(n_5512),
.B1(n_474),
.B2(n_477),
.Y(n_5516)
);

OAI31xp33_ASAP7_75t_SL g5517 ( 
.A1(n_5516),
.A2(n_473),
.A3(n_478),
.B(n_479),
.Y(n_5517)
);

AOI22xp5_ASAP7_75t_L g5518 ( 
.A1(n_5515),
.A2(n_479),
.B1(n_480),
.B2(n_481),
.Y(n_5518)
);

AOI21xp5_ASAP7_75t_L g5519 ( 
.A1(n_5515),
.A2(n_480),
.B(n_482),
.Y(n_5519)
);

AO22x2_ASAP7_75t_L g5520 ( 
.A1(n_5519),
.A2(n_483),
.B1(n_485),
.B2(n_486),
.Y(n_5520)
);

OAI21x1_ASAP7_75t_L g5521 ( 
.A1(n_5518),
.A2(n_5517),
.B(n_486),
.Y(n_5521)
);

OAI21x1_ASAP7_75t_L g5522 ( 
.A1(n_5519),
.A2(n_483),
.B(n_488),
.Y(n_5522)
);

AOI22xp5_ASAP7_75t_L g5523 ( 
.A1(n_5519),
.A2(n_489),
.B1(n_490),
.B2(n_491),
.Y(n_5523)
);

AOI31xp33_ASAP7_75t_L g5524 ( 
.A1(n_5523),
.A2(n_489),
.A3(n_490),
.B(n_492),
.Y(n_5524)
);

O2A1O1Ixp33_ASAP7_75t_L g5525 ( 
.A1(n_5520),
.A2(n_494),
.B(n_495),
.C(n_497),
.Y(n_5525)
);

AOI21xp5_ASAP7_75t_L g5526 ( 
.A1(n_5521),
.A2(n_495),
.B(n_499),
.Y(n_5526)
);

AOI21xp5_ASAP7_75t_L g5527 ( 
.A1(n_5522),
.A2(n_499),
.B(n_501),
.Y(n_5527)
);

INVx1_ASAP7_75t_L g5528 ( 
.A(n_5522),
.Y(n_5528)
);

AOI22x1_ASAP7_75t_L g5529 ( 
.A1(n_5528),
.A2(n_501),
.B1(n_502),
.B2(n_503),
.Y(n_5529)
);

AOI22xp33_ASAP7_75t_SL g5530 ( 
.A1(n_5526),
.A2(n_5527),
.B1(n_5524),
.B2(n_5525),
.Y(n_5530)
);

AOI22xp5_ASAP7_75t_L g5531 ( 
.A1(n_5526),
.A2(n_504),
.B1(n_505),
.B2(n_506),
.Y(n_5531)
);

OAI21xp5_ASAP7_75t_L g5532 ( 
.A1(n_5526),
.A2(n_506),
.B(n_508),
.Y(n_5532)
);

OAI22xp5_ASAP7_75t_L g5533 ( 
.A1(n_5524),
.A2(n_509),
.B1(n_511),
.B2(n_513),
.Y(n_5533)
);

OAI22xp33_ASAP7_75t_L g5534 ( 
.A1(n_5524),
.A2(n_509),
.B1(n_513),
.B2(n_516),
.Y(n_5534)
);

OA22x2_ASAP7_75t_L g5535 ( 
.A1(n_5528),
.A2(n_517),
.B1(n_518),
.B2(n_519),
.Y(n_5535)
);

OAI22xp33_ASAP7_75t_L g5536 ( 
.A1(n_5524),
.A2(n_517),
.B1(n_519),
.B2(n_520),
.Y(n_5536)
);

AOI22xp5_ASAP7_75t_L g5537 ( 
.A1(n_5526),
.A2(n_521),
.B1(n_522),
.B2(n_523),
.Y(n_5537)
);

OAI22xp33_ASAP7_75t_L g5538 ( 
.A1(n_5524),
.A2(n_523),
.B1(n_524),
.B2(n_525),
.Y(n_5538)
);

OAI22xp33_ASAP7_75t_L g5539 ( 
.A1(n_5524),
.A2(n_526),
.B1(n_527),
.B2(n_530),
.Y(n_5539)
);

AO21x2_ASAP7_75t_L g5540 ( 
.A1(n_5532),
.A2(n_527),
.B(n_530),
.Y(n_5540)
);

NAND3xp33_ASAP7_75t_L g5541 ( 
.A(n_5530),
.B(n_531),
.C(n_532),
.Y(n_5541)
);

OA21x2_ASAP7_75t_L g5542 ( 
.A1(n_5531),
.A2(n_531),
.B(n_532),
.Y(n_5542)
);

AOI21xp5_ASAP7_75t_L g5543 ( 
.A1(n_5534),
.A2(n_1708),
.B(n_1706),
.Y(n_5543)
);

NAND2x1p5_ASAP7_75t_L g5544 ( 
.A(n_5537),
.B(n_1708),
.Y(n_5544)
);

OAI21xp5_ASAP7_75t_L g5545 ( 
.A1(n_5533),
.A2(n_536),
.B(n_537),
.Y(n_5545)
);

OAI22xp5_ASAP7_75t_L g5546 ( 
.A1(n_5536),
.A2(n_536),
.B1(n_537),
.B2(n_538),
.Y(n_5546)
);

OA21x2_ASAP7_75t_L g5547 ( 
.A1(n_5529),
.A2(n_538),
.B(n_539),
.Y(n_5547)
);

INVx1_ASAP7_75t_SL g5548 ( 
.A(n_5540),
.Y(n_5548)
);

AOI22x1_ASAP7_75t_L g5549 ( 
.A1(n_5543),
.A2(n_5539),
.B1(n_5538),
.B2(n_5535),
.Y(n_5549)
);

INVx1_ASAP7_75t_L g5550 ( 
.A(n_5547),
.Y(n_5550)
);

INVx1_ASAP7_75t_L g5551 ( 
.A(n_5544),
.Y(n_5551)
);

INVxp67_ASAP7_75t_L g5552 ( 
.A(n_5542),
.Y(n_5552)
);

AOI221xp5_ASAP7_75t_L g5553 ( 
.A1(n_5552),
.A2(n_5545),
.B1(n_5546),
.B2(n_5541),
.C(n_539),
.Y(n_5553)
);

AOI221xp5_ASAP7_75t_L g5554 ( 
.A1(n_5550),
.A2(n_614),
.B1(n_619),
.B2(n_620),
.C(n_621),
.Y(n_5554)
);

AOI22xp5_ASAP7_75t_L g5555 ( 
.A1(n_5548),
.A2(n_624),
.B1(n_625),
.B2(n_629),
.Y(n_5555)
);

AOI21xp5_ASAP7_75t_L g5556 ( 
.A1(n_5553),
.A2(n_5551),
.B(n_5549),
.Y(n_5556)
);

AOI211xp5_ASAP7_75t_L g5557 ( 
.A1(n_5556),
.A2(n_5554),
.B(n_5555),
.C(n_2230),
.Y(n_5557)
);


endmodule