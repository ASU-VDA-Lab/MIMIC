module fake_jpeg_6588_n_108 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_7),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx5_ASAP7_75t_SL g31 ( 
.A(n_30),
.Y(n_31)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_29),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_20),
.B1(n_14),
.B2(n_17),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_15),
.B1(n_16),
.B2(n_11),
.Y(n_49)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_38),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_46),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_14),
.B1(n_17),
.B2(n_11),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_13),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_40),
.B1(n_48),
.B2(n_33),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_15),
.B1(n_22),
.B2(n_21),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_33),
.B1(n_39),
.B2(n_13),
.Y(n_57)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_21),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_24),
.C(n_39),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_59),
.C(n_63),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_57),
.B1(n_47),
.B2(n_51),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_0),
.Y(n_56)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_24),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_65),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_19),
.C(n_32),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_69),
.B(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_75),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_49),
.C(n_32),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_12),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

OA21x2_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_57),
.B(n_53),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_71),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_19),
.B(n_53),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_80),
.C(n_67),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_72),
.A2(n_32),
.B1(n_19),
.B2(n_21),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_79),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_12),
.B(n_2),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_68),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_90),
.B1(n_79),
.B2(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_73),
.C(n_84),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

AOI221xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_76),
.B1(n_77),
.B2(n_83),
.C(n_82),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_12),
.B1(n_2),
.B2(n_1),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_85),
.C(n_76),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_94),
.Y(n_102)
);

FAx1_ASAP7_75t_SL g101 ( 
.A(n_98),
.B(n_95),
.CI(n_7),
.CON(n_101),
.SN(n_101)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_92),
.B(n_5),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_6),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_101),
.B(n_102),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_97),
.B1(n_96),
.B2(n_1),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_8),
.B(n_9),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

OAI21x1_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_103),
.B(n_102),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_8),
.Y(n_108)
);


endmodule