module fake_jpeg_1288_n_447 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_447);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_447;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_2),
.B(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_17),
.B(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_72),
.Y(n_95)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g138 ( 
.A(n_50),
.Y(n_138)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_0),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_53),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_54),
.B(n_60),
.Y(n_122)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_24),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_1),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_17),
.B(n_15),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_19),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_85),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_21),
.Y(n_85)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_90),
.Y(n_102)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_21),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_92),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_22),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_93),
.B(n_94),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_64),
.A2(n_30),
.B1(n_22),
.B2(n_36),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_104),
.A2(n_106),
.B1(n_108),
.B2(n_113),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_57),
.A2(n_41),
.B1(n_18),
.B2(n_43),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_66),
.A2(n_22),
.B1(n_30),
.B2(n_36),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_51),
.A2(n_18),
.B1(n_27),
.B2(n_43),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_69),
.A2(n_36),
.B1(n_30),
.B2(n_43),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_119),
.A2(n_120),
.B1(n_125),
.B2(n_131),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_63),
.A2(n_42),
.B1(n_39),
.B2(n_27),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_53),
.A2(n_36),
.B1(n_30),
.B2(n_44),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_53),
.A2(n_44),
.B1(n_32),
.B2(n_29),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_60),
.A2(n_32),
.B(n_29),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_68),
.C(n_20),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_65),
.A2(n_27),
.B1(n_42),
.B2(n_39),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_136),
.A2(n_140),
.B1(n_147),
.B2(n_86),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_78),
.A2(n_18),
.B1(n_42),
.B2(n_39),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_60),
.A2(n_38),
.B1(n_45),
.B2(n_33),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_142),
.A2(n_26),
.B1(n_20),
.B2(n_47),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_61),
.A2(n_38),
.B1(n_45),
.B2(n_33),
.Y(n_147)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_150),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_151),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_52),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g225 ( 
.A(n_153),
.B(n_168),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_58),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_156),
.B(n_161),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_97),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_157),
.B(n_165),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_158),
.A2(n_145),
.B1(n_37),
.B2(n_146),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_95),
.B(n_26),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_163),
.Y(n_208)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_111),
.B(n_121),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_122),
.B(n_87),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_77),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_164),
.B(n_173),
.Y(n_219)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_102),
.B(n_49),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_172),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_55),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_169),
.Y(n_235)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_171),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_98),
.B(n_90),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_101),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_13),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_174),
.B(n_175),
.Y(n_237)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

BUFx8_ASAP7_75t_L g203 ( 
.A(n_176),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_97),
.B(n_11),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_177),
.Y(n_217)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_117),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_178),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_139),
.B(n_56),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_185),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_96),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_105),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_183),
.A2(n_187),
.B1(n_192),
.B2(n_195),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g232 ( 
.A1(n_184),
.A2(n_198),
.B1(n_23),
.B2(n_37),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_149),
.B(n_74),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_128),
.B(n_109),
.Y(n_186)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_200),
.Y(n_218)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_99),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_89),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_189),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_113),
.B(n_71),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_112),
.B(n_11),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_190),
.A2(n_193),
.B1(n_141),
.B2(n_135),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_134),
.B(n_12),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_191),
.B(n_196),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_99),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_103),
.B(n_11),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_110),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_106),
.B(n_82),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_4),
.Y(n_236)
);

AO22x1_ASAP7_75t_SL g198 ( 
.A1(n_119),
.A2(n_59),
.B1(n_83),
.B2(n_81),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_104),
.B(n_80),
.C(n_93),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_129),
.C(n_137),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_123),
.B(n_88),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_108),
.B1(n_76),
.B2(n_67),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_202),
.A2(n_228),
.B1(n_196),
.B2(n_195),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_188),
.A2(n_94),
.B1(n_120),
.B2(n_136),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_205),
.A2(n_212),
.B1(n_220),
.B2(n_233),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_236),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_197),
.A2(n_140),
.B1(n_129),
.B2(n_137),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_156),
.B(n_135),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_216),
.B(n_229),
.C(n_230),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_189),
.A2(n_70),
.B1(n_73),
.B2(n_75),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_152),
.A2(n_103),
.B1(n_141),
.B2(n_123),
.Y(n_221)
);

OAI21xp33_ASAP7_75t_SL g278 ( 
.A1(n_221),
.A2(n_226),
.B(n_232),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_154),
.A2(n_145),
.B(n_84),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_222),
.A2(n_4),
.B(n_5),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_223),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_199),
.A2(n_23),
.B1(n_37),
.B2(n_3),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_167),
.B(n_37),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_165),
.B(n_37),
.C(n_23),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_158),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_198),
.A2(n_10),
.B1(n_5),
.B2(n_6),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_241),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_276)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_201),
.B(n_172),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_244),
.B(n_245),
.Y(n_281)
);

A2O1A1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_168),
.B(n_153),
.C(n_186),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_206),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_246),
.B(n_249),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_201),
.B(n_168),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_247),
.B(n_255),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_227),
.A2(n_153),
.B(n_186),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_248),
.A2(n_272),
.B(n_273),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_252),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_200),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_263),
.C(n_213),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_223),
.A2(n_198),
.B1(n_187),
.B2(n_192),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_254),
.A2(n_271),
.B1(n_218),
.B2(n_245),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_160),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_166),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_256),
.B(n_259),
.Y(n_303)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_257),
.Y(n_300)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_258),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_203),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_225),
.Y(n_260)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_260),
.Y(n_306)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_261),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_200),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_170),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_268),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_157),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_265),
.A2(n_209),
.B(n_225),
.Y(n_290)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_266),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_219),
.B(n_150),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_267),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_208),
.B(n_182),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_238),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_270),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_204),
.B(n_180),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_205),
.A2(n_162),
.B1(n_183),
.B2(n_151),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_218),
.A2(n_7),
.B(n_8),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_274),
.A2(n_279),
.B(n_214),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_222),
.B1(n_215),
.B2(n_228),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_231),
.B(n_7),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_237),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_218),
.B(n_10),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_251),
.A2(n_202),
.B1(n_209),
.B2(n_232),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_280),
.B(n_283),
.Y(n_316)
);

AOI22x1_ASAP7_75t_L g282 ( 
.A1(n_275),
.A2(n_212),
.B1(n_241),
.B2(n_220),
.Y(n_282)
);

AO22x1_ASAP7_75t_SL g333 ( 
.A1(n_282),
.A2(n_252),
.B1(n_266),
.B2(n_276),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_250),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_288),
.A2(n_309),
.B1(n_279),
.B2(n_259),
.Y(n_317)
);

NAND2xp33_ASAP7_75t_R g338 ( 
.A(n_290),
.B(n_9),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_296),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_264),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_232),
.B1(n_211),
.B2(n_225),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_297),
.A2(n_298),
.B1(n_307),
.B2(n_312),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_251),
.A2(n_232),
.B1(n_213),
.B2(n_230),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_213),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_304),
.C(n_250),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_249),
.A2(n_207),
.B(n_210),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_302),
.A2(n_274),
.B(n_243),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_262),
.B(n_235),
.C(n_210),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_305),
.B(n_273),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_278),
.A2(n_242),
.B1(n_224),
.B2(n_203),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_244),
.B(n_277),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_8),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_275),
.A2(n_203),
.B1(n_224),
.B2(n_10),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_250),
.A2(n_247),
.B1(n_260),
.B2(n_263),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_313),
.B(n_314),
.C(n_323),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_315),
.A2(n_319),
.B(n_322),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_317),
.A2(n_283),
.B1(n_282),
.B2(n_307),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_291),
.B(n_261),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_318),
.B(n_327),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_288),
.A2(n_279),
.B1(n_248),
.B2(n_246),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_320),
.Y(n_351)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_321),
.Y(n_352)
);

OA21x2_ASAP7_75t_L g322 ( 
.A1(n_281),
.A2(n_265),
.B(n_257),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_299),
.B(n_253),
.C(n_255),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_265),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_324),
.B(n_281),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_325),
.Y(n_341)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_301),
.Y(n_326)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_326),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_295),
.B(n_269),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_291),
.B(n_258),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_332),
.Y(n_344)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_301),
.Y(n_330)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_330),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_303),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_335),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_8),
.C(n_9),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_334),
.B(n_305),
.C(n_306),
.Y(n_363)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_284),
.Y(n_336)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_336),
.Y(n_343)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_284),
.Y(n_337)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_337),
.Y(n_355)
);

XOR2x1_ASAP7_75t_L g349 ( 
.A(n_338),
.B(n_290),
.Y(n_349)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_292),
.Y(n_339)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_339),
.Y(n_360)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_292),
.Y(n_340)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_340),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_342),
.A2(n_316),
.B1(n_331),
.B2(n_322),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_289),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_329),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_348),
.B(n_349),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_316),
.A2(n_331),
.B1(n_280),
.B2(n_286),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_356),
.A2(n_317),
.B(n_293),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_329),
.A2(n_282),
.B1(n_296),
.B2(n_298),
.Y(n_357)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_357),
.Y(n_372)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_330),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_359),
.B(n_363),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_335),
.B(n_294),
.Y(n_361)
);

NOR2x1_ASAP7_75t_L g376 ( 
.A(n_361),
.B(n_294),
.Y(n_376)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_321),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_300),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_313),
.B(n_304),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_347),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_354),
.B(n_314),
.C(n_323),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_366),
.B(n_370),
.C(n_380),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_369),
.A2(n_371),
.B1(n_378),
.B2(n_379),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_324),
.C(n_286),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_375),
.Y(n_394)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_374),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_319),
.Y(n_375)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_376),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_345),
.B(n_322),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_382),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_350),
.A2(n_325),
.B1(n_333),
.B2(n_289),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_345),
.A2(n_303),
.B(n_293),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_306),
.C(n_297),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_341),
.B(n_285),
.C(n_302),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_349),
.C(n_334),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_344),
.B(n_308),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_383),
.B(n_346),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_285),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_384),
.B(n_362),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_341),
.A2(n_340),
.B(n_339),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_385),
.B(n_355),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_387),
.B(n_400),
.Y(n_406)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_388),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_389),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_366),
.B(n_337),
.C(n_361),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_393),
.C(n_396),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_368),
.B(n_351),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g404 ( 
.A(n_391),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_373),
.B(n_359),
.C(n_358),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_372),
.A2(n_350),
.B1(n_333),
.B2(n_360),
.Y(n_395)
);

INVxp33_ASAP7_75t_L g414 ( 
.A(n_395),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_358),
.C(n_364),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_376),
.B(n_343),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_401),
.Y(n_403)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_378),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_402),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_399),
.A2(n_367),
.B(n_371),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_407),
.A2(n_362),
.B(n_360),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_386),
.B(n_380),
.C(n_375),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_408),
.B(n_410),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_386),
.B(n_384),
.C(n_377),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_394),
.B(n_369),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_411),
.B(n_393),
.C(n_412),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_390),
.B(n_381),
.C(n_382),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_412),
.B(n_396),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_425),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_418),
.B(n_419),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_398),
.C(n_394),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_413),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_422),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_404),
.A2(n_392),
.B1(n_397),
.B2(n_395),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_421),
.B(n_423),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_409),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_405),
.B(n_398),
.C(n_400),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_415),
.B(n_387),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_424),
.B(n_406),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_406),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_429),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_420),
.B(n_403),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_430),
.B(n_431),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g431 ( 
.A(n_422),
.B(n_410),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_433),
.B(n_411),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_434),
.B(n_435),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_432),
.B(n_408),
.C(n_414),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_426),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_437),
.A2(n_436),
.B(n_428),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_438),
.A2(n_428),
.B(n_414),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_439),
.A2(n_437),
.B(n_355),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_441),
.B(n_352),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_442),
.B(n_443),
.C(n_343),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_444),
.B(n_440),
.Y(n_445)
);

AOI221xp5_ASAP7_75t_L g446 ( 
.A1(n_445),
.A2(n_353),
.B1(n_326),
.B2(n_300),
.C(n_311),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_446),
.A2(n_309),
.B(n_311),
.Y(n_447)
);


endmodule