module fake_jpeg_30672_n_12 (n_0, n_3, n_2, n_1, n_12);

input n_0;
input n_3;
input n_2;
input n_1;

output n_12;

wire n_11;
wire n_10;
wire n_4;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

INVx1_ASAP7_75t_L g4 ( 
.A(n_3),
.Y(n_4)
);

BUFx5_ASAP7_75t_L g5 ( 
.A(n_0),
.Y(n_5)
);

INVx5_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_SL g7 ( 
.A(n_4),
.B(n_0),
.Y(n_7)
);

AOI22xp5_ASAP7_75t_L g9 ( 
.A1(n_7),
.A2(n_8),
.B1(n_0),
.B2(n_1),
.Y(n_9)
);

O2A1O1Ixp33_ASAP7_75t_L g8 ( 
.A1(n_4),
.A2(n_3),
.B(n_1),
.C(n_2),
.Y(n_8)
);

OAI22xp5_ASAP7_75t_L g10 ( 
.A1(n_9),
.A2(n_6),
.B1(n_5),
.B2(n_2),
.Y(n_10)
);

OAI21xp5_ASAP7_75t_L g11 ( 
.A1(n_10),
.A2(n_9),
.B(n_6),
.Y(n_11)
);

AOI211xp5_ASAP7_75t_L g12 ( 
.A1(n_11),
.A2(n_6),
.B(n_5),
.C(n_2),
.Y(n_12)
);


endmodule