module fake_jpeg_6211_n_245 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_245);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_245;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_34),
.B(n_35),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_13),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_17),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_48),
.Y(n_66)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_37),
.B(n_40),
.Y(n_49)
);

FAx1_ASAP7_75t_SL g70 ( 
.A(n_49),
.B(n_60),
.CI(n_37),
.CON(n_70),
.SN(n_70)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_57),
.B(n_58),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_20),
.B(n_14),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_27),
.B(n_28),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_56),
.B1(n_54),
.B2(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_36),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_79),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_37),
.B1(n_27),
.B2(n_28),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_78),
.B1(n_46),
.B2(n_19),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_14),
.Y(n_90)
);

BUFx24_ASAP7_75t_SL g71 ( 
.A(n_51),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_36),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_76),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_74),
.A2(n_21),
.B(n_15),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_45),
.B1(n_38),
.B2(n_16),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_46),
.B1(n_45),
.B2(n_38),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_36),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_34),
.B1(n_41),
.B2(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_59),
.Y(n_88)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_34),
.B1(n_46),
.B2(n_41),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_92),
.B1(n_94),
.B2(n_78),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_96),
.B(n_72),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_64),
.A2(n_34),
.B1(n_46),
.B2(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_16),
.B1(n_79),
.B2(n_75),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_21),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_98),
.B(n_65),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_103),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_104),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_73),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_113),
.B(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_83),
.B1(n_97),
.B2(n_93),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_86),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_87),
.B(n_76),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_81),
.C(n_74),
.Y(n_123)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_115),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_117),
.B(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_118),
.A2(n_67),
.B1(n_45),
.B2(n_38),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_119),
.A2(n_122),
.B1(n_128),
.B2(n_134),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_89),
.B1(n_68),
.B2(n_90),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_125),
.C(n_131),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_81),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_64),
.B1(n_94),
.B2(n_96),
.Y(n_128)
);

AOI211xp5_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_66),
.B(n_70),
.C(n_77),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_137),
.B1(n_109),
.B2(n_111),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_85),
.C(n_77),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_85),
.C(n_66),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_133),
.C(n_135),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_95),
.C(n_55),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_84),
.B1(n_67),
.B2(n_16),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_67),
.C(n_38),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_140),
.B(n_144),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_121),
.B(n_99),
.Y(n_141)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_102),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_110),
.B1(n_116),
.B2(n_103),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_152),
.B1(n_156),
.B2(n_158),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_155),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_118),
.B1(n_100),
.B2(n_101),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_104),
.Y(n_153)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_101),
.Y(n_154)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_126),
.B1(n_129),
.B2(n_122),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_115),
.B1(n_45),
.B2(n_21),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_127),
.B1(n_19),
.B2(n_21),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_158),
.A2(n_20),
.B(n_18),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_124),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_139),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_42),
.C(n_107),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_42),
.C(n_33),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_156),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_160),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_168),
.C(n_173),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_166),
.A2(n_172),
.B1(n_176),
.B2(n_179),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_127),
.Y(n_168)
);

FAx1_ASAP7_75t_SL g184 ( 
.A(n_169),
.B(n_151),
.CI(n_146),
.CON(n_184),
.SN(n_184)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_42),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_151),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_80),
.B1(n_42),
.B2(n_19),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_42),
.B1(n_19),
.B2(n_20),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_152),
.B1(n_145),
.B2(n_148),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_189),
.B1(n_22),
.B2(n_14),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g181 ( 
.A(n_174),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_195),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_184),
.B(n_187),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_190),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_59),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_188),
.B(n_191),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_176),
.A2(n_82),
.B1(n_22),
.B2(n_18),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_17),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_192),
.A2(n_164),
.B1(n_177),
.B2(n_167),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_82),
.C(n_32),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_194),
.C(n_173),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_17),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_200),
.C(n_201),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_171),
.C(n_172),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_24),
.C(n_15),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_32),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_202),
.B(n_205),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_0),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_32),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_192),
.A2(n_22),
.B1(n_24),
.B2(n_15),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_11),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_185),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_218),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_213),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_224)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_215),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_31),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_217),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_199),
.B(n_1),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_25),
.Y(n_218)
);

OAI21x1_ASAP7_75t_L g219 ( 
.A1(n_218),
.A2(n_198),
.B(n_207),
.Y(n_219)
);

AOI31xp33_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_201),
.A3(n_2),
.B(n_3),
.Y(n_220)
);

NOR2x1_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_226),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_209),
.B(n_1),
.CI(n_4),
.CON(n_225),
.SN(n_225)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_25),
.B(n_30),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_211),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_9),
.C(n_6),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_4),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_26),
.B(n_5),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_231),
.Y(n_235)
);

AOI21x1_ASAP7_75t_L g233 ( 
.A1(n_229),
.A2(n_225),
.B(n_227),
.Y(n_233)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_233),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_232),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_236),
.C(n_237),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_222),
.B(n_5),
.Y(n_236)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

AOI222xp33_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_235),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_242)
);

NAND3xp33_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_243),
.C(n_8),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_4),
.A3(n_6),
.B1(n_8),
.B2(n_9),
.C1(n_241),
.C2(n_219),
.Y(n_243)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_244),
.Y(n_245)
);


endmodule