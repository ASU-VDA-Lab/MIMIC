module fake_ariane_3333_n_1025 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1025);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1025;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_1016;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_462;
wire n_670;
wire n_607;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_731;
wire n_754;
wire n_336;
wire n_665;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_320;
wire n_309;
wire n_559;
wire n_331;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_839;
wire n_928;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_677;
wire n_614;
wire n_604;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_699;
wire n_727;
wire n_590;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_1015;
wire n_644;
wire n_536;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_705;
wire n_630;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_809;
wire n_628;
wire n_461;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_741;
wire n_747;
wire n_772;
wire n_527;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_676;
wire n_708;
wire n_308;
wire n_551;
wire n_417;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_680;
wire n_571;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_755;
wire n_593;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_664;
wire n_629;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_999;
wire n_998;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_751;
wire n_615;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_28),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_148),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_95),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_10),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_197),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_185),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_182),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_133),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_121),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_67),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_172),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_83),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_131),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_154),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_46),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_38),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_106),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_40),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_32),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_108),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_24),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_164),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_85),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_115),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_79),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_36),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_127),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_132),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_184),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_73),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_98),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_196),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_13),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_209),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_9),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_212),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_110),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_28),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_124),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_3),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_64),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_147),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_90),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_213),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_70),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_129),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_168),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_103),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_31),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_43),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_160),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_123),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_136),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_15),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_215),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_114),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_89),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_199),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_175),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_101),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_20),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_179),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_26),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_76),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_25),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_202),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_23),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_18),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_86),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_195),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_87),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_93),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_180),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_25),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_157),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_19),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_211),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_210),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_174),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_99),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_205),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_29),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_116),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_53),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_170),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_176),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_104),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_173),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_155),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_82),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_71),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_137),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_77),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_187),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_111),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_6),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_203),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_78),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_274),
.B(n_0),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_233),
.B(n_0),
.Y(n_321)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_258),
.Y(n_322)
);

BUFx8_ASAP7_75t_SL g323 ( 
.A(n_234),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_258),
.Y(n_324)
);

BUFx8_ASAP7_75t_SL g325 ( 
.A(n_234),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_280),
.B(n_1),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_261),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_258),
.Y(n_328)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_258),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_261),
.Y(n_330)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_319),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_319),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_299),
.B(n_1),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_288),
.B(n_2),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_2),
.Y(n_335)
);

AND2x4_ASAP7_75t_L g336 ( 
.A(n_231),
.B(n_3),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_220),
.B(n_4),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_311),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_228),
.B(n_239),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_319),
.Y(n_340)
);

BUFx8_ASAP7_75t_SL g341 ( 
.A(n_261),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_288),
.B(n_4),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_319),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_231),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_238),
.B(n_5),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_238),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_261),
.Y(n_347)
);

BUFx8_ASAP7_75t_SL g348 ( 
.A(n_289),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_289),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_289),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_223),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_289),
.Y(n_352)
);

BUFx8_ASAP7_75t_SL g353 ( 
.A(n_219),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_241),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_260),
.Y(n_356)
);

AND2x6_ASAP7_75t_L g357 ( 
.A(n_260),
.B(n_33),
.Y(n_357)
);

AND2x4_ASAP7_75t_L g358 ( 
.A(n_270),
.B(n_5),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_305),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_295),
.Y(n_360)
);

INVx5_ASAP7_75t_L g361 ( 
.A(n_285),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_305),
.Y(n_362)
);

AND2x6_ASAP7_75t_L g363 ( 
.A(n_243),
.B(n_34),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_222),
.B(n_6),
.Y(n_364)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_266),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_266),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_240),
.Y(n_367)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_302),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_245),
.B(n_7),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_222),
.B(n_7),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_247),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_248),
.B(n_8),
.Y(n_372)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_302),
.Y(n_373)
);

BUFx12f_ASAP7_75t_L g374 ( 
.A(n_242),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_282),
.B(n_8),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_254),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_351),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_338),
.A2(n_317),
.B1(n_256),
.B2(n_275),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_333),
.A2(n_259),
.B1(n_297),
.B2(n_284),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_L g380 ( 
.A1(n_321),
.A2(n_303),
.B1(n_262),
.B2(n_298),
.Y(n_380)
);

AND2x2_ASAP7_75t_SL g381 ( 
.A(n_364),
.B(n_249),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_354),
.Y(n_382)
);

OR2x6_ASAP7_75t_L g383 ( 
.A(n_374),
.B(n_265),
.Y(n_383)
);

OAI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_321),
.A2(n_314),
.B1(n_306),
.B2(n_271),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_327),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_349),
.Y(n_386)
);

AO22x2_ASAP7_75t_L g387 ( 
.A1(n_326),
.A2(n_269),
.B1(n_272),
.B2(n_279),
.Y(n_387)
);

OA22x2_ASAP7_75t_L g388 ( 
.A1(n_360),
.A2(n_281),
.B1(n_293),
.B2(n_296),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_370),
.A2(n_300),
.B1(n_304),
.B2(n_313),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_366),
.B(n_221),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_326),
.A2(n_316),
.B1(n_315),
.B2(n_312),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_366),
.B(n_224),
.Y(n_392)
);

OAI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_320),
.A2(n_310),
.B1(n_309),
.B2(n_308),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_344),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_365),
.B(n_225),
.Y(n_395)
);

OAI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_333),
.A2(n_335),
.B1(n_366),
.B2(n_358),
.Y(n_396)
);

NAND2xp33_ASAP7_75t_SL g397 ( 
.A(n_334),
.B(n_226),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_227),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_229),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_344),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_335),
.A2(n_307),
.B1(n_301),
.B2(n_294),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_375),
.A2(n_292),
.B1(n_291),
.B2(n_290),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_344),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_365),
.B(n_230),
.Y(n_404)
);

AO22x2_ASAP7_75t_L g405 ( 
.A1(n_342),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_367),
.A2(n_287),
.B1(n_283),
.B2(n_278),
.Y(n_406)
);

AO22x2_ASAP7_75t_L g407 ( 
.A1(n_336),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_232),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_368),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_356),
.Y(n_410)
);

OAI22xp33_ASAP7_75t_L g411 ( 
.A1(n_374),
.A2(n_277),
.B1(n_276),
.B2(n_273),
.Y(n_411)
);

AO22x2_ASAP7_75t_L g412 ( 
.A1(n_336),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_412)
);

OA22x2_ASAP7_75t_L g413 ( 
.A1(n_376),
.A2(n_268),
.B1(n_267),
.B2(n_264),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_336),
.A2(n_263),
.B1(n_257),
.B2(n_255),
.Y(n_414)
);

OA22x2_ASAP7_75t_L g415 ( 
.A1(n_358),
.A2(n_253),
.B1(n_252),
.B2(n_251),
.Y(n_415)
);

OAI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_358),
.A2(n_339),
.B1(n_372),
.B2(n_337),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_327),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_327),
.Y(n_418)
);

OAI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_345),
.A2(n_250),
.B1(n_246),
.B2(n_244),
.Y(n_419)
);

OR2x6_ASAP7_75t_L g420 ( 
.A(n_353),
.B(n_355),
.Y(n_420)
);

OAI22xp33_ASAP7_75t_L g421 ( 
.A1(n_368),
.A2(n_237),
.B1(n_236),
.B2(n_235),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_345),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_368),
.B(n_16),
.Y(n_423)
);

AO22x2_ASAP7_75t_L g424 ( 
.A1(n_345),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_356),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_373),
.B(n_20),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_347),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_373),
.B(n_21),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_373),
.B(n_21),
.Y(n_429)
);

OAI22xp33_ASAP7_75t_SL g430 ( 
.A1(n_373),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_361),
.B(n_35),
.Y(n_431)
);

OAI22xp33_ASAP7_75t_SL g432 ( 
.A1(n_369),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_432)
);

BUFx10_ASAP7_75t_L g433 ( 
.A(n_344),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_353),
.Y(n_434)
);

OAI22xp33_ASAP7_75t_L g435 ( 
.A1(n_355),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_381),
.B(n_371),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_403),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_377),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_434),
.B(n_323),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_382),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_378),
.B(n_323),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_385),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_416),
.A2(n_363),
.B(n_357),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_417),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_418),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_379),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_401),
.B(n_325),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_410),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_410),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_406),
.B(n_413),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_425),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_425),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_390),
.A2(n_363),
.B(n_357),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_403),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_392),
.B(n_371),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_394),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_400),
.Y(n_458)
);

INVxp33_ASAP7_75t_L g459 ( 
.A(n_387),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_433),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_433),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_386),
.Y(n_462)
);

XNOR2x2_ASAP7_75t_L g463 ( 
.A(n_405),
.B(n_325),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_388),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_393),
.B(n_346),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_423),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_420),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_426),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_SL g469 ( 
.A(n_428),
.B(n_346),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_429),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_386),
.Y(n_471)
);

AND2x2_ASAP7_75t_SL g472 ( 
.A(n_422),
.B(n_369),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_399),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_420),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_386),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_391),
.B(n_341),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

CKINVDCx14_ASAP7_75t_R g478 ( 
.A(n_383),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_398),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_383),
.B(n_346),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_404),
.B(n_346),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_R g482 ( 
.A(n_396),
.B(n_330),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_415),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_409),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_395),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_389),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_397),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_408),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_414),
.B(n_402),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_384),
.A2(n_380),
.B(n_419),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_407),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_421),
.B(n_361),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_407),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_412),
.Y(n_494)
);

AND2x6_ASAP7_75t_L g495 ( 
.A(n_431),
.B(n_363),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_412),
.B(n_356),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_424),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_424),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_411),
.B(n_361),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_405),
.B(n_356),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_432),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_435),
.B(n_359),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_430),
.B(n_341),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_377),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_377),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_416),
.B(n_361),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_390),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_403),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_377),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_377),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_377),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_377),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_462),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_449),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_450),
.Y(n_515)
);

NOR2xp67_ASAP7_75t_L g516 ( 
.A(n_473),
.B(n_361),
.Y(n_516)
);

INVxp33_ASAP7_75t_L g517 ( 
.A(n_439),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_R g518 ( 
.A(n_478),
.B(n_467),
.Y(n_518)
);

AND2x6_ASAP7_75t_L g519 ( 
.A(n_496),
.B(n_363),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_436),
.B(n_359),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_452),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_456),
.B(n_359),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_480),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_453),
.Y(n_524)
);

BUFx12f_ASAP7_75t_SL g525 ( 
.A(n_489),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_481),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_R g527 ( 
.A(n_478),
.B(n_363),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_454),
.A2(n_357),
.B(n_330),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_443),
.A2(n_473),
.B(n_488),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_442),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_486),
.B(n_348),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_444),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_462),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_456),
.B(n_359),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_437),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_507),
.B(n_466),
.Y(n_536)
);

INVxp67_ASAP7_75t_SL g537 ( 
.A(n_461),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_502),
.B(n_362),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_468),
.B(n_362),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_470),
.B(n_362),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_498),
.B(n_362),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_479),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_482),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_445),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_501),
.B(n_347),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_491),
.B(n_494),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_438),
.B(n_322),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_497),
.B(n_347),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_440),
.B(n_504),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_464),
.B(n_350),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_477),
.B(n_357),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_472),
.B(n_350),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_482),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_448),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_457),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_508),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_460),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_471),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_495),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_472),
.B(n_350),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_500),
.Y(n_561)
);

AND2x2_ASAP7_75t_SL g562 ( 
.A(n_503),
.B(n_357),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_505),
.B(n_322),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_459),
.B(n_322),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_459),
.B(n_509),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_495),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_510),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_499),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_458),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_511),
.B(n_329),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_455),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_512),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_475),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_469),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_499),
.B(n_329),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_506),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_490),
.B(n_329),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_485),
.B(n_30),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_465),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_487),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_490),
.B(n_332),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_487),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_506),
.B(n_332),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_493),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_483),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_495),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_484),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_451),
.B(n_332),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_495),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_492),
.B(n_349),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_495),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_492),
.B(n_348),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_469),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_493),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_474),
.B(n_349),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_446),
.A2(n_352),
.B1(n_349),
.B2(n_343),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_446),
.B(n_31),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_467),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_447),
.B(n_352),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_463),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_580),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_573),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_514),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_529),
.B(n_352),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_526),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_526),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_538),
.B(n_352),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_580),
.Y(n_608)
);

BUFx12f_ASAP7_75t_L g609 ( 
.A(n_582),
.Y(n_609)
);

OR2x6_ASAP7_75t_L g610 ( 
.A(n_582),
.B(n_476),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_572),
.Y(n_611)
);

BUFx4f_ASAP7_75t_L g612 ( 
.A(n_595),
.Y(n_612)
);

BUFx2_ASAP7_75t_SL g613 ( 
.A(n_595),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_572),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_546),
.B(n_32),
.Y(n_615)
);

BUFx12f_ASAP7_75t_L g616 ( 
.A(n_542),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_514),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_588),
.B(n_441),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_541),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_573),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_538),
.B(n_576),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_521),
.Y(n_622)
);

NAND2x1_ASAP7_75t_SL g623 ( 
.A(n_531),
.B(n_37),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_541),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_SL g625 ( 
.A(n_559),
.B(n_566),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_588),
.B(n_523),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_518),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_SL g628 ( 
.A(n_559),
.B(n_331),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_568),
.B(n_331),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_586),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_586),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_573),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_586),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_521),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_576),
.B(n_324),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_520),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_543),
.B(n_331),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_515),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_553),
.B(n_331),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_520),
.B(n_324),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_546),
.B(n_39),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_564),
.B(n_324),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_565),
.B(n_41),
.Y(n_643)
);

INVx6_ASAP7_75t_L g644 ( 
.A(n_526),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_L g645 ( 
.A(n_586),
.B(n_324),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_573),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_524),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_552),
.B(n_328),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_523),
.B(n_331),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_552),
.B(n_328),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_560),
.B(n_598),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_524),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_525),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_565),
.B(n_42),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_560),
.B(n_542),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_586),
.Y(n_656)
);

NOR2x1p5_ASAP7_75t_L g657 ( 
.A(n_537),
.B(n_343),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_589),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_515),
.Y(n_659)
);

BUFx12f_ASAP7_75t_L g660 ( 
.A(n_599),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_550),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_550),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_525),
.B(n_328),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_585),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_564),
.B(n_328),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_574),
.Y(n_666)
);

OR2x6_ASAP7_75t_L g667 ( 
.A(n_578),
.B(n_340),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_609),
.B(n_578),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_626),
.B(n_597),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_601),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_644),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_611),
.Y(n_672)
);

INVx3_ASAP7_75t_SL g673 ( 
.A(n_627),
.Y(n_673)
);

INVx5_ASAP7_75t_L g674 ( 
.A(n_644),
.Y(n_674)
);

BUFx5_ASAP7_75t_L g675 ( 
.A(n_641),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_602),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_603),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_616),
.Y(n_678)
);

OR2x6_ASAP7_75t_L g679 ( 
.A(n_613),
.B(n_578),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_608),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_666),
.B(n_557),
.Y(n_681)
);

INVxp67_ASAP7_75t_SL g682 ( 
.A(n_641),
.Y(n_682)
);

CKINVDCx16_ASAP7_75t_R g683 ( 
.A(n_610),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_653),
.Y(n_684)
);

CKINVDCx11_ASAP7_75t_R g685 ( 
.A(n_610),
.Y(n_685)
);

BUFx4_ASAP7_75t_SL g686 ( 
.A(n_610),
.Y(n_686)
);

BUFx12f_ASAP7_75t_L g687 ( 
.A(n_660),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_651),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_614),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_666),
.B(n_567),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_612),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_612),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_615),
.Y(n_693)
);

BUFx12f_ASAP7_75t_L g694 ( 
.A(n_615),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_644),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_643),
.Y(n_696)
);

INVxp33_ASAP7_75t_L g697 ( 
.A(n_655),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_655),
.B(n_567),
.Y(n_698)
);

BUFx12f_ASAP7_75t_L g699 ( 
.A(n_643),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_664),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_638),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_602),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_659),
.Y(n_703)
);

CKINVDCx14_ASAP7_75t_R g704 ( 
.A(n_618),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_650),
.Y(n_705)
);

INVx3_ASAP7_75t_SL g706 ( 
.A(n_654),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_654),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_636),
.A2(n_574),
.B1(n_578),
.B2(n_562),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_617),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_636),
.B(n_522),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_622),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_634),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_658),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_602),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_620),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_620),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_648),
.Y(n_717)
);

INVxp67_ASAP7_75t_SL g718 ( 
.A(n_658),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_661),
.B(n_599),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_619),
.B(n_522),
.Y(n_720)
);

BUFx12f_ASAP7_75t_L g721 ( 
.A(n_667),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_663),
.Y(n_722)
);

BUFx12f_ASAP7_75t_L g723 ( 
.A(n_685),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_677),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_672),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_669),
.B(n_600),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_691),
.Y(n_727)
);

INVx5_ASAP7_75t_L g728 ( 
.A(n_699),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_682),
.A2(n_681),
.B1(n_696),
.B2(n_690),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_689),
.Y(n_730)
);

BUFx8_ASAP7_75t_L g731 ( 
.A(n_687),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_677),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_701),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_687),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_686),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_704),
.A2(n_600),
.B1(n_579),
.B2(n_562),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_704),
.A2(n_562),
.B1(n_561),
.B2(n_584),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_703),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_706),
.A2(n_667),
.B1(n_549),
.B2(n_606),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_685),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_699),
.A2(n_584),
.B1(n_594),
.B2(n_647),
.Y(n_741)
);

INVx1_ASAP7_75t_SL g742 ( 
.A(n_670),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_719),
.A2(n_594),
.B1(n_652),
.B2(n_569),
.Y(n_743)
);

BUFx4f_ASAP7_75t_SL g744 ( 
.A(n_673),
.Y(n_744)
);

BUFx10_ASAP7_75t_L g745 ( 
.A(n_678),
.Y(n_745)
);

CKINVDCx11_ASAP7_75t_R g746 ( 
.A(n_673),
.Y(n_746)
);

OAI22x1_ASAP7_75t_L g747 ( 
.A1(n_706),
.A2(n_596),
.B1(n_592),
.B2(n_663),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_700),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_707),
.A2(n_667),
.B1(n_605),
.B2(n_606),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_709),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_691),
.Y(n_751)
);

BUFx8_ASAP7_75t_SL g752 ( 
.A(n_684),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_684),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_709),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_688),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_693),
.B(n_548),
.Y(n_756)
);

BUFx4f_ASAP7_75t_SL g757 ( 
.A(n_694),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_711),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_718),
.A2(n_625),
.B(n_604),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_674),
.Y(n_760)
);

NAND2x1p5_ASAP7_75t_L g761 ( 
.A(n_674),
.B(n_605),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_SL g762 ( 
.A1(n_679),
.A2(n_566),
.B(n_559),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_711),
.Y(n_763)
);

INVx6_ASAP7_75t_L g764 ( 
.A(n_674),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_694),
.B(n_548),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_712),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_681),
.A2(n_624),
.B1(n_629),
.B2(n_536),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_690),
.A2(n_629),
.B1(n_662),
.B2(n_519),
.Y(n_768)
);

BUFx12f_ASAP7_75t_L g769 ( 
.A(n_668),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_712),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_697),
.A2(n_569),
.B1(n_555),
.B2(n_532),
.Y(n_771)
);

CKINVDCx11_ASAP7_75t_R g772 ( 
.A(n_683),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_725),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_726),
.A2(n_675),
.B1(n_668),
.B2(n_679),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_729),
.A2(n_697),
.B1(n_698),
.B2(n_708),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_736),
.A2(n_675),
.B1(n_668),
.B2(n_679),
.Y(n_776)
);

INVx1_ASAP7_75t_SL g777 ( 
.A(n_742),
.Y(n_777)
);

OAI222xp33_ASAP7_75t_L g778 ( 
.A1(n_737),
.A2(n_596),
.B1(n_717),
.B2(n_722),
.C1(n_705),
.C2(n_710),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_755),
.B(n_680),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_748),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_730),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_741),
.A2(n_675),
.B1(n_532),
.B2(n_517),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_SL g783 ( 
.A1(n_767),
.A2(n_623),
.B(n_593),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_752),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_760),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_760),
.Y(n_786)
);

AOI222xp33_ASAP7_75t_L g787 ( 
.A1(n_756),
.A2(n_585),
.B1(n_545),
.B2(n_720),
.C1(n_544),
.C2(n_554),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_747),
.A2(n_675),
.B1(n_555),
.B2(n_649),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_735),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_733),
.Y(n_790)
);

BUFx12f_ASAP7_75t_L g791 ( 
.A(n_731),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_738),
.Y(n_792)
);

OAI21xp33_ASAP7_75t_L g793 ( 
.A1(n_771),
.A2(n_587),
.B(n_540),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_746),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_750),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_743),
.A2(n_675),
.B1(n_554),
.B2(n_530),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_753),
.B(n_695),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_SL g798 ( 
.A1(n_739),
.A2(n_675),
.B1(n_721),
.B2(n_519),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_755),
.A2(n_544),
.B1(n_530),
.B2(n_657),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_764),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_739),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_765),
.A2(n_771),
.B1(n_758),
.B2(n_763),
.Y(n_802)
);

CKINVDCx6p67_ASAP7_75t_R g803 ( 
.A(n_723),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_754),
.A2(n_692),
.B1(n_721),
.B2(n_587),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_744),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_SL g806 ( 
.A1(n_728),
.A2(n_519),
.B1(n_692),
.B2(n_621),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_766),
.A2(n_621),
.B1(n_534),
.B2(n_519),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_SL g808 ( 
.A1(n_768),
.A2(n_593),
.B(n_575),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_724),
.A2(n_770),
.B1(n_732),
.B2(n_769),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_727),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_749),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_749),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_742),
.A2(n_674),
.B1(n_695),
.B2(n_671),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_744),
.A2(n_671),
.B1(n_516),
.B2(n_713),
.Y(n_814)
);

BUFx4f_ASAP7_75t_SL g815 ( 
.A(n_731),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_772),
.A2(n_534),
.B1(n_519),
.B2(n_639),
.Y(n_816)
);

NAND3xp33_ASAP7_75t_L g817 ( 
.A(n_728),
.B(n_581),
.C(n_577),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_727),
.Y(n_818)
);

AOI222xp33_ASAP7_75t_L g819 ( 
.A1(n_757),
.A2(n_545),
.B1(n_519),
.B2(n_539),
.C1(n_571),
.C2(n_665),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_740),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_SL g821 ( 
.A1(n_728),
.A2(n_519),
.B1(n_527),
.B2(n_528),
.Y(n_821)
);

OAI21xp33_ASAP7_75t_L g822 ( 
.A1(n_734),
.A2(n_563),
.B(n_547),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_727),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_757),
.A2(n_637),
.B1(n_639),
.B2(n_590),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_751),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_751),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_728),
.A2(n_637),
.B1(n_590),
.B2(n_571),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_761),
.A2(n_671),
.B1(n_516),
.B2(n_713),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_782),
.A2(n_751),
.B1(n_573),
.B2(n_642),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_780),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_800),
.B(n_676),
.Y(n_831)
);

OAI22xp33_ASAP7_75t_L g832 ( 
.A1(n_783),
.A2(n_764),
.B1(n_761),
.B2(n_713),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_824),
.A2(n_764),
.B1(n_702),
.B2(n_715),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_775),
.A2(n_665),
.B1(n_642),
.B2(n_535),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_777),
.B(n_702),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_779),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_780),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_781),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_787),
.A2(n_556),
.B1(n_535),
.B2(n_583),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_781),
.B(n_715),
.Y(n_840)
);

OA21x2_ASAP7_75t_L g841 ( 
.A1(n_788),
.A2(n_759),
.B(n_635),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_809),
.A2(n_556),
.B1(n_535),
.B2(n_607),
.Y(n_842)
);

OAI21xp33_ASAP7_75t_SL g843 ( 
.A1(n_801),
.A2(n_786),
.B(n_785),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_773),
.B(n_716),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_801),
.A2(n_716),
.B1(n_759),
.B2(n_676),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_790),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_816),
.A2(n_714),
.B1(n_676),
.B2(n_620),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_792),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_SL g849 ( 
.A1(n_811),
.A2(n_528),
.B1(n_551),
.B2(n_632),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_819),
.A2(n_556),
.B1(n_607),
.B2(n_558),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_812),
.B(n_676),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_795),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_SL g853 ( 
.A1(n_817),
.A2(n_551),
.B1(n_646),
.B2(n_632),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_802),
.A2(n_558),
.B1(n_640),
.B2(n_646),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_SL g855 ( 
.A1(n_778),
.A2(n_551),
.B1(n_646),
.B2(n_632),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_776),
.A2(n_714),
.B1(n_558),
.B2(n_762),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_798),
.A2(n_640),
.B1(n_551),
.B2(n_513),
.Y(n_857)
);

OA21x2_ASAP7_75t_L g858 ( 
.A1(n_808),
.A2(n_635),
.B(n_570),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_810),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_SL g860 ( 
.A(n_791),
.B(n_745),
.Y(n_860)
);

NAND4xp25_ASAP7_75t_SL g861 ( 
.A(n_784),
.B(n_745),
.C(n_45),
.D(n_47),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_797),
.B(n_818),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_796),
.A2(n_714),
.B1(n_656),
.B2(n_630),
.Y(n_863)
);

AOI222xp33_ASAP7_75t_L g864 ( 
.A1(n_774),
.A2(n_513),
.B1(n_533),
.B2(n_645),
.C1(n_714),
.C2(n_340),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_823),
.B(n_825),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_798),
.A2(n_513),
.B1(n_533),
.B2(n_656),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_826),
.Y(n_867)
);

OAI22xp33_ASAP7_75t_L g868 ( 
.A1(n_815),
.A2(n_625),
.B1(n_631),
.B2(n_630),
.Y(n_868)
);

NAND3xp33_ASAP7_75t_L g869 ( 
.A(n_822),
.B(n_533),
.C(n_340),
.Y(n_869)
);

OAI22xp33_ASAP7_75t_L g870 ( 
.A1(n_803),
.A2(n_633),
.B1(n_631),
.B2(n_566),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_793),
.A2(n_633),
.B1(n_591),
.B2(n_589),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_SL g872 ( 
.A1(n_813),
.A2(n_800),
.B1(n_814),
.B2(n_828),
.Y(n_872)
);

AOI222xp33_ASAP7_75t_L g873 ( 
.A1(n_804),
.A2(n_799),
.B1(n_827),
.B2(n_807),
.C1(n_800),
.C2(n_805),
.Y(n_873)
);

OAI221xp5_ASAP7_75t_SL g874 ( 
.A1(n_832),
.A2(n_806),
.B1(n_821),
.B2(n_785),
.C(n_786),
.Y(n_874)
);

OAI21xp33_ASAP7_75t_L g875 ( 
.A1(n_843),
.A2(n_794),
.B(n_806),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_855),
.A2(n_821),
.B1(n_820),
.B2(n_789),
.Y(n_876)
);

NAND3xp33_ASAP7_75t_L g877 ( 
.A(n_872),
.B(n_800),
.C(n_343),
.Y(n_877)
);

NAND3xp33_ASAP7_75t_L g878 ( 
.A(n_872),
.B(n_343),
.C(n_340),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_SL g879 ( 
.A1(n_861),
.A2(n_591),
.B(n_48),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_862),
.B(n_44),
.Y(n_880)
);

AOI221xp5_ASAP7_75t_L g881 ( 
.A1(n_836),
.A2(n_846),
.B1(n_852),
.B2(n_838),
.C(n_830),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_837),
.B(n_49),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_855),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_848),
.B(n_54),
.Y(n_884)
);

NAND3xp33_ASAP7_75t_L g885 ( 
.A(n_867),
.B(n_628),
.C(n_56),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_SL g886 ( 
.A1(n_873),
.A2(n_55),
.B(n_57),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_840),
.B(n_58),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_854),
.A2(n_628),
.B1(n_60),
.B2(n_61),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_835),
.B(n_844),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_851),
.B(n_59),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_865),
.B(n_62),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_859),
.B(n_218),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_SL g893 ( 
.A(n_860),
.B(n_63),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_845),
.B(n_217),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_834),
.A2(n_839),
.B1(n_849),
.B2(n_869),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_858),
.B(n_65),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_866),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_897)
);

OAI21xp33_ASAP7_75t_L g898 ( 
.A1(n_853),
.A2(n_72),
.B(n_74),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_858),
.B(n_75),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_831),
.B(n_216),
.Y(n_900)
);

NOR3xp33_ASAP7_75t_SL g901 ( 
.A(n_868),
.B(n_80),
.C(n_81),
.Y(n_901)
);

NAND3xp33_ASAP7_75t_L g902 ( 
.A(n_853),
.B(n_84),
.C(n_88),
.Y(n_902)
);

AOI21xp33_ASAP7_75t_L g903 ( 
.A1(n_856),
.A2(n_91),
.B(n_92),
.Y(n_903)
);

OAI221xp5_ASAP7_75t_L g904 ( 
.A1(n_833),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.C(n_100),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_868),
.B(n_102),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_849),
.B(n_214),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_881),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_889),
.B(n_841),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_886),
.A2(n_847),
.B1(n_870),
.B2(n_863),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_899),
.B(n_841),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_896),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_890),
.B(n_870),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_896),
.B(n_857),
.Y(n_913)
);

NAND3xp33_ASAP7_75t_L g914 ( 
.A(n_882),
.B(n_850),
.C(n_842),
.Y(n_914)
);

INVxp67_ASAP7_75t_SL g915 ( 
.A(n_882),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_875),
.B(n_829),
.Y(n_916)
);

OR2x2_ASAP7_75t_L g917 ( 
.A(n_874),
.B(n_871),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_890),
.B(n_880),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_887),
.B(n_105),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_884),
.Y(n_920)
);

NAND4xp75_ASAP7_75t_L g921 ( 
.A(n_901),
.B(n_864),
.C(n_109),
.D(n_112),
.Y(n_921)
);

NAND3xp33_ASAP7_75t_SL g922 ( 
.A(n_879),
.B(n_107),
.C(n_113),
.Y(n_922)
);

AO21x2_ASAP7_75t_L g923 ( 
.A1(n_892),
.A2(n_117),
.B(n_118),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_884),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_876),
.B(n_119),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_905),
.B(n_120),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_908),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_918),
.B(n_893),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_915),
.B(n_895),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_907),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_911),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_911),
.B(n_906),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_924),
.Y(n_933)
);

XNOR2xp5_ASAP7_75t_L g934 ( 
.A(n_918),
.B(n_877),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_910),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_920),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_910),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_920),
.B(n_894),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_913),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_913),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_912),
.B(n_895),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_928),
.Y(n_942)
);

XNOR2xp5_ASAP7_75t_L g943 ( 
.A(n_934),
.B(n_925),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_941),
.A2(n_916),
.B1(n_925),
.B2(n_922),
.Y(n_944)
);

XOR2x2_ASAP7_75t_L g945 ( 
.A(n_929),
.B(n_930),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_939),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_937),
.Y(n_947)
);

XNOR2x1_ASAP7_75t_L g948 ( 
.A(n_940),
.B(n_917),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_937),
.Y(n_949)
);

OA22x2_ASAP7_75t_L g950 ( 
.A1(n_943),
.A2(n_940),
.B1(n_927),
.B2(n_935),
.Y(n_950)
);

AOI22x1_ASAP7_75t_SL g951 ( 
.A1(n_945),
.A2(n_933),
.B1(n_935),
.B2(n_936),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_946),
.Y(n_952)
);

XOR2x2_ASAP7_75t_L g953 ( 
.A(n_948),
.B(n_914),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_944),
.A2(n_909),
.B1(n_917),
.B2(n_932),
.Y(n_954)
);

AOI22x1_ASAP7_75t_L g955 ( 
.A1(n_947),
.A2(n_938),
.B1(n_926),
.B2(n_916),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_942),
.A2(n_938),
.B1(n_921),
.B2(n_926),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_947),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_952),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_957),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_954),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_955),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_950),
.Y(n_962)
);

NAND4xp75_ASAP7_75t_L g963 ( 
.A(n_962),
.B(n_951),
.C(n_956),
.D(n_953),
.Y(n_963)
);

NAND4xp75_ASAP7_75t_L g964 ( 
.A(n_961),
.B(n_951),
.C(n_900),
.D(n_891),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_958),
.Y(n_965)
);

OAI322xp33_ASAP7_75t_L g966 ( 
.A1(n_960),
.A2(n_949),
.A3(n_931),
.B1(n_919),
.B2(n_883),
.C1(n_904),
.C2(n_878),
.Y(n_966)
);

AOI311xp33_ASAP7_75t_L g967 ( 
.A1(n_959),
.A2(n_949),
.A3(n_897),
.B(n_903),
.C(n_931),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_965),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_966),
.Y(n_969)
);

AOI221xp5_ASAP7_75t_L g970 ( 
.A1(n_963),
.A2(n_959),
.B1(n_898),
.B2(n_923),
.C(n_902),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_964),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_967),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_968),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_969),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_972),
.B(n_971),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_970),
.A2(n_888),
.B1(n_885),
.B2(n_923),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_970),
.A2(n_923),
.B1(n_888),
.B2(n_126),
.Y(n_977)
);

AO22x2_ASAP7_75t_L g978 ( 
.A1(n_972),
.A2(n_122),
.B1(n_125),
.B2(n_128),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_968),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_973),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_979),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_975),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_977),
.A2(n_130),
.B1(n_134),
.B2(n_135),
.Y(n_983)
);

NOR2x1_ASAP7_75t_L g984 ( 
.A(n_974),
.B(n_138),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_978),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_976),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_985),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_SL g988 ( 
.A1(n_982),
.A2(n_142),
.B(n_143),
.Y(n_988)
);

NAND4xp25_ASAP7_75t_L g989 ( 
.A(n_980),
.B(n_981),
.C(n_986),
.D(n_984),
.Y(n_989)
);

OR2x6_ASAP7_75t_L g990 ( 
.A(n_983),
.B(n_144),
.Y(n_990)
);

AND4x1_ASAP7_75t_L g991 ( 
.A(n_982),
.B(n_145),
.C(n_146),
.D(n_149),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_980),
.B(n_150),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_980),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_980),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_980),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_992),
.B(n_151),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_993),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_994),
.A2(n_152),
.B1(n_153),
.B2(n_156),
.Y(n_998)
);

AO22x2_ASAP7_75t_L g999 ( 
.A1(n_995),
.A2(n_158),
.B1(n_159),
.B2(n_161),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_990),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_989),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_SL g1002 ( 
.A1(n_988),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_1002)
);

INVxp67_ASAP7_75t_SL g1003 ( 
.A(n_987),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_991),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_997),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_999),
.Y(n_1006)
);

AO22x2_ASAP7_75t_L g1007 ( 
.A1(n_1004),
.A2(n_169),
.B1(n_171),
.B2(n_177),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_1003),
.A2(n_178),
.B1(n_181),
.B2(n_183),
.Y(n_1008)
);

INVxp67_ASAP7_75t_SL g1009 ( 
.A(n_996),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_999),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_1001),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1009),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_1005),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1006),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_1010),
.B(n_1000),
.Y(n_1015)
);

OAI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_1013),
.A2(n_1011),
.B1(n_998),
.B2(n_1002),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_1012),
.A2(n_1008),
.B1(n_1007),
.B2(n_193),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1017),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1016),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_1018),
.A2(n_1014),
.B1(n_1015),
.B2(n_194),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_1019),
.A2(n_191),
.B1(n_192),
.B2(n_198),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1020),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1021),
.Y(n_1023)
);

AOI221xp5_ASAP7_75t_L g1024 ( 
.A1(n_1022),
.A2(n_200),
.B1(n_201),
.B2(n_204),
.C(n_206),
.Y(n_1024)
);

AOI211xp5_ASAP7_75t_L g1025 ( 
.A1(n_1024),
.A2(n_1023),
.B(n_207),
.C(n_208),
.Y(n_1025)
);


endmodule