module fake_jpeg_14868_n_128 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_128);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx24_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_31),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_33),
.B(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_39),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_2),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_44),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_3),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_16),
.Y(n_52)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_21),
.B(n_4),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_5),
.C(n_8),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_27),
.A2(n_4),
.B1(n_5),
.B2(n_10),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_14),
.B1(n_19),
.B2(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_13),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_60),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_27),
.B1(n_21),
.B2(n_17),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_54),
.B1(n_30),
.B2(n_29),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_53),
.Y(n_73)
);

NOR2x1_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_63),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_18),
.B1(n_19),
.B2(n_24),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_69),
.B1(n_56),
.B2(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_13),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_24),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_6),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_68),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_59),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_55),
.B1(n_84),
.B2(n_70),
.Y(n_96)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_32),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_76),
.C(n_83),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_35),
.B(n_6),
.C(n_44),
.Y(n_75)
);

FAx1_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_62),
.CI(n_46),
.CON(n_91),
.SN(n_91)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_35),
.C(n_36),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_60),
.B(n_61),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_48),
.B(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_86),
.Y(n_100)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_84),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_48),
.C(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_51),
.B(n_57),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_63),
.B(n_46),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_90),
.B(n_96),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_87),
.B(n_89),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_85),
.A2(n_77),
.B1(n_76),
.B2(n_83),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_95),
.B1(n_96),
.B2(n_73),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_55),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_94),
.B(n_88),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_82),
.A2(n_55),
.B1(n_65),
.B2(n_81),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_72),
.C(n_78),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_104),
.C(n_106),
.Y(n_113)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_SL g110 ( 
.A(n_108),
.B(n_109),
.C(n_91),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_92),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_88),
.C(n_109),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_114),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_106),
.C(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_121),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_116),
.A2(n_103),
.B1(n_91),
.B2(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_120),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_97),
.C(n_93),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_98),
.C(n_123),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_126),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_122),
.B(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);


endmodule