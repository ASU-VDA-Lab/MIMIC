module fake_jpeg_11134_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx5_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_6),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

AO22x1_ASAP7_75t_SL g19 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_19)
);

A2O1A1O1Ixp25_ASAP7_75t_L g38 ( 
.A1(n_19),
.A2(n_1),
.B(n_4),
.C(n_23),
.D(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_15),
.A2(n_17),
.B1(n_14),
.B2(n_10),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_17),
.B1(n_18),
.B2(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_28),
.B1(n_26),
.B2(n_24),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_35),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_19),
.Y(n_42)
);

FAx1_ASAP7_75t_SL g40 ( 
.A(n_19),
.B(n_22),
.CI(n_29),
.CON(n_40),
.SN(n_40)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_37),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_31),
.B1(n_34),
.B2(n_39),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_35),
.B(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_51),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_41),
.B1(n_34),
.B2(n_43),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_42),
.B1(n_40),
.B2(n_44),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_42),
.B1(n_47),
.B2(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_54),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_50),
.B(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_52),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_57),
.A2(n_58),
.B(n_41),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_59),
.A2(n_39),
.B(n_36),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_36),
.Y(n_61)
);


endmodule