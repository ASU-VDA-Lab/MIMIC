module fake_netlist_5_2580_n_656 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_656);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_656;

wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_619;
wire n_408;
wire n_376;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_483;
wire n_544;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_280;
wire n_590;
wire n_629;
wire n_378;
wire n_551;
wire n_581;
wire n_382;
wire n_554;
wire n_254;
wire n_583;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_455;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_507;
wire n_497;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_506;
wire n_610;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_307;
wire n_633;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_546;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_264;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_584;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_311;
wire n_208;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_638;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_627;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_180;
wire n_560;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_572;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_269;
wire n_529;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_644;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_262;
wire n_238;
wire n_639;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_278;

INVx2_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_68),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_89),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_25),
.Y(n_146)
);

BUFx2_ASAP7_75t_SL g147 ( 
.A(n_103),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_75),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_56),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_107),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_18),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_21),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_30),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_41),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_91),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_35),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_95),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_108),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_34),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_122),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_22),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_33),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_102),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_106),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_24),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_70),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_66),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_13),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_13),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_20),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_60),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_9),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_15),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_61),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_52),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_36),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_80),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_12),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_43),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_11),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_11),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_137),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_71),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_8),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_77),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_94),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_129),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_121),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_50),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_23),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_39),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_64),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_47),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_74),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_59),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_16),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_40),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_9),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_26),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_67),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_132),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_0),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_0),
.Y(n_219)
);

BUFx8_ASAP7_75t_SL g220 ( 
.A(n_149),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_1),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_1),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_2),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_143),
.Y(n_224)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_143),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_152),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_174),
.Y(n_228)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_152),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_176),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_2),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_151),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_185),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_153),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_155),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_184),
.B(n_3),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_158),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_160),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_186),
.B(n_3),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_4),
.Y(n_240)
);

CKINVDCx6p67_ASAP7_75t_R g241 ( 
.A(n_149),
.Y(n_241)
);

BUFx8_ASAP7_75t_L g242 ( 
.A(n_161),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_163),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_165),
.Y(n_244)
);

CKINVDCx6p67_ASAP7_75t_R g245 ( 
.A(n_150),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_173),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_188),
.B(n_4),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_178),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_147),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_179),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_187),
.B(n_5),
.Y(n_251)
);

AND2x4_ASAP7_75t_L g252 ( 
.A(n_195),
.B(n_14),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_5),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

AND2x4_ASAP7_75t_L g255 ( 
.A(n_210),
.B(n_17),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_150),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_144),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_145),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_168),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_221),
.A2(n_168),
.B1(n_192),
.B2(n_207),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_175),
.B1(n_208),
.B2(n_205),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_146),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_219),
.A2(n_172),
.B1(n_202),
.B2(n_201),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_148),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_220),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_154),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g267 ( 
.A1(n_228),
.A2(n_211),
.B1(n_200),
.B2(n_198),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_L g268 ( 
.A1(n_222),
.A2(n_197),
.B1(n_196),
.B2(n_193),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_156),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_157),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_231),
.A2(n_189),
.B1(n_183),
.B2(n_182),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_L g273 ( 
.A1(n_236),
.A2(n_180),
.B1(n_171),
.B2(n_170),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_256),
.A2(n_169),
.B1(n_167),
.B2(n_166),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_164),
.B1(n_162),
.B2(n_159),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_227),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_R g277 ( 
.A1(n_215),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_19),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_227),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_219),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_220),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_227),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_248),
.B(n_10),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_223),
.B(n_12),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_216),
.B(n_27),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_216),
.B(n_28),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_223),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_240),
.A2(n_253),
.B1(n_247),
.B2(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_256),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_240),
.A2(n_37),
.B1(n_38),
.B2(n_42),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_227),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_247),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_249),
.B(n_48),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_257),
.B(n_49),
.Y(n_294)
);

NOR2x1p5_ASAP7_75t_L g295 ( 
.A(n_241),
.B(n_51),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_253),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_249),
.B(n_57),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_252),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_218),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_218),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_249),
.B(n_65),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_249),
.B(n_69),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_241),
.A2(n_245),
.B1(n_255),
.B2(n_252),
.Y(n_303)
);

AO22x2_ASAP7_75t_L g304 ( 
.A1(n_252),
.A2(n_72),
.B1(n_73),
.B2(n_76),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_R g305 ( 
.A1(n_217),
.A2(n_78),
.B1(n_81),
.B2(n_82),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_R g306 ( 
.A1(n_226),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_218),
.B(n_87),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_218),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_245),
.A2(n_88),
.B1(n_90),
.B2(n_93),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_L g310 ( 
.A1(n_234),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_255),
.A2(n_100),
.B1(n_101),
.B2(n_104),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_269),
.B(n_270),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_265),
.B(n_257),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_271),
.B(n_257),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_264),
.B(n_266),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_260),
.Y(n_317)
);

BUFx6f_ASAP7_75t_SL g318 ( 
.A(n_281),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_300),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_274),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_285),
.B(n_229),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_282),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_260),
.B(n_257),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_279),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_261),
.B(n_263),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_262),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_289),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_257),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_286),
.B(n_225),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_249),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_105),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_288),
.B(n_235),
.Y(n_335)
);

HAxp5_ASAP7_75t_SL g336 ( 
.A(n_309),
.B(n_244),
.CON(n_336),
.SN(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_307),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_283),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_278),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_284),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_293),
.Y(n_341)
);

INVx4_ASAP7_75t_SL g342 ( 
.A(n_297),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_298),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_311),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_301),
.Y(n_345)
);

INVx4_ASAP7_75t_SL g346 ( 
.A(n_305),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_304),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_263),
.A2(n_237),
.B(n_243),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_261),
.B(n_242),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_304),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_273),
.B(n_225),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_275),
.B(n_109),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_272),
.B(n_237),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_287),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_268),
.B(n_225),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_302),
.Y(n_356)
);

XNOR2x2_ASAP7_75t_L g357 ( 
.A(n_280),
.B(n_214),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_295),
.B(n_213),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_292),
.Y(n_360)
);

BUFx8_ASAP7_75t_L g361 ( 
.A(n_277),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_294),
.B(n_225),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_296),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_310),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_306),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_267),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_299),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_299),
.Y(n_368)
);

INVx4_ASAP7_75t_SL g369 ( 
.A(n_274),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_299),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_285),
.A2(n_225),
.B(n_229),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_264),
.B(n_242),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_282),
.Y(n_373)
);

XOR2x2_ASAP7_75t_L g374 ( 
.A(n_260),
.B(n_242),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_264),
.B(n_238),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_299),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_299),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_312),
.B(n_238),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_324),
.Y(n_379)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_342),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_111),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_329),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_373),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_348),
.B(n_243),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_348),
.B(n_214),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_315),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_316),
.B(n_250),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_254),
.Y(n_388)
);

OR2x2_ASAP7_75t_SL g389 ( 
.A(n_365),
.B(n_366),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_353),
.B(n_213),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_326),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_340),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_367),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_337),
.B(n_246),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_357),
.Y(n_396)
);

AND2x2_ASAP7_75t_SL g397 ( 
.A(n_327),
.B(n_254),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_328),
.B(n_250),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_325),
.B(n_246),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_335),
.B(n_338),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_333),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_364),
.Y(n_402)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_342),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_319),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_359),
.B(n_246),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_356),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_341),
.A2(n_229),
.B(n_224),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_359),
.B(n_224),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_347),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_345),
.B(n_254),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_339),
.B(n_224),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_363),
.B(n_250),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_322),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_368),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_323),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_370),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_344),
.B(n_250),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_377),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_376),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_313),
.Y(n_420)
);

AND2x6_ASAP7_75t_L g421 ( 
.A(n_350),
.B(n_254),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_318),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_354),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_351),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_358),
.B(n_254),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_360),
.B(n_229),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_321),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_321),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_317),
.B(n_229),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_330),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_331),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_331),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_320),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_372),
.B(n_114),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_362),
.A2(n_115),
.B(n_116),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_349),
.B(n_117),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_332),
.B(n_118),
.Y(n_438)
);

AND2x2_ASAP7_75t_SL g439 ( 
.A(n_336),
.B(n_119),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_332),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_346),
.B(n_120),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_382),
.Y(n_442)
);

OR2x6_ASAP7_75t_L g443 ( 
.A(n_403),
.B(n_318),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_382),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_422),
.Y(n_445)
);

OR2x6_ASAP7_75t_L g446 ( 
.A(n_403),
.B(n_334),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_369),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_416),
.B(n_369),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_384),
.B(n_346),
.Y(n_449)
);

BUFx12f_ASAP7_75t_L g450 ( 
.A(n_422),
.Y(n_450)
);

OR2x6_ASAP7_75t_L g451 ( 
.A(n_403),
.B(n_352),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_389),
.B(n_374),
.Y(n_452)
);

NAND2x1p5_ASAP7_75t_L g453 ( 
.A(n_380),
.B(n_371),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_379),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_387),
.B(n_123),
.Y(n_455)
);

INVx6_ASAP7_75t_L g456 ( 
.A(n_393),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_380),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_400),
.B(n_126),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_423),
.B(n_361),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_402),
.B(n_361),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_430),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_409),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_400),
.B(n_378),
.Y(n_463)
);

OR2x6_ASAP7_75t_L g464 ( 
.A(n_380),
.B(n_128),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_380),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_415),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_391),
.B(n_130),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_389),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_415),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_384),
.B(n_133),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_378),
.B(n_134),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_406),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_404),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_406),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_391),
.B(n_135),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_425),
.B(n_397),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_390),
.B(n_136),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_430),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_396),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_404),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_390),
.B(n_139),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_425),
.B(n_140),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_392),
.B(n_423),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_413),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_412),
.B(n_141),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_463),
.B(n_417),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_417),
.Y(n_487)
);

BUFx4f_ASAP7_75t_L g488 ( 
.A(n_457),
.Y(n_488)
);

NAND2x1p5_ASAP7_75t_L g489 ( 
.A(n_457),
.B(n_381),
.Y(n_489)
);

INVx6_ASAP7_75t_SL g490 ( 
.A(n_443),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_456),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_444),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_483),
.B(n_434),
.Y(n_493)
);

INVx5_ASAP7_75t_L g494 ( 
.A(n_457),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_449),
.B(n_424),
.Y(n_495)
);

AO21x1_ASAP7_75t_L g496 ( 
.A1(n_476),
.A2(n_437),
.B(n_470),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_465),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_465),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_456),
.Y(n_499)
);

BUFx12f_ASAP7_75t_L g500 ( 
.A(n_443),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_465),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_472),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_454),
.Y(n_503)
);

BUFx2_ASAP7_75t_SL g504 ( 
.A(n_444),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_442),
.Y(n_505)
);

BUFx6f_ASAP7_75t_SL g506 ( 
.A(n_443),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_468),
.Y(n_507)
);

INVx8_ASAP7_75t_L g508 ( 
.A(n_464),
.Y(n_508)
);

INVx3_ASAP7_75t_SL g509 ( 
.A(n_445),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_466),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_447),
.B(n_448),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_472),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_479),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_469),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_449),
.Y(n_515)
);

INVx6_ASAP7_75t_L g516 ( 
.A(n_505),
.Y(n_516)
);

BUFx8_ASAP7_75t_SL g517 ( 
.A(n_507),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_493),
.A2(n_439),
.B1(n_452),
.B2(n_478),
.Y(n_518)
);

BUFx12f_ASAP7_75t_L g519 ( 
.A(n_500),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_515),
.A2(n_439),
.B1(n_461),
.B2(n_478),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_486),
.A2(n_439),
.B1(n_485),
.B2(n_381),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_510),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_486),
.A2(n_441),
.B(n_460),
.Y(n_523)
);

OAI22xp33_ASAP7_75t_L g524 ( 
.A1(n_513),
.A2(n_431),
.B1(n_451),
.B2(n_434),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_495),
.A2(n_381),
.B1(n_435),
.B2(n_447),
.Y(n_525)
);

NAND2x1p5_ASAP7_75t_L g526 ( 
.A(n_494),
.B(n_472),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_492),
.A2(n_431),
.B1(n_446),
.B2(n_451),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_491),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_510),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_495),
.A2(n_381),
.B1(n_435),
.B2(n_448),
.Y(n_530)
);

INVx6_ASAP7_75t_L g531 ( 
.A(n_505),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_491),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_514),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_503),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_503),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_494),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_487),
.Y(n_537)
);

BUFx12f_ASAP7_75t_L g538 ( 
.A(n_500),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_509),
.Y(n_539)
);

OAI22xp33_ASAP7_75t_L g540 ( 
.A1(n_508),
.A2(n_451),
.B1(n_386),
.B2(n_446),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_509),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_494),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_536),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_525),
.B(n_397),
.Y(n_544)
);

OAI21xp33_ASAP7_75t_SL g545 ( 
.A1(n_530),
.A2(n_397),
.B(n_438),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_536),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_521),
.A2(n_424),
.B1(n_458),
.B2(n_426),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_SL g548 ( 
.A1(n_527),
.A2(n_508),
.B1(n_441),
.B2(n_504),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_542),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_518),
.A2(n_489),
.B1(n_440),
.B2(n_508),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_527),
.A2(n_426),
.B1(n_459),
.B2(n_471),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_520),
.A2(n_426),
.B1(n_508),
.B2(n_477),
.Y(n_552)
);

BUFx4f_ASAP7_75t_SL g553 ( 
.A(n_539),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_SL g554 ( 
.A1(n_537),
.A2(n_506),
.B1(n_464),
.B2(n_446),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_524),
.A2(n_426),
.B1(n_481),
.B2(n_496),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_529),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_522),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_540),
.A2(n_426),
.B1(n_393),
.B2(n_394),
.Y(n_558)
);

BUFx4f_ASAP7_75t_SL g559 ( 
.A(n_541),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_519),
.A2(n_394),
.B1(n_419),
.B2(n_428),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_538),
.A2(n_419),
.B1(n_428),
.B2(n_433),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_534),
.B(n_385),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_SL g563 ( 
.A1(n_523),
.A2(n_506),
.B1(n_464),
.B2(n_436),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_516),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_516),
.A2(n_419),
.B1(n_433),
.B2(n_398),
.Y(n_565)
);

AOI222xp33_ASAP7_75t_L g566 ( 
.A1(n_523),
.A2(n_418),
.B1(n_420),
.B2(n_395),
.C1(n_484),
.C2(n_473),
.Y(n_566)
);

BUFx4f_ASAP7_75t_SL g567 ( 
.A(n_532),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_535),
.B(n_385),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_531),
.A2(n_418),
.B1(n_429),
.B2(n_432),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_531),
.A2(n_489),
.B1(n_488),
.B2(n_480),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_533),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_526),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_SL g573 ( 
.A1(n_542),
.A2(n_506),
.B1(n_470),
.B2(n_399),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_566),
.A2(n_399),
.B1(n_395),
.B2(n_411),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_557),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_SL g576 ( 
.A1(n_545),
.A2(n_455),
.B1(n_475),
.B2(n_467),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_551),
.A2(n_548),
.B1(n_558),
.B2(n_554),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_562),
.B(n_511),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_550),
.A2(n_467),
.B1(n_475),
.B2(n_482),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_563),
.A2(n_490),
.B1(n_511),
.B2(n_488),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_556),
.B(n_511),
.Y(n_581)
);

OAI22xp33_ASAP7_75t_L g582 ( 
.A1(n_544),
.A2(n_414),
.B1(n_490),
.B2(n_450),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_544),
.A2(n_429),
.B1(n_432),
.B2(n_411),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_571),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_555),
.A2(n_413),
.B1(n_414),
.B2(n_405),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_SL g586 ( 
.A1(n_570),
.A2(n_438),
.B1(n_488),
.B2(n_494),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_562),
.B(n_462),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_547),
.A2(n_405),
.B1(n_408),
.B2(n_401),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_557),
.Y(n_589)
);

OAI211xp5_ASAP7_75t_L g590 ( 
.A1(n_560),
.A2(n_409),
.B(n_528),
.C(n_388),
.Y(n_590)
);

OAI22xp33_ASAP7_75t_L g591 ( 
.A1(n_553),
.A2(n_490),
.B1(n_532),
.B2(n_391),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_556),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_561),
.A2(n_532),
.B1(n_499),
.B2(n_526),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_568),
.Y(n_594)
);

INVxp67_ASAP7_75t_SL g595 ( 
.A(n_568),
.Y(n_595)
);

OAI22xp33_ASAP7_75t_L g596 ( 
.A1(n_559),
.A2(n_499),
.B1(n_406),
.B2(n_474),
.Y(n_596)
);

NAND3xp33_ASAP7_75t_L g597 ( 
.A(n_577),
.B(n_552),
.C(n_573),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_587),
.B(n_564),
.Y(n_598)
);

NAND2x1_ASAP7_75t_L g599 ( 
.A(n_589),
.B(n_546),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_595),
.B(n_572),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_584),
.Y(n_601)
);

NAND4xp25_ASAP7_75t_L g602 ( 
.A(n_574),
.B(n_569),
.C(n_565),
.D(n_408),
.Y(n_602)
);

OAI221xp5_ASAP7_75t_L g603 ( 
.A1(n_579),
.A2(n_401),
.B1(n_383),
.B2(n_546),
.C(n_543),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_594),
.B(n_546),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_578),
.B(n_543),
.Y(n_605)
);

AOI221xp5_ASAP7_75t_L g606 ( 
.A1(n_582),
.A2(n_383),
.B1(n_427),
.B2(n_379),
.C(n_406),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_575),
.B(n_543),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_592),
.B(n_549),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_581),
.B(n_549),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_591),
.B(n_580),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_586),
.B(n_549),
.Y(n_611)
);

OR2x2_ASAP7_75t_L g612 ( 
.A(n_601),
.B(n_583),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_597),
.A2(n_576),
.B1(n_574),
.B2(n_585),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_600),
.B(n_590),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_607),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_L g616 ( 
.A(n_597),
.B(n_585),
.C(n_593),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_604),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_609),
.B(n_596),
.Y(n_618)
);

NAND4xp75_ASAP7_75t_L g619 ( 
.A(n_610),
.B(n_427),
.C(n_567),
.D(n_517),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_615),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_617),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_612),
.Y(n_622)
);

NAND4xp75_ASAP7_75t_L g623 ( 
.A(n_618),
.B(n_611),
.C(n_608),
.D(n_606),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_614),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_616),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_613),
.B(n_598),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_622),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_L g628 ( 
.A(n_626),
.B(n_619),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_622),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_624),
.B(n_605),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_621),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_627),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_631),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_629),
.Y(n_634)
);

AOI22x1_ASAP7_75t_L g635 ( 
.A1(n_628),
.A2(n_625),
.B1(n_620),
.B2(n_623),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_630),
.Y(n_636)
);

OAI322xp33_ASAP7_75t_L g637 ( 
.A1(n_635),
.A2(n_626),
.A3(n_630),
.B1(n_603),
.B2(n_599),
.C1(n_602),
.C2(n_410),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_633),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_632),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_639),
.A2(n_636),
.B1(n_634),
.B2(n_588),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_638),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_641),
.A2(n_637),
.B1(n_636),
.B2(n_588),
.Y(n_642)
);

AOI31xp33_ASAP7_75t_L g643 ( 
.A1(n_642),
.A2(n_640),
.A3(n_453),
.B(n_407),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_643),
.A2(n_421),
.B1(n_502),
.B2(n_406),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_644),
.A2(n_421),
.B1(n_498),
.B2(n_497),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_645),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_646),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_647),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_SL g649 ( 
.A1(n_648),
.A2(n_421),
.B1(n_498),
.B2(n_497),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_649),
.Y(n_650)
);

OAI22xp33_ASAP7_75t_L g651 ( 
.A1(n_650),
.A2(n_498),
.B1(n_497),
.B2(n_512),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_650),
.A2(n_512),
.B1(n_421),
.B2(n_498),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_652),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_651),
.Y(n_654)
);

AOI221xp5_ASAP7_75t_L g655 ( 
.A1(n_654),
.A2(n_497),
.B1(n_512),
.B2(n_501),
.C(n_502),
.Y(n_655)
);

AOI211xp5_ASAP7_75t_L g656 ( 
.A1(n_655),
.A2(n_653),
.B(n_512),
.C(n_142),
.Y(n_656)
);


endmodule