module fake_aes_1033_n_42 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_42);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_33;
wire n_30;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
NAND2xp33_ASAP7_75t_L g11 ( .A(n_3), .B(n_4), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_1), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_10), .Y(n_13) );
NOR2xp33_ASAP7_75t_R g14 ( .A(n_5), .B(n_9), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_5), .B(n_2), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_1), .B(n_4), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_3), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_18), .B(n_0), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_13), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_12), .B(n_2), .Y(n_22) );
AOI22xp5_ASAP7_75t_L g23 ( .A1(n_11), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_23) );
OR2x2_ASAP7_75t_L g24 ( .A(n_17), .B(n_6), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_19), .Y(n_25) );
NOR2x1p5_ASAP7_75t_L g26 ( .A(n_24), .B(n_17), .Y(n_26) );
OAI22xp5_ASAP7_75t_SL g27 ( .A1(n_23), .A2(n_15), .B1(n_16), .B2(n_14), .Y(n_27) );
AND2x4_ASAP7_75t_L g28 ( .A(n_19), .B(n_20), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_25), .Y(n_29) );
AND4x1_ASAP7_75t_L g30 ( .A(n_27), .B(n_23), .C(n_22), .D(n_21), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
INVx2_ASAP7_75t_SL g32 ( .A(n_31), .Y(n_32) );
HB1xp67_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_33), .B(n_26), .Y(n_34) );
OR2x2_ASAP7_75t_L g35 ( .A(n_32), .B(n_25), .Y(n_35) );
AND2x4_ASAP7_75t_L g36 ( .A(n_34), .B(n_30), .Y(n_36) );
NOR2x1_ASAP7_75t_L g37 ( .A(n_35), .B(n_28), .Y(n_37) );
OAI22xp5_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_32), .B1(n_29), .B2(n_28), .Y(n_38) );
INVx2_ASAP7_75t_L g39 ( .A(n_37), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_36), .Y(n_40) );
BUFx2_ASAP7_75t_L g41 ( .A(n_39), .Y(n_41) );
OAI22xp5_ASAP7_75t_L g42 ( .A1(n_41), .A2(n_40), .B1(n_39), .B2(n_38), .Y(n_42) );
endmodule