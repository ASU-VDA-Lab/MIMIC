module fake_jpeg_11203_n_578 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_578);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_578;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_0),
.B(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_57),
.Y(n_150)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_58),
.Y(n_156)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_60),
.Y(n_175)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_23),
.B(n_10),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_67),
.B(n_70),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_23),
.B(n_10),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_25),
.A2(n_11),
.B1(n_17),
.B2(n_16),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_82),
.A2(n_25),
.B1(n_20),
.B2(n_27),
.Y(n_135)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_83),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_40),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_104),
.Y(n_115)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_89),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_93),
.Y(n_168)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_44),
.B(n_11),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_95),
.B(n_99),
.Y(n_169)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_97),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_44),
.B(n_9),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_108),
.Y(n_134)
);

BUFx8_ASAP7_75t_L g106 ( 
.A(n_20),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_107),
.Y(n_128)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_20),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_25),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_67),
.B(n_24),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_131),
.B(n_143),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_135),
.A2(n_27),
.B1(n_31),
.B2(n_72),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_70),
.B(n_24),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_24),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_148),
.B(n_165),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_58),
.A2(n_46),
.B1(n_41),
.B2(n_40),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_149),
.A2(n_155),
.B1(n_158),
.B2(n_167),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_47),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_152),
.B(n_160),
.Y(n_215)
);

AO22x1_ASAP7_75t_SL g155 ( 
.A1(n_82),
.A2(n_40),
.B1(n_38),
.B2(n_31),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_65),
.A2(n_41),
.B1(n_46),
.B2(n_53),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_64),
.B(n_47),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_106),
.B(n_53),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_33),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_68),
.B(n_49),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_128),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_66),
.B(n_45),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_90),
.A2(n_46),
.B1(n_41),
.B2(n_31),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_79),
.B(n_42),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_172),
.B(n_176),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_71),
.B(n_47),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_173),
.B(n_32),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_80),
.B(n_45),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_27),
.B(n_36),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_177),
.A2(n_21),
.B(n_35),
.Y(n_261)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_178),
.Y(n_267)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_180),
.Y(n_250)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_182),
.Y(n_284)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_183),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_149),
.A2(n_85),
.B1(n_93),
.B2(n_97),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_184),
.A2(n_187),
.B1(n_197),
.B2(n_213),
.Y(n_258)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_185),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_96),
.B1(n_98),
.B2(n_89),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_186),
.A2(n_117),
.B1(n_175),
.B2(n_145),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_100),
.B1(n_60),
.B2(n_57),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_137),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_188),
.Y(n_291)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

INVx3_ASAP7_75t_SL g285 ( 
.A(n_191),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_210),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_193),
.Y(n_294)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_194),
.Y(n_286)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_196),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_123),
.A2(n_42),
.B1(n_33),
.B2(n_45),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_198),
.Y(n_262)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_199),
.Y(n_248)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_200),
.Y(n_269)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_130),
.Y(n_201)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_201),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_202),
.B(n_205),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_204),
.A2(n_21),
.B1(n_52),
.B2(n_36),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_126),
.B(n_140),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_115),
.B(n_53),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_206),
.Y(n_266)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_120),
.Y(n_208)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_208),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_146),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_209),
.Y(n_263)
);

AND2x2_ASAP7_75t_SL g210 ( 
.A(n_124),
.B(n_31),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_134),
.Y(n_211)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_211),
.Y(n_282)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_212),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_42),
.B1(n_33),
.B2(n_46),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_214),
.B(n_219),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_155),
.A2(n_19),
.B1(n_51),
.B2(n_48),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_217),
.A2(n_220),
.B1(n_222),
.B2(n_52),
.Y(n_281)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_171),
.Y(n_218)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_218),
.Y(n_295)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_146),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_119),
.A2(n_19),
.B1(n_51),
.B2(n_48),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_163),
.B(n_38),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_221),
.B(n_224),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_116),
.A2(n_38),
.B1(n_36),
.B2(n_35),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_139),
.B(n_19),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_223),
.Y(n_273)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_127),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_130),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_225),
.B(n_226),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_116),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_157),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_227),
.Y(n_242)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_228),
.Y(n_244)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_153),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_229),
.Y(n_271)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_150),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_230),
.A2(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_231),
.A2(n_122),
.B1(n_114),
.B2(n_39),
.Y(n_243)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_153),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_232),
.Y(n_246)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_151),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_233),
.Y(n_270)
);

O2A1O1Ixp33_ASAP7_75t_SL g234 ( 
.A1(n_142),
.A2(n_16),
.B(n_18),
.C(n_17),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_234),
.A2(n_43),
.B(n_39),
.C(n_34),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_144),
.B(n_32),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_238),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_122),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_129),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_133),
.B(n_32),
.Y(n_238)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_129),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_114),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_240),
.A2(n_43),
.B1(n_39),
.B2(n_34),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_243),
.B(n_0),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_249),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_297)
);

AO22x1_ASAP7_75t_SL g251 ( 
.A1(n_181),
.A2(n_117),
.B1(n_119),
.B2(n_145),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_251),
.B(n_201),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_141),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_253),
.B(n_264),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_216),
.A2(n_136),
.B1(n_132),
.B2(n_156),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_186),
.A2(n_136),
.B1(n_132),
.B2(n_156),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_204),
.A2(n_175),
.B1(n_113),
.B2(n_48),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_260),
.A2(n_288),
.B1(n_222),
.B2(n_210),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_261),
.A2(n_287),
.B(n_292),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_190),
.B(n_122),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_177),
.A2(n_113),
.B(n_52),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_268),
.A2(n_221),
.B(n_219),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_SL g277 ( 
.A(n_207),
.B(n_51),
.C(n_43),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_277),
.B(n_287),
.Y(n_346)
);

AO21x1_ASAP7_75t_L g347 ( 
.A1(n_278),
.A2(n_277),
.B(n_265),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_280),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_230),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_184),
.A2(n_34),
.B1(n_35),
.B2(n_21),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_283),
.A2(n_285),
.B1(n_242),
.B2(n_273),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_203),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_203),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_214),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_257),
.A2(n_236),
.B1(n_194),
.B2(n_226),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_298),
.A2(n_310),
.B1(n_321),
.B2(n_341),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_263),
.Y(n_299)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_299),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_300),
.B(n_342),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_258),
.A2(n_205),
.B1(n_210),
.B2(n_191),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_301),
.A2(n_302),
.B1(n_311),
.B2(n_312),
.Y(n_349)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_258),
.A2(n_234),
.B1(n_228),
.B2(n_237),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_253),
.B(n_264),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_303),
.B(n_295),
.C(n_289),
.Y(n_359)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_248),
.Y(n_304)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_252),
.B(n_192),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_305),
.B(n_327),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_306),
.A2(n_291),
.B1(n_286),
.B2(n_296),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_307),
.A2(n_319),
.B(n_335),
.Y(n_373)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_255),
.Y(n_308)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_308),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_294),
.A2(n_209),
.B1(n_239),
.B2(n_225),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_281),
.A2(n_224),
.B1(n_208),
.B2(n_199),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_243),
.A2(n_196),
.B1(n_188),
.B2(n_240),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_313),
.A2(n_315),
.B1(n_325),
.B2(n_338),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_0),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_314),
.B(n_318),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_251),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_274),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_316),
.B(n_322),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_279),
.B(n_9),
.Y(n_318)
);

XNOR2x2_ASAP7_75t_L g319 ( 
.A(n_241),
.B(n_9),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_255),
.Y(n_320)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_320),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_294),
.A2(n_8),
.B1(n_14),
.B2(n_5),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_268),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_323),
.Y(n_354)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_245),
.Y(n_324)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_324),
.Y(n_376)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_245),
.Y(n_326)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_326),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_267),
.B(n_5),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_262),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_328),
.B(n_332),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_241),
.B(n_4),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_329),
.B(n_331),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_251),
.A2(n_6),
.B1(n_12),
.B2(n_13),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_330),
.A2(n_285),
.B1(n_244),
.B2(n_275),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_267),
.B(n_6),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_262),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_241),
.B(n_4),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_333),
.B(n_343),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_261),
.A2(n_18),
.B(n_6),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_335),
.A2(n_344),
.B(n_291),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_282),
.B(n_6),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_337),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_274),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_266),
.A2(n_4),
.B1(n_13),
.B2(n_12),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_282),
.B(n_13),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_339),
.B(n_340),
.Y(n_379)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_269),
.Y(n_340)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_248),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_269),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_266),
.B(n_278),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_265),
.A2(n_272),
.B(n_292),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_242),
.B(n_244),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_345),
.Y(n_390)
);

XNOR2x1_ASAP7_75t_SL g353 ( 
.A(n_346),
.B(n_265),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_284),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_345),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_350),
.B(n_383),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_353),
.B(n_333),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_355),
.A2(n_367),
.B1(n_372),
.B2(n_377),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_301),
.A2(n_256),
.B1(n_254),
.B2(n_288),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_357),
.A2(n_388),
.B1(n_297),
.B2(n_324),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_359),
.B(n_374),
.C(n_378),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_343),
.A2(n_274),
.B(n_270),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_362),
.A2(n_385),
.B(n_331),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_366),
.A2(n_368),
.B(n_371),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_322),
.A2(n_285),
.B1(n_286),
.B2(n_289),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_307),
.A2(n_259),
.B(n_276),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_311),
.A2(n_295),
.B1(n_276),
.B2(n_250),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_373),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_303),
.B(n_334),
.C(n_305),
.Y(n_374)
);

AO22x1_ASAP7_75t_L g375 ( 
.A1(n_347),
.A2(n_247),
.B1(n_250),
.B2(n_293),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_375),
.A2(n_382),
.B(n_360),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_300),
.A2(n_247),
.B1(n_293),
.B2(n_290),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_246),
.C(n_271),
.Y(n_378)
);

BUFx8_ASAP7_75t_L g381 ( 
.A(n_316),
.Y(n_381)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_381),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_325),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_317),
.A2(n_263),
.B1(n_296),
.B2(n_259),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_336),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_386),
.B(n_391),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_306),
.A2(n_271),
.B1(n_290),
.B2(n_284),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_297),
.A2(n_347),
.B1(n_330),
.B2(n_306),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_389),
.A2(n_315),
.B1(n_312),
.B2(n_323),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_339),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_369),
.Y(n_392)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_392),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_364),
.B(n_318),
.Y(n_395)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_395),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_396),
.A2(n_417),
.B1(n_420),
.B2(n_377),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_369),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_397),
.B(n_401),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_329),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_412),
.C(n_422),
.Y(n_434)
);

XNOR2x1_ASAP7_75t_L g399 ( 
.A(n_359),
.B(n_346),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_399),
.B(n_406),
.Y(n_442)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_361),
.Y(n_400)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_400),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_367),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_379),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_402),
.B(n_429),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_405),
.A2(n_408),
.B1(n_421),
.B2(n_404),
.Y(n_459)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_361),
.Y(n_407)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_407),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_389),
.A2(n_337),
.B1(n_314),
.B2(n_326),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_363),
.Y(n_409)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_409),
.Y(n_452)
);

AO21x1_ASAP7_75t_L g410 ( 
.A1(n_360),
.A2(n_319),
.B(n_309),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_410),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_353),
.B(n_319),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_411),
.B(n_373),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_365),
.B(n_344),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_350),
.B(n_320),
.Y(n_413)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_413),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_414),
.A2(n_426),
.B(n_381),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_382),
.A2(n_308),
.B1(n_309),
.B2(n_327),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_352),
.A2(n_382),
.B(n_371),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_418),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_342),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_424),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_349),
.A2(n_328),
.B1(n_332),
.B2(n_340),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_360),
.A2(n_304),
.B1(n_341),
.B2(n_338),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_378),
.B(n_299),
.C(n_365),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_352),
.B(n_299),
.C(n_362),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_425),
.C(n_428),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_386),
.B(n_391),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_364),
.B(n_358),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_358),
.B(n_360),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_363),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_430),
.B(n_431),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_403),
.B(n_375),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_432),
.A2(n_438),
.B1(n_454),
.B2(n_457),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_427),
.A2(n_366),
.B(n_375),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_435),
.A2(n_449),
.B(n_416),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_408),
.A2(n_349),
.B1(n_383),
.B2(n_357),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_437),
.A2(n_439),
.B1(n_444),
.B2(n_448),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_396),
.A2(n_355),
.B1(n_372),
.B2(n_354),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_393),
.A2(n_351),
.B1(n_370),
.B2(n_368),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_379),
.Y(n_441)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_441),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_393),
.A2(n_351),
.B1(n_370),
.B2(n_356),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_419),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_445),
.B(n_447),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_394),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_404),
.A2(n_388),
.B1(n_376),
.B2(n_380),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_420),
.A2(n_376),
.B1(n_380),
.B2(n_387),
.Y(n_454)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_394),
.Y(n_455)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_455),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_417),
.A2(n_387),
.B1(n_348),
.B2(n_384),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_459),
.A2(n_424),
.B1(n_405),
.B2(n_426),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_403),
.B(n_381),
.C(n_348),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_460),
.B(n_461),
.C(n_422),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_399),
.B(n_381),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_464),
.B(n_454),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_434),
.B(n_398),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_465),
.B(n_466),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_434),
.B(n_412),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_444),
.A2(n_427),
.B1(n_423),
.B2(n_414),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_467),
.A2(n_477),
.B1(n_448),
.B2(n_433),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_472),
.A2(n_435),
.B(n_453),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_460),
.B(n_428),
.C(n_406),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_473),
.B(n_474),
.C(n_479),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_425),
.C(n_418),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_436),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_475),
.B(n_481),
.Y(n_506)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_443),
.Y(n_476)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_476),
.Y(n_491)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_443),
.Y(n_478)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_478),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_440),
.B(n_411),
.C(n_415),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_436),
.Y(n_480)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_480),
.Y(n_496)
);

XOR2x2_ASAP7_75t_L g481 ( 
.A(n_431),
.B(n_410),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_432),
.A2(n_421),
.B1(n_416),
.B2(n_415),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_483),
.A2(n_488),
.B1(n_439),
.B2(n_437),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_461),
.B(n_384),
.C(n_442),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_484),
.B(n_486),
.C(n_490),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_462),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_485),
.B(n_487),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_442),
.B(n_384),
.C(n_456),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_430),
.B(n_451),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_487),
.B(n_466),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_458),
.A2(n_447),
.B1(n_438),
.B2(n_456),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_441),
.Y(n_489)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_489),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_453),
.B(n_449),
.C(n_458),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_493),
.B(n_513),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_472),
.A2(n_445),
.B(n_457),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_494),
.B(n_508),
.Y(n_518)
);

XNOR2x1_ASAP7_75t_L g528 ( 
.A(n_495),
.B(n_501),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_482),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_497),
.B(n_509),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_499),
.B(n_503),
.C(n_464),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_470),
.B(n_446),
.Y(n_502)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_502),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_465),
.B(n_446),
.C(n_450),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_450),
.Y(n_504)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_504),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_469),
.A2(n_452),
.B1(n_483),
.B2(n_463),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_469),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_477),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_510),
.B(n_511),
.Y(n_533)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_490),
.Y(n_511)
);

FAx1_ASAP7_75t_SL g512 ( 
.A(n_474),
.B(n_452),
.CI(n_481),
.CON(n_512),
.SN(n_512)
);

FAx1_ASAP7_75t_SL g530 ( 
.A(n_512),
.B(n_503),
.CI(n_498),
.CON(n_530),
.SN(n_530)
);

CKINVDCx14_ASAP7_75t_R g527 ( 
.A(n_514),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_515),
.B(n_524),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_505),
.B(n_479),
.C(n_473),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_517),
.B(n_523),
.C(n_531),
.Y(n_536)
);

INVx11_ASAP7_75t_L g519 ( 
.A(n_502),
.Y(n_519)
);

INVx11_ASAP7_75t_L g547 ( 
.A(n_519),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_509),
.A2(n_471),
.B1(n_486),
.B2(n_467),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_522),
.A2(n_526),
.B1(n_506),
.B2(n_493),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_505),
.B(n_468),
.C(n_484),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_500),
.B(n_468),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_513),
.B(n_471),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_525),
.B(n_529),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_510),
.A2(n_507),
.B1(n_496),
.B2(n_504),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_494),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_530),
.B(n_512),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_499),
.B(n_500),
.C(n_498),
.Y(n_531)
);

INVx6_ASAP7_75t_L g534 ( 
.A(n_519),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_534),
.B(n_535),
.Y(n_553)
);

BUFx24_ASAP7_75t_SL g535 ( 
.A(n_530),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_531),
.B(n_508),
.C(n_495),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_537),
.B(n_538),
.Y(n_557)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_520),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_539),
.B(n_544),
.Y(n_554)
);

NAND3xp33_ASAP7_75t_SL g541 ( 
.A(n_532),
.B(n_507),
.C(n_496),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_541),
.A2(n_542),
.B(n_543),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_533),
.A2(n_512),
.B(n_491),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_516),
.B(n_491),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_SL g545 ( 
.A(n_516),
.B(n_492),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_545),
.B(n_518),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_528),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_546),
.B(n_530),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_527),
.B(n_492),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_548),
.B(n_521),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_536),
.B(n_549),
.C(n_537),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_550),
.B(n_556),
.Y(n_561)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_551),
.Y(n_565)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_552),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_549),
.B(n_517),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_558),
.B(n_524),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_543),
.A2(n_515),
.B(n_523),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_559),
.B(n_560),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_534),
.B(n_526),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_551),
.A2(n_539),
.B(n_540),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_563),
.A2(n_564),
.B(n_566),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_557),
.B(n_536),
.C(n_554),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_567),
.A2(n_555),
.B1(n_554),
.B2(n_553),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_568),
.B(n_569),
.Y(n_572)
);

NOR2x1_ASAP7_75t_L g569 ( 
.A(n_562),
.B(n_547),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_564),
.A2(n_560),
.B(n_544),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_571),
.A2(n_561),
.B(n_565),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_573),
.B(n_570),
.C(n_563),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_574),
.B(n_572),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_575),
.B(n_547),
.C(n_545),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_576),
.A2(n_528),
.B(n_518),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_577),
.A2(n_522),
.B(n_525),
.Y(n_578)
);


endmodule