module fake_jpeg_30990_n_524 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_524);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_524;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_53),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_55),
.Y(n_120)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_17),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_60),
.B(n_77),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_70),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_35),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_75),
.Y(n_132)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_25),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_19),
.B(n_0),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_19),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_79),
.B(n_85),
.Y(n_149)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_20),
.B(n_1),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_93),
.Y(n_122)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_94),
.Y(n_119)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_20),
.B(n_1),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_24),
.C(n_45),
.Y(n_107)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_107),
.B(n_148),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_55),
.A2(n_81),
.B1(n_50),
.B2(n_89),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_109),
.A2(n_112),
.B1(n_121),
.B2(n_127),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_37),
.B1(n_21),
.B2(n_43),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_62),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_116),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_56),
.A2(n_37),
.B1(n_21),
.B2(n_43),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_95),
.A2(n_37),
.B1(n_21),
.B2(n_43),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_53),
.A2(n_47),
.B1(n_27),
.B2(n_40),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_130),
.A2(n_145),
.B1(n_150),
.B2(n_152),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_58),
.A2(n_21),
.B1(n_37),
.B2(n_40),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_134),
.A2(n_64),
.B1(n_65),
.B2(n_82),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_78),
.A2(n_22),
.B1(n_45),
.B2(n_44),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_86),
.A2(n_22),
.B1(n_44),
.B2(n_36),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_88),
.A2(n_24),
.B1(n_30),
.B2(n_36),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_90),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_99),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_52),
.A2(n_30),
.B1(n_48),
.B2(n_34),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_155),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_208)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_80),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_92),
.A2(n_37),
.B1(n_21),
.B2(n_47),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_160),
.A2(n_68),
.B1(n_70),
.B2(n_72),
.Y(n_167)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_162),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_153),
.A2(n_94),
.B1(n_97),
.B2(n_93),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_163),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_112),
.A2(n_69),
.B1(n_76),
.B2(n_90),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g257 ( 
.A1(n_164),
.A2(n_167),
.B(n_177),
.Y(n_257)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_166),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_40),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g265 ( 
.A(n_168),
.B(n_197),
.C(n_203),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_147),
.A2(n_61),
.B1(n_54),
.B2(n_59),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_169),
.A2(n_186),
.B1(n_205),
.B2(n_141),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_170),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_118),
.A2(n_71),
.B1(n_63),
.B2(n_98),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_172),
.A2(n_181),
.B1(n_218),
.B2(n_6),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_173),
.Y(n_239)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_176),
.Y(n_240)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_127),
.B1(n_121),
.B2(n_134),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_179),
.Y(n_255)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_180),
.Y(n_269)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_190),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_47),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_184),
.B(n_202),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_66),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_206),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_34),
.B1(n_28),
.B2(n_27),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_109),
.Y(n_190)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_106),
.Y(n_192)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_192),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_120),
.B(n_42),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_194),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_108),
.B(n_42),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_126),
.Y(n_195)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_195),
.Y(n_238)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_196),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_138),
.B(n_34),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_101),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_200),
.Y(n_232)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_140),
.Y(n_199)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_199),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_101),
.B(n_42),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_201),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_116),
.B(n_28),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_117),
.B(n_28),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_125),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_204),
.B(n_207),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_110),
.A2(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_101),
.B(n_2),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_125),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_208),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_124),
.B(n_4),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_104),
.C(n_144),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_131),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_210),
.B(n_213),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_123),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_139),
.A2(n_159),
.B1(n_128),
.B2(n_122),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_212),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_123),
.B(n_42),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_129),
.Y(n_214)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_214),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_119),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_215),
.Y(n_242)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_133),
.Y(n_217)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_217),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_119),
.A2(n_42),
.B1(n_5),
.B2(n_6),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_102),
.Y(n_219)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_136),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_220),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_123),
.B(n_4),
.Y(n_221)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_221),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_166),
.A2(n_115),
.B(n_137),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_228),
.A2(n_173),
.B(n_181),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_231),
.B(n_185),
.Y(n_287)
);

BUFx4f_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_233),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_234),
.B(n_251),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_191),
.A2(n_135),
.B1(n_102),
.B2(n_142),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_236),
.A2(n_243),
.B1(n_250),
.B2(n_267),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_171),
.B(n_115),
.C(n_135),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_241),
.B(n_164),
.C(n_177),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_191),
.A2(n_142),
.B1(n_7),
.B2(n_8),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_190),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_202),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_261),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_216),
.A2(n_7),
.B1(n_10),
.B2(n_13),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_260),
.A2(n_184),
.B1(n_208),
.B2(n_163),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_173),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_211),
.Y(n_266)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_266),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_273),
.A2(n_276),
.B1(n_302),
.B2(n_304),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_168),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_275),
.B(n_280),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_244),
.A2(n_177),
.B1(n_209),
.B2(n_164),
.Y(n_276)
);

NAND3xp33_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_221),
.C(n_206),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_277),
.B(n_290),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_165),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_282),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_224),
.A2(n_177),
.B(n_175),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_279),
.A2(n_252),
.B(n_246),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_232),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_175),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_233),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_283),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_284),
.A2(n_255),
.B(n_252),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_231),
.B(n_204),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_285),
.B(n_293),
.Y(n_342)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_222),
.Y(n_286)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_287),
.B(n_311),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_289),
.B(n_313),
.C(n_318),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_233),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_244),
.A2(n_220),
.B1(n_207),
.B2(n_196),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_291),
.A2(n_254),
.B1(n_227),
.B2(n_258),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_222),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_292),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_242),
.B(n_185),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_228),
.B(n_164),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_294),
.B(n_271),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_253),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_295),
.B(n_306),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_255),
.Y(n_297)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_297),
.Y(n_331)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_298),
.Y(n_351)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_299),
.Y(n_336)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_272),
.Y(n_300)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_300),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_237),
.A2(n_201),
.B1(n_178),
.B2(n_180),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_230),
.B(n_217),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_303),
.B(n_305),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_237),
.A2(n_162),
.B1(n_219),
.B2(n_199),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_230),
.B(n_241),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_226),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_239),
.B(n_261),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_307),
.B(n_308),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_265),
.B(n_189),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_272),
.Y(n_309)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_309),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_239),
.B(n_218),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_310),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_247),
.B(n_214),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_251),
.A2(n_170),
.B1(n_176),
.B2(n_195),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_312),
.A2(n_315),
.B1(n_276),
.B2(n_274),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_247),
.B(n_182),
.C(n_174),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_236),
.B(n_10),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_314),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_257),
.A2(n_192),
.B1(n_13),
.B2(n_14),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_234),
.A2(n_10),
.B1(n_13),
.B2(n_15),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_316),
.A2(n_260),
.B1(n_254),
.B2(n_248),
.Y(n_322)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_268),
.Y(n_317)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_317),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_268),
.B(n_15),
.C(n_16),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_320),
.A2(n_322),
.B1(n_323),
.B2(n_329),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_289),
.A2(n_257),
.B1(n_250),
.B2(n_249),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_324),
.Y(n_390)
);

XOR2x1_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_223),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_328),
.A2(n_332),
.B(n_339),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_281),
.A2(n_249),
.B1(n_238),
.B2(n_240),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_294),
.A2(n_235),
.B(n_266),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_340),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_294),
.A2(n_248),
.B1(n_246),
.B2(n_229),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_341),
.A2(n_346),
.B1(n_284),
.B2(n_281),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_279),
.A2(n_235),
.B(n_225),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_307),
.Y(n_366)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_286),
.Y(n_348)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_348),
.Y(n_364)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_298),
.Y(n_349)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_349),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_285),
.B(n_262),
.C(n_269),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_303),
.C(n_313),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_274),
.A2(n_240),
.B1(n_238),
.B2(n_229),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_354),
.A2(n_359),
.B1(n_296),
.B2(n_283),
.Y(n_372)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_299),
.Y(n_355)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_355),
.Y(n_374)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_300),
.Y(n_356)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_356),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_288),
.B(n_245),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_358),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_274),
.A2(n_245),
.B1(n_269),
.B2(n_15),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_360),
.B(n_365),
.C(n_367),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_345),
.B(n_295),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_362),
.B(n_363),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_327),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_330),
.C(n_347),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_366),
.A2(n_344),
.B(n_339),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_350),
.B(n_287),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_326),
.B(n_278),
.Y(n_368)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_347),
.B(n_282),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_370),
.B(n_324),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_342),
.B(n_288),
.Y(n_371)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_371),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_372),
.A2(n_376),
.B1(n_392),
.B2(n_357),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_323),
.A2(n_312),
.B1(n_315),
.B2(n_273),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_375),
.A2(n_386),
.B1(n_393),
.B2(n_335),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_330),
.B(n_308),
.C(n_293),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_380),
.C(n_382),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_333),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_385),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_353),
.B(n_311),
.C(n_292),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_358),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_381),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_342),
.B(n_302),
.C(n_309),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_346),
.A2(n_314),
.B1(n_316),
.B2(n_310),
.Y(n_383)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_383),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_358),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_345),
.A2(n_304),
.B1(n_290),
.B2(n_317),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_326),
.B(n_296),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_387),
.Y(n_403)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_336),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_388),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_334),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_391),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_335),
.A2(n_318),
.B1(n_301),
.B2(n_16),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_322),
.A2(n_301),
.B1(n_329),
.B2(n_332),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_394),
.A2(n_396),
.B1(n_397),
.B2(n_405),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_367),
.B(n_352),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_412),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_375),
.A2(n_352),
.B1(n_354),
.B2(n_359),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_373),
.A2(n_361),
.B1(n_393),
.B2(n_385),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_398),
.B(n_410),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_399),
.A2(n_400),
.B1(n_364),
.B2(n_384),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_372),
.A2(n_324),
.B1(n_357),
.B2(n_319),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_404),
.B(n_406),
.Y(n_430)
);

A2O1A1Ixp33_ASAP7_75t_SL g405 ( 
.A1(n_389),
.A2(n_340),
.B(n_328),
.C(n_321),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_365),
.B(n_360),
.Y(n_406)
);

OAI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_390),
.A2(n_343),
.B1(n_355),
.B2(n_336),
.Y(n_409)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_409),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_387),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_380),
.B(n_325),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_370),
.B(n_351),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_413),
.B(n_369),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_389),
.A2(n_337),
.B(n_338),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_416),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_366),
.A2(n_390),
.B(n_378),
.Y(n_417)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_417),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_382),
.B(n_368),
.C(n_377),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_419),
.B(n_421),
.C(n_386),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_373),
.B(n_337),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_404),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_331),
.C(n_338),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_428),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_331),
.C(n_379),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_426),
.B(n_441),
.C(n_431),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_418),
.Y(n_427)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_427),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_401),
.B(n_392),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_431),
.B(n_434),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_401),
.B(n_369),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_391),
.Y(n_435)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_435),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_436),
.B(n_443),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_395),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_444),
.Y(n_451)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_415),
.Y(n_439)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_439),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_423),
.Y(n_440)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_440),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_388),
.C(n_364),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_422),
.Y(n_442)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_442),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_420),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_412),
.B(n_374),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_445),
.B(n_413),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_399),
.A2(n_374),
.B1(n_384),
.B2(n_349),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_446),
.B(n_396),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_408),
.B(n_343),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_348),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_433),
.A2(n_400),
.B1(n_403),
.B2(n_407),
.Y(n_449)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_449),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_448),
.Y(n_452)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_452),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_433),
.A2(n_429),
.B1(n_435),
.B2(n_440),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_461),
.Y(n_470)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_438),
.A2(n_416),
.B(n_405),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_456),
.B(n_468),
.Y(n_478)
);

AOI21xp33_ASAP7_75t_L g457 ( 
.A1(n_426),
.A2(n_402),
.B(n_405),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_457),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_SL g463 ( 
.A1(n_432),
.A2(n_405),
.B1(n_397),
.B2(n_398),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_463),
.A2(n_467),
.B1(n_421),
.B2(n_430),
.Y(n_475)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_424),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_465),
.B(n_425),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_466),
.B(n_469),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_441),
.B(n_419),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_449),
.A2(n_394),
.B1(n_428),
.B2(n_445),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_472),
.B(n_473),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_450),
.A2(n_455),
.B(n_453),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_474),
.A2(n_475),
.B(n_478),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_434),
.C(n_437),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_476),
.B(n_483),
.C(n_459),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_430),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_483),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_450),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_479),
.B(n_480),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_425),
.C(n_444),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_462),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_484),
.B(n_485),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_469),
.A2(n_356),
.B1(n_414),
.B2(n_462),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_486),
.B(n_494),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_471),
.B(n_451),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_493),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_476),
.B(n_459),
.C(n_464),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_490),
.B(n_491),
.C(n_477),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_478),
.B(n_451),
.C(n_466),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_492),
.B(n_497),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_470),
.B(n_458),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_470),
.A2(n_460),
.B(n_414),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_495),
.Y(n_499)
);

NOR2xp67_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_458),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_496),
.B(n_498),
.Y(n_502)
);

XOR2x2_ASAP7_75t_SL g497 ( 
.A(n_472),
.B(n_460),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_506),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_481),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_504),
.B(n_505),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_484),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_486),
.B(n_473),
.C(n_480),
.Y(n_506)
);

AOI21x1_ASAP7_75t_L g508 ( 
.A1(n_500),
.A2(n_502),
.B(n_501),
.Y(n_508)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_508),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_507),
.A2(n_497),
.B(n_489),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_511),
.B(n_485),
.Y(n_517)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_507),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_512),
.B(n_513),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_479),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_503),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_516),
.B(n_517),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_514),
.A2(n_513),
.B(n_510),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_519),
.B(n_515),
.C(n_517),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_518),
.Y(n_521)
);

BUFx24_ASAP7_75t_SL g522 ( 
.A(n_521),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_482),
.B1(n_490),
.B2(n_491),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_523),
.B(n_482),
.Y(n_524)
);


endmodule