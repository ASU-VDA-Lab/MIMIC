module fake_jpeg_15913_n_63 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_63);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_63;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

AOI21xp5_ASAP7_75t_L g10 ( 
.A1(n_2),
.A2(n_7),
.B(n_4),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_19),
.C(n_18),
.Y(n_24)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_SL g23 ( 
.A1(n_22),
.A2(n_11),
.B(n_16),
.C(n_17),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_23),
.A2(n_22),
.B1(n_18),
.B2(n_12),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_19),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_20),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_10),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_16),
.B(n_17),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_9),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_33),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_35),
.B1(n_0),
.B2(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_22),
.B1(n_17),
.B2(n_16),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_40),
.B(n_30),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_17),
.B(n_16),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_46),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_30),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_48),
.C(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_42),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_43),
.B(n_3),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_31),
.B(n_2),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_43),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_52),
.C(n_3),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_3),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_55),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_49),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_50),
.Y(n_57)
);

MAJx2_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_55),
.C(n_6),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_5),
.B1(n_8),
.B2(n_57),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_60),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_8),
.Y(n_63)
);


endmodule