module fake_jpeg_189_n_545 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_545);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_545;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_0),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_18),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_12),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_58),
.Y(n_146)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_59),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_32),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_60),
.B(n_65),
.Y(n_134)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_63),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_30),
.B(n_16),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_64),
.B(n_66),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_44),
.B(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_31),
.B(n_15),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_67),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_69),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_27),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_70),
.B(n_77),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_28),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_72),
.B(n_76),
.Y(n_143)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_75),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_28),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_14),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_78),
.B(n_99),
.Y(n_156)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_80),
.Y(n_201)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_81),
.Y(n_171)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_88),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_89),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_90),
.Y(n_202)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_91),
.Y(n_175)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx6_ASAP7_75t_SL g142 ( 
.A(n_94),
.Y(n_142)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_96),
.B(n_115),
.Y(n_158)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_98),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_44),
.B(n_14),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_100),
.Y(n_187)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_101),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_102),
.Y(n_203)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_107),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_110),
.Y(n_188)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_111),
.Y(n_196)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_34),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_113),
.Y(n_207)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_37),
.Y(n_114)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_114),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_53),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_29),
.Y(n_116)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_29),
.Y(n_117)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_117),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_25),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_SL g154 ( 
.A1(n_118),
.A2(n_45),
.B(n_51),
.Y(n_154)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_40),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_125),
.Y(n_137)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_40),
.Y(n_120)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_53),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_2),
.Y(n_161)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_40),
.Y(n_122)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_41),
.B(n_2),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_2),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_40),
.Y(n_124)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_124),
.Y(n_197)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_41),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_126),
.B(n_168),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_42),
.B1(n_50),
.B2(n_39),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_138),
.A2(n_205),
.B1(n_148),
.B2(n_172),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_98),
.A2(n_42),
.B1(n_50),
.B2(n_39),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_139),
.A2(n_151),
.B1(n_186),
.B2(n_127),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_83),
.A2(n_38),
.B1(n_55),
.B2(n_46),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_148),
.A2(n_166),
.B1(n_172),
.B2(n_185),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_100),
.A2(n_51),
.B1(n_46),
.B2(n_34),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_71),
.B(n_2),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_152),
.B(n_199),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_154),
.A2(n_157),
.B(n_10),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_161),
.B(n_169),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_94),
.A2(n_45),
.B(n_5),
.C(n_6),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g280 ( 
.A1(n_162),
.A2(n_154),
.B(n_142),
.C(n_192),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_67),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_105),
.B(n_109),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_105),
.B(n_14),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_107),
.A2(n_112),
.B1(n_75),
.B2(n_92),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_109),
.B(n_4),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_174),
.B(n_178),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_119),
.B(n_95),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_114),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_181),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_79),
.A2(n_93),
.B1(n_86),
.B2(n_90),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_84),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_73),
.B(n_12),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_192),
.B(n_193),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_101),
.B(n_4),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_108),
.B(n_7),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_194),
.B(n_127),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_116),
.B(n_7),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_124),
.B(n_8),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_204),
.B(n_206),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_88),
.A2(n_8),
.B1(n_10),
.B2(n_89),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_69),
.B1(n_80),
.B2(n_138),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_104),
.B(n_8),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_106),
.B(n_10),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_210),
.B(n_131),
.Y(n_246)
);

INVx4_ASAP7_75t_SL g211 ( 
.A(n_142),
.Y(n_211)
);

INVx3_ASAP7_75t_SL g309 ( 
.A(n_211),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_165),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_212),
.B(n_231),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_137),
.B(n_128),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g304 ( 
.A(n_213),
.B(n_281),
.Y(n_304)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_214),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_137),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_215),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_216),
.B(n_248),
.Y(n_282)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_133),
.Y(n_218)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_218),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_156),
.B(n_80),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_219),
.B(n_224),
.Y(n_295)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_149),
.Y(n_220)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_220),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_222),
.A2(n_259),
.B1(n_277),
.B2(n_268),
.Y(n_319)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_223),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_136),
.B(n_162),
.Y(n_224)
);

INVx11_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_225),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_226),
.A2(n_221),
.B1(n_260),
.B2(n_262),
.Y(n_316)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_147),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_227),
.Y(n_328)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_147),
.Y(n_228)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_228),
.Y(n_310)
);

INVx3_ASAP7_75t_SL g229 ( 
.A(n_155),
.Y(n_229)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_229),
.Y(n_315)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_230),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_158),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_139),
.A2(n_187),
.B1(n_184),
.B2(n_203),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_232),
.A2(n_236),
.B1(n_278),
.B2(n_254),
.Y(n_294)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_184),
.A2(n_187),
.B1(n_145),
.B2(n_130),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_171),
.Y(n_237)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_237),
.Y(n_318)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_133),
.Y(n_238)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_238),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_143),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_239),
.B(n_254),
.Y(n_299)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_242),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_243),
.B(n_246),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_249),
.Y(n_284)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_163),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_245),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_146),
.B(n_159),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_247),
.B(n_255),
.Y(n_301)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_163),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_134),
.B(n_177),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_170),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_253),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_135),
.A2(n_180),
.B1(n_132),
.B2(n_183),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_252),
.A2(n_258),
.B1(n_263),
.B2(n_270),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_164),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_195),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_140),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_182),
.B(n_196),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_256),
.B(n_257),
.Y(n_300)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_170),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_135),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_173),
.A2(n_188),
.B(n_209),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_260),
.A2(n_213),
.B(n_236),
.Y(n_305)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_150),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_261),
.B(n_264),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_141),
.B(n_153),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_262),
.B(n_268),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_132),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_183),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_180),
.B(n_190),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_265),
.Y(n_311)
);

AOI21xp33_ASAP7_75t_L g267 ( 
.A1(n_200),
.A2(n_176),
.B(n_201),
.Y(n_267)
);

AOI32xp33_ASAP7_75t_L g326 ( 
.A1(n_267),
.A2(n_273),
.A3(n_211),
.B1(n_228),
.B2(n_227),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_144),
.B(n_179),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_150),
.B(n_190),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_269),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_144),
.A2(n_179),
.B1(n_201),
.B2(n_189),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_160),
.B(n_189),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_271),
.A2(n_211),
.B1(n_263),
.B2(n_244),
.Y(n_293)
);

AND2x2_ASAP7_75t_SL g272 ( 
.A(n_160),
.B(n_195),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_215),
.C(n_213),
.Y(n_288)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_191),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_273),
.B(n_274),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_208),
.B(n_202),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_208),
.B(n_202),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_276),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_129),
.B(n_155),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_129),
.A2(n_205),
.B1(n_206),
.B2(n_138),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_176),
.A2(n_151),
.B1(n_152),
.B2(n_139),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_278),
.A2(n_275),
.B1(n_276),
.B2(n_239),
.Y(n_320)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_176),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_280),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_137),
.B(n_152),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_288),
.B(n_320),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_217),
.A2(n_224),
.B1(n_226),
.B2(n_232),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_291),
.A2(n_325),
.B1(n_315),
.B2(n_309),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_293),
.B(n_326),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_219),
.A2(n_281),
.B1(n_277),
.B2(n_241),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_296),
.A2(n_297),
.B1(n_303),
.B2(n_316),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_240),
.B1(n_251),
.B2(n_234),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_251),
.A2(n_280),
.B1(n_259),
.B2(n_233),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_305),
.A2(n_327),
.B(n_312),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_247),
.B(n_237),
.C(n_242),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_304),
.C(n_303),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_319),
.A2(n_322),
.B1(n_324),
.B2(n_330),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_272),
.A2(n_235),
.B1(n_245),
.B2(n_257),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_272),
.A2(n_248),
.B1(n_250),
.B2(n_255),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_230),
.A2(n_214),
.B1(n_229),
.B2(n_258),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_326),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_220),
.A2(n_218),
.B1(n_238),
.B2(n_223),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_229),
.A2(n_261),
.B1(n_266),
.B2(n_253),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_332),
.A2(n_333),
.B1(n_309),
.B2(n_322),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_266),
.A2(n_263),
.B1(n_225),
.B2(n_264),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_279),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_335),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_336),
.A2(n_337),
.B(n_341),
.Y(n_383)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_287),
.Y(n_338)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_338),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_339),
.B(n_374),
.Y(n_377)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_287),
.Y(n_340)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_340),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_327),
.A2(n_295),
.B(n_314),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_318),
.Y(n_342)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_342),
.Y(n_385)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_318),
.Y(n_343)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_343),
.Y(n_389)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_334),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_344),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_295),
.B(n_313),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_345),
.B(n_349),
.Y(n_398)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_321),
.Y(n_346)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_346),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_313),
.B(n_306),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_347),
.B(n_348),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_306),
.B(n_296),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_331),
.B(n_307),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_321),
.Y(n_350)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_319),
.A2(n_304),
.B1(n_305),
.B2(n_301),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_352),
.A2(n_366),
.B1(n_372),
.B2(n_361),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_299),
.A2(n_311),
.B(n_282),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_353),
.A2(n_323),
.B(n_289),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_311),
.B(n_331),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_354),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_294),
.A2(n_333),
.B(n_312),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_355),
.A2(n_289),
.B(n_364),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_301),
.B(n_300),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_367),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_328),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_358),
.B(n_369),
.Y(n_382)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_362),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_288),
.A2(n_297),
.B1(n_282),
.B2(n_324),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_363),
.A2(n_364),
.B1(n_361),
.B2(n_339),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_282),
.A2(n_332),
.B1(n_304),
.B2(n_330),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_284),
.B(n_290),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_365),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_285),
.A2(n_293),
.B1(n_283),
.B2(n_286),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_286),
.B(n_292),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_317),
.B(n_298),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_368),
.B(n_375),
.Y(n_404)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_298),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_283),
.B(n_309),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_370),
.B(n_373),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_310),
.B(n_308),
.C(n_329),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_371),
.B(n_375),
.C(n_374),
.Y(n_394)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_308),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_310),
.B(n_334),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_329),
.B(n_315),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_360),
.A2(n_302),
.B(n_323),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_376),
.A2(n_380),
.B(n_386),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_336),
.A2(n_302),
.B(n_289),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_368),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_387),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_388),
.A2(n_359),
.B1(n_362),
.B2(n_372),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_341),
.B(n_352),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_390),
.B(n_404),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_361),
.A2(n_355),
.B1(n_351),
.B2(n_348),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_391),
.A2(n_392),
.B1(n_359),
.B2(n_346),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_394),
.B(n_405),
.C(n_406),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_337),
.A2(n_360),
.B(n_356),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_SL g430 ( 
.A(n_396),
.B(n_369),
.C(n_373),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_356),
.B(n_347),
.C(n_345),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_363),
.C(n_351),
.Y(n_406)
);

NOR2x1_ASAP7_75t_L g407 ( 
.A(n_337),
.B(n_357),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_353),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_382),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_410),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_398),
.B(n_367),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_411),
.B(n_433),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_403),
.Y(n_413)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_413),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_366),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_414),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_415),
.A2(n_431),
.B1(n_389),
.B2(n_397),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_377),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_416),
.B(n_421),
.Y(n_449)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_382),
.Y(n_417)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_417),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_403),
.Y(n_418)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_418),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_419),
.A2(n_420),
.B(n_385),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_408),
.A2(n_358),
.B1(n_340),
.B2(n_342),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_338),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_377),
.B(n_371),
.C(n_343),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_428),
.C(n_432),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_424),
.A2(n_387),
.B1(n_390),
.B2(n_391),
.Y(n_443)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_378),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_425),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_350),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_426),
.B(n_427),
.Y(n_437)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_379),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_377),
.B(n_406),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_380),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_408),
.A2(n_344),
.B1(n_388),
.B2(n_390),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_406),
.B(n_396),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_398),
.B(n_399),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_381),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_434),
.B(n_393),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_400),
.B(n_383),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_385),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_428),
.B(n_394),
.C(n_392),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_438),
.B(n_444),
.C(n_448),
.Y(n_466)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_439),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_426),
.B(n_384),
.Y(n_440)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_440),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_417),
.B(n_401),
.Y(n_441)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_441),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_414),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_416),
.B(n_394),
.C(n_383),
.Y(n_444)
);

XOR2x1_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_407),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_445),
.B(n_446),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_423),
.B(n_404),
.C(n_407),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_424),
.A2(n_387),
.B1(n_401),
.B2(n_395),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_459),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_453),
.A2(n_454),
.B1(n_437),
.B2(n_440),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_412),
.B(n_376),
.C(n_386),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_430),
.C(n_409),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_457),
.B(n_421),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_458),
.A2(n_429),
.B(n_409),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_409),
.A2(n_414),
.B1(n_419),
.B2(n_422),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_461),
.A2(n_479),
.B1(n_459),
.B2(n_470),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_463),
.A2(n_458),
.B(n_452),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_402),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_464),
.B(n_468),
.Y(n_485)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_454),
.Y(n_465)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_465),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_467),
.B(n_472),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_450),
.B(n_412),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_448),
.B(n_435),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_478),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_449),
.B(n_432),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_474),
.B(n_480),
.C(n_446),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_449),
.B(n_431),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_476),
.B(n_436),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_441),
.B(n_420),
.Y(n_477)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_477),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_447),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_438),
.B(n_429),
.C(n_427),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_447),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_481),
.B(n_460),
.Y(n_483)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_483),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_480),
.B(n_460),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_486),
.B(n_491),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_487),
.B(n_473),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_455),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_488),
.B(n_490),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_489),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_444),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_492),
.A2(n_495),
.B1(n_470),
.B2(n_471),
.Y(n_500)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_465),
.Y(n_495)
);

BUFx12_ASAP7_75t_L g496 ( 
.A(n_467),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_496),
.B(n_472),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_462),
.A2(n_453),
.B1(n_437),
.B2(n_451),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_497),
.A2(n_443),
.B1(n_479),
.B2(n_461),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_499),
.B(n_507),
.Y(n_512)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_500),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_485),
.B(n_462),
.Y(n_501)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_501),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_502),
.A2(n_492),
.B1(n_489),
.B2(n_471),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_436),
.C(n_476),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_504),
.B(n_505),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_491),
.B(n_474),
.C(n_461),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_490),
.B(n_473),
.C(n_463),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_506),
.B(n_487),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_482),
.A2(n_477),
.B(n_475),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_510),
.B(n_494),
.Y(n_511)
);

AOI21x1_ASAP7_75t_L g528 ( 
.A1(n_511),
.A2(n_517),
.B(n_484),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_516),
.B(n_445),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_498),
.A2(n_497),
.B(n_475),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_518),
.B(n_519),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_498),
.A2(n_484),
.B1(n_495),
.B2(n_457),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_508),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_521),
.Y(n_524)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_503),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_513),
.A2(n_509),
.B(n_505),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_523),
.A2(n_512),
.B(n_496),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_514),
.B(n_506),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_525),
.B(n_526),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_504),
.C(n_519),
.Y(n_526)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_527),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_528),
.A2(n_517),
.B(n_515),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_507),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_529),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_531),
.B(n_533),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_526),
.B(n_521),
.Y(n_533)
);

INVxp33_ASAP7_75t_L g539 ( 
.A(n_535),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_534),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_536),
.B(n_537),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_530),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g541 ( 
.A1(n_539),
.A2(n_522),
.B(n_532),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_541),
.A2(n_540),
.B(n_538),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_542),
.A2(n_524),
.B(n_529),
.Y(n_543)
);

OAI21x1_ASAP7_75t_L g544 ( 
.A1(n_543),
.A2(n_512),
.B(n_527),
.Y(n_544)
);

MAJx2_ASAP7_75t_L g545 ( 
.A(n_544),
.B(n_493),
.C(n_442),
.Y(n_545)
);


endmodule