module real_aes_18363_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_1034;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1457;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_0), .A2(n_71), .B1(n_570), .B2(n_864), .Y(n_863) );
INVxp33_ASAP7_75t_SL g902 ( .A(n_0), .Y(n_902) );
CKINVDCx5p33_ASAP7_75t_R g1006 ( .A(n_1), .Y(n_1006) );
XOR2xp5_ASAP7_75t_L g1027 ( .A(n_2), .B(n_1028), .Y(n_1027) );
CKINVDCx5p33_ASAP7_75t_R g1131 ( .A(n_3), .Y(n_1131) );
AOI221xp5_ASAP7_75t_L g988 ( .A1(n_4), .A2(n_86), .B1(n_475), .B2(n_827), .C(n_989), .Y(n_988) );
AOI22xp33_ASAP7_75t_SL g1023 ( .A1(n_4), .A2(n_137), .B1(n_583), .B2(n_861), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1497 ( .A1(n_5), .A2(n_228), .B1(n_692), .B2(n_1038), .Y(n_1497) );
AOI22xp33_ASAP7_75t_L g1508 ( .A1(n_5), .A2(n_196), .B1(n_955), .B2(n_1509), .Y(n_1508) );
INVx1_ASAP7_75t_L g737 ( .A(n_6), .Y(n_737) );
INVx1_ASAP7_75t_L g694 ( .A(n_7), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_7), .A2(n_147), .B1(n_425), .B2(n_474), .C(n_718), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g797 ( .A1(n_8), .A2(n_219), .B1(n_367), .B2(n_798), .C(n_799), .Y(n_797) );
INVx1_ASAP7_75t_L g832 ( .A(n_8), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_9), .A2(n_40), .B1(n_692), .B2(n_1038), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_9), .A2(n_223), .B1(n_538), .B2(n_1060), .Y(n_1059) );
INVx1_ASAP7_75t_L g801 ( .A(n_10), .Y(n_801) );
AOI221xp5_ASAP7_75t_L g834 ( .A1(n_10), .A2(n_152), .B1(n_770), .B2(n_835), .C(n_836), .Y(n_834) );
AOI22xp5_ASAP7_75t_SL g1240 ( .A1(n_11), .A2(n_267), .B1(n_1220), .B2(n_1227), .Y(n_1240) );
XNOR2x2_ASAP7_75t_L g1429 ( .A(n_11), .B(n_1430), .Y(n_1429) );
AOI22xp33_ASAP7_75t_L g1476 ( .A1(n_11), .A2(n_1477), .B1(n_1482), .B2(n_1519), .Y(n_1476) );
AOI21xp33_ASAP7_75t_L g756 ( .A1(n_12), .A2(n_357), .B(n_629), .Y(n_756) );
INVx1_ASAP7_75t_L g787 ( .A(n_12), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_13), .A2(n_74), .B1(n_399), .B2(n_499), .Y(n_498) );
OAI22xp33_ASAP7_75t_L g588 ( .A1(n_13), .A2(n_36), .B1(n_589), .B2(n_592), .Y(n_588) );
INVx1_ASAP7_75t_L g331 ( .A(n_14), .Y(n_331) );
OAI221xp5_ASAP7_75t_SL g451 ( .A1(n_14), .A2(n_270), .B1(n_452), .B2(n_456), .C(n_461), .Y(n_451) );
INVx1_ASAP7_75t_L g296 ( .A(n_15), .Y(n_296) );
AND2x2_ASAP7_75t_L g394 ( .A(n_15), .B(n_235), .Y(n_394) );
AND2x2_ASAP7_75t_L g419 ( .A(n_15), .B(n_420), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_15), .B(n_306), .Y(n_532) );
OAI22xp33_ASAP7_75t_L g1443 ( .A1(n_16), .A2(n_53), .B1(n_1444), .B2(n_1448), .Y(n_1443) );
INVx1_ASAP7_75t_L g1463 ( .A(n_16), .Y(n_1463) );
INVx2_ASAP7_75t_L g1215 ( .A(n_17), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_17), .B(n_1216), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_17), .B(n_109), .Y(n_1223) );
INVx1_ASAP7_75t_L g1493 ( .A(n_18), .Y(n_1493) );
OAI221xp5_ASAP7_75t_L g1513 ( .A1(n_18), .A2(n_170), .B1(n_452), .B2(n_1514), .C(n_1515), .Y(n_1513) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_19), .A2(n_237), .B1(n_560), .B2(n_564), .Y(n_676) );
INVxp67_ASAP7_75t_SL g723 ( .A(n_19), .Y(n_723) );
OAI222xp33_ASAP7_75t_L g974 ( .A1(n_20), .A2(n_153), .B1(n_456), .B2(n_975), .C1(n_976), .C2(n_980), .Y(n_974) );
INVx1_ASAP7_75t_L g1012 ( .A(n_20), .Y(n_1012) );
AOI22xp5_ASAP7_75t_SL g1250 ( .A1(n_21), .A2(n_138), .B1(n_1220), .B2(n_1227), .Y(n_1250) );
XNOR2x2_ASAP7_75t_L g792 ( .A(n_22), .B(n_793), .Y(n_792) );
OAI21xp5_ASAP7_75t_L g1065 ( .A1(n_23), .A2(n_398), .B(n_1066), .Y(n_1065) );
AOI22xp5_ASAP7_75t_SL g1260 ( .A1(n_24), .A2(n_258), .B1(n_1217), .B2(n_1222), .Y(n_1260) );
INVx1_ASAP7_75t_L g748 ( .A(n_25), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_25), .A2(n_148), .B1(n_774), .B2(n_777), .Y(n_773) );
INVx1_ASAP7_75t_L g636 ( .A(n_26), .Y(n_636) );
INVx1_ASAP7_75t_L g1063 ( .A(n_27), .Y(n_1063) );
AOI221xp5_ASAP7_75t_L g866 ( .A1(n_28), .A2(n_79), .B1(n_617), .B2(n_758), .C(n_867), .Y(n_866) );
AOI22xp33_ASAP7_75t_SL g907 ( .A1(n_28), .A2(n_31), .B1(n_776), .B2(n_777), .Y(n_907) );
CKINVDCx5p33_ASAP7_75t_R g938 ( .A(n_29), .Y(n_938) );
INVx1_ASAP7_75t_L g1046 ( .A(n_30), .Y(n_1046) );
AOI22xp33_ASAP7_75t_SL g859 ( .A1(n_31), .A2(n_136), .B1(n_570), .B2(n_680), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g1086 ( .A(n_32), .Y(n_1086) );
INVx1_ASAP7_75t_L g995 ( .A(n_33), .Y(n_995) );
AOI22xp33_ASAP7_75t_SL g1437 ( .A1(n_34), .A2(n_167), .B1(n_583), .B2(n_867), .Y(n_1437) );
INVxp67_ASAP7_75t_SL g1468 ( .A(n_34), .Y(n_1468) );
INVx1_ASAP7_75t_L g870 ( .A(n_35), .Y(n_870) );
OA222x2_ASAP7_75t_L g888 ( .A1(n_35), .A2(n_177), .B1(n_275), .B2(n_707), .C1(n_889), .C2(n_891), .Y(n_888) );
OAI211xp5_ASAP7_75t_L g486 ( .A1(n_36), .A2(n_487), .B(n_490), .C(n_533), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g1211 ( .A1(n_37), .A2(n_188), .B1(n_1212), .B2(n_1217), .Y(n_1211) );
INVx1_ASAP7_75t_L g803 ( .A(n_38), .Y(n_803) );
AOI221xp5_ASAP7_75t_L g826 ( .A1(n_38), .A2(n_77), .B1(n_827), .B2(n_829), .C(n_831), .Y(n_826) );
AOI221xp5_ASAP7_75t_L g860 ( .A1(n_39), .A2(n_222), .B1(n_629), .B2(n_861), .C(n_862), .Y(n_860) );
INVx1_ASAP7_75t_L g905 ( .A(n_39), .Y(n_905) );
AOI221xp5_ASAP7_75t_L g1051 ( .A1(n_40), .A2(n_125), .B1(n_770), .B2(n_1052), .C(n_1053), .Y(n_1051) );
OAI221xp5_ASAP7_75t_L g812 ( .A1(n_41), .A2(n_66), .B1(n_552), .B2(n_554), .C(n_556), .Y(n_812) );
INVxp67_ASAP7_75t_SL g821 ( .A(n_41), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_42), .A2(n_80), .B1(n_367), .B2(n_368), .Y(n_366) );
INVxp67_ASAP7_75t_SL g465 ( .A(n_42), .Y(n_465) );
INVxp67_ASAP7_75t_SL g981 ( .A(n_43), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_43), .A2(n_86), .B1(n_583), .B2(n_861), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1303 ( .A1(n_44), .A2(n_102), .B1(n_1220), .B2(n_1237), .Y(n_1303) );
OAI211xp5_ASAP7_75t_SL g733 ( .A1(n_45), .A2(n_734), .B(n_735), .C(n_738), .Y(n_733) );
INVx1_ASAP7_75t_L g763 ( .A(n_45), .Y(n_763) );
OAI22xp33_ASAP7_75t_L g1140 ( .A1(n_46), .A2(n_179), .B1(n_552), .B2(n_554), .Y(n_1140) );
OAI22xp5_ASAP7_75t_L g1154 ( .A1(n_46), .A2(n_83), .B1(n_664), .B2(n_666), .Y(n_1154) );
AOI22xp5_ASAP7_75t_L g1219 ( .A1(n_47), .A2(n_189), .B1(n_1220), .B2(n_1222), .Y(n_1219) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_48), .A2(n_116), .B1(n_679), .B2(n_683), .C(n_685), .Y(n_678) );
INVx1_ASAP7_75t_L g713 ( .A(n_48), .Y(n_713) );
INVx1_ASAP7_75t_L g979 ( .A(n_49), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_49), .A2(n_245), .B1(n_569), .B2(n_684), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g1040 ( .A1(n_50), .A2(n_112), .B1(n_682), .B2(n_884), .Y(n_1040) );
AOI221xp5_ASAP7_75t_L g1058 ( .A1(n_50), .A2(n_82), .B1(n_436), .B2(n_473), .C(n_896), .Y(n_1058) );
INVx1_ASAP7_75t_L g338 ( .A(n_51), .Y(n_338) );
INVx1_ASAP7_75t_L g348 ( .A(n_51), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g1228 ( .A1(n_52), .A2(n_90), .B1(n_1212), .B2(n_1220), .Y(n_1228) );
INVx1_ASAP7_75t_L g1462 ( .A(n_53), .Y(n_1462) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_54), .A2(n_100), .B1(n_691), .B2(n_692), .C(n_693), .Y(n_690) );
INVx1_ASAP7_75t_L g721 ( .A(n_54), .Y(n_721) );
CKINVDCx5p33_ASAP7_75t_R g1078 ( .A(n_55), .Y(n_1078) );
INVx1_ASAP7_75t_L g622 ( .A(n_56), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g1089 ( .A(n_57), .Y(n_1089) );
AOI22xp5_ASAP7_75t_L g1230 ( .A1(n_58), .A2(n_274), .B1(n_1212), .B2(n_1217), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_59), .A2(n_249), .B1(n_560), .B2(n_564), .Y(n_559) );
INVxp67_ASAP7_75t_SL g595 ( .A(n_59), .Y(n_595) );
INVx1_ASAP7_75t_L g289 ( .A(n_60), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_61), .A2(n_224), .B1(n_560), .B2(n_564), .Y(n_811) );
INVx1_ASAP7_75t_L g825 ( .A(n_61), .Y(n_825) );
INVx2_ASAP7_75t_L g328 ( .A(n_62), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_63), .A2(n_245), .B1(n_538), .B2(n_991), .Y(n_990) );
AOI22xp5_ASAP7_75t_L g1020 ( .A1(n_63), .A2(n_159), .B1(n_684), .B2(n_1021), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_64), .A2(n_229), .B1(n_798), .B2(n_862), .Y(n_1170) );
AOI221xp5_ASAP7_75t_L g1190 ( .A1(n_64), .A2(n_173), .B1(n_1191), .B2(n_1194), .C(n_1195), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_65), .A2(n_201), .B1(n_589), .B2(n_592), .Y(n_796) );
INVx1_ASAP7_75t_L g823 ( .A(n_65), .Y(n_823) );
INVx1_ASAP7_75t_L g845 ( .A(n_66), .Y(n_845) );
INVx1_ASAP7_75t_L g1129 ( .A(n_67), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g1150 ( .A1(n_67), .A2(n_233), .B1(n_538), .B2(n_776), .Y(n_1150) );
AOI22xp5_ASAP7_75t_L g1261 ( .A1(n_68), .A2(n_73), .B1(n_1212), .B2(n_1220), .Y(n_1261) );
CKINVDCx5p33_ASAP7_75t_R g1139 ( .A(n_69), .Y(n_1139) );
AOI21xp33_ASAP7_75t_L g627 ( .A1(n_70), .A2(n_628), .B(n_629), .Y(n_627) );
INVxp67_ASAP7_75t_L g650 ( .A(n_70), .Y(n_650) );
INVxp67_ASAP7_75t_SL g906 ( .A(n_71), .Y(n_906) );
INVx1_ASAP7_75t_L g1094 ( .A(n_72), .Y(n_1094) );
OAI221xp5_ASAP7_75t_L g551 ( .A1(n_74), .A2(n_124), .B1(n_552), .B2(n_554), .C(n_556), .Y(n_551) );
AOI22xp33_ASAP7_75t_SL g1174 ( .A1(n_75), .A2(n_117), .B1(n_342), .B2(n_1169), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_75), .A2(n_145), .B1(n_439), .B2(n_441), .Y(n_1196) );
INVx1_ASAP7_75t_L g696 ( .A(n_76), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g804 ( .A1(n_77), .A2(n_220), .B1(n_798), .B2(n_805), .C(n_806), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_78), .A2(n_253), .B1(n_357), .B2(n_372), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_78), .A2(n_226), .B1(n_439), .B2(n_441), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g895 ( .A1(n_79), .A2(n_222), .B1(n_896), .B2(n_898), .C(n_899), .Y(n_895) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_80), .A2(n_99), .B1(n_423), .B2(n_429), .C(n_436), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g1159 ( .A(n_81), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_82), .A2(n_234), .B1(n_1035), .B2(n_1036), .Y(n_1034) );
OAI221xp5_ASAP7_75t_L g1136 ( .A1(n_83), .A2(n_178), .B1(n_755), .B2(n_1137), .C(n_1138), .Y(n_1136) );
INVx1_ASAP7_75t_L g882 ( .A(n_84), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g886 ( .A(n_84), .B(n_487), .Y(n_886) );
OAI222xp33_ASAP7_75t_L g1100 ( .A1(n_85), .A2(n_130), .B1(n_246), .B2(n_563), .C1(n_695), .C2(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g1114 ( .A(n_85), .Y(n_1114) );
AOI22xp5_ASAP7_75t_L g1226 ( .A1(n_87), .A2(n_200), .B1(n_1217), .B2(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g760 ( .A(n_88), .Y(n_760) );
CKINVDCx5p33_ASAP7_75t_R g1180 ( .A(n_89), .Y(n_1180) );
INVx1_ASAP7_75t_L g525 ( .A(n_91), .Y(n_525) );
AOI221xp5_ASAP7_75t_L g749 ( .A1(n_92), .A2(n_140), .B1(n_617), .B2(n_750), .C(n_751), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_92), .A2(n_208), .B1(n_416), .B2(n_774), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g1164 ( .A(n_93), .Y(n_1164) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_94), .A2(n_192), .B1(n_589), .B2(n_592), .Y(n_637) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_94), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g1452 ( .A1(n_95), .A2(n_134), .B1(n_398), .B2(n_917), .Y(n_1452) );
INVx1_ASAP7_75t_L g883 ( .A(n_96), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_96), .A2(n_197), .B1(n_399), .B2(n_499), .Y(n_908) );
INVx1_ASAP7_75t_L g1088 ( .A(n_97), .Y(n_1088) );
AOI221xp5_ASAP7_75t_L g1105 ( .A1(n_97), .A2(n_154), .B1(n_751), .B2(n_798), .C(n_1106), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g1495 ( .A1(n_98), .A2(n_122), .B1(n_583), .B2(n_884), .Y(n_1495) );
AOI221xp5_ASAP7_75t_L g1505 ( .A1(n_98), .A2(n_280), .B1(n_898), .B2(n_1506), .C(n_1507), .Y(n_1505) );
AOI22xp33_ASAP7_75t_SL g383 ( .A1(n_99), .A2(n_172), .B1(n_342), .B2(n_384), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_100), .A2(n_203), .B1(n_425), .B2(n_474), .C(n_712), .Y(n_711) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_101), .Y(n_291) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_101), .B(n_289), .Y(n_1213) );
CKINVDCx5p33_ASAP7_75t_R g941 ( .A(n_103), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_104), .A2(n_168), .B1(n_372), .B2(n_758), .Y(n_933) );
AOI22xp5_ASAP7_75t_L g960 ( .A1(n_104), .A2(n_106), .B1(n_774), .B2(n_777), .Y(n_960) );
INVx1_ASAP7_75t_L g599 ( .A(n_105), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g1235 ( .A1(n_105), .A2(n_171), .B1(n_1212), .B2(n_1217), .Y(n_1235) );
INVx1_ASAP7_75t_L g943 ( .A(n_106), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g1441 ( .A1(n_107), .A2(n_132), .B1(n_684), .B2(n_1439), .Y(n_1441) );
AOI221xp5_ASAP7_75t_L g1471 ( .A1(n_107), .A2(n_181), .B1(n_835), .B2(n_1472), .C(n_1474), .Y(n_1471) );
INVx1_ASAP7_75t_L g355 ( .A(n_108), .Y(n_355) );
INVx1_ASAP7_75t_L g1216 ( .A(n_109), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_109), .B(n_1215), .Y(n_1221) );
AOI22xp5_ASAP7_75t_L g1241 ( .A1(n_110), .A2(n_198), .B1(n_1212), .B2(n_1217), .Y(n_1241) );
AOI22xp5_ASAP7_75t_L g911 ( .A1(n_111), .A2(n_912), .B1(n_913), .B2(n_967), .Y(n_911) );
INVx1_ASAP7_75t_L g967 ( .A(n_111), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_112), .A2(n_234), .B1(n_777), .B2(n_991), .Y(n_1054) );
OAI22xp33_ASAP7_75t_L g689 ( .A1(n_113), .A2(n_163), .B1(n_589), .B2(n_592), .Y(n_689) );
INVxp67_ASAP7_75t_SL g725 ( .A(n_113), .Y(n_725) );
AOI22xp33_ASAP7_75t_SL g1166 ( .A1(n_114), .A2(n_145), .B1(n_1167), .B2(n_1169), .Y(n_1166) );
AOI221xp5_ASAP7_75t_L g1183 ( .A1(n_114), .A2(n_117), .B1(n_436), .B2(n_1184), .C(n_1187), .Y(n_1183) );
CKINVDCx5p33_ASAP7_75t_R g1160 ( .A(n_115), .Y(n_1160) );
INVx1_ASAP7_75t_L g719 ( .A(n_116), .Y(n_719) );
INVx2_ASAP7_75t_L g330 ( .A(n_118), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_118), .B(n_328), .Y(n_354) );
INVx1_ASAP7_75t_L g382 ( .A(n_118), .Y(n_382) );
INVx1_ASAP7_75t_L g624 ( .A(n_119), .Y(n_624) );
INVx1_ASAP7_75t_L g1095 ( .A(n_120), .Y(n_1095) );
OAI22xp33_ASAP7_75t_L g1103 ( .A1(n_120), .A2(n_166), .B1(n_552), .B2(n_554), .Y(n_1103) );
CKINVDCx5p33_ASAP7_75t_R g1124 ( .A(n_121), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1518 ( .A1(n_122), .A2(n_269), .B1(n_991), .B2(n_1509), .Y(n_1518) );
INVxp67_ASAP7_75t_SL g754 ( .A(n_123), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_123), .A2(n_140), .B1(n_768), .B2(n_771), .Y(n_767) );
INVxp67_ASAP7_75t_SL g540 ( .A(n_124), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_125), .A2(n_223), .B1(n_692), .B2(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_L g1435 ( .A(n_126), .Y(n_1435) );
OAI221xp5_ASAP7_75t_L g1464 ( .A1(n_126), .A2(n_205), .B1(n_1465), .B2(n_1466), .C(n_1467), .Y(n_1464) );
OAI22xp5_ASAP7_75t_L g1488 ( .A1(n_127), .A2(n_157), .B1(n_917), .B2(n_997), .Y(n_1488) );
AOI221xp5_ASAP7_75t_L g526 ( .A1(n_128), .A2(n_149), .B1(n_515), .B2(n_527), .C(n_529), .Y(n_526) );
AOI221xp5_ASAP7_75t_L g582 ( .A1(n_128), .A2(n_162), .B1(n_570), .B2(n_583), .C(n_584), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g1496 ( .A1(n_129), .A2(n_196), .B1(n_378), .B2(n_1038), .Y(n_1496) );
AOI21xp33_ASAP7_75t_L g1517 ( .A1(n_129), .A2(n_1053), .B(n_1506), .Y(n_1517) );
OAI221xp5_ASAP7_75t_L g1091 ( .A1(n_130), .A2(n_166), .B1(n_492), .B2(n_664), .C(n_666), .Y(n_1091) );
INVx1_ASAP7_75t_L g1069 ( .A(n_131), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1456 ( .A1(n_132), .A2(n_183), .B1(n_956), .B2(n_1457), .Y(n_1456) );
INVx1_ASAP7_75t_L g523 ( .A(n_133), .Y(n_523) );
AOI221xp5_ASAP7_75t_L g567 ( .A1(n_133), .A2(n_279), .B1(n_568), .B2(n_570), .C(n_571), .Y(n_567) );
OAI211xp5_ASAP7_75t_L g1454 ( .A1(n_134), .A2(n_414), .B(n_1455), .C(n_1461), .Y(n_1454) );
OAI221xp5_ASAP7_75t_L g675 ( .A1(n_135), .A2(n_207), .B1(n_552), .B2(n_554), .C(n_556), .Y(n_675) );
OAI21xp33_ASAP7_75t_L g706 ( .A1(n_135), .A2(n_492), .B(n_707), .Y(n_706) );
INVxp67_ASAP7_75t_SL g900 ( .A(n_136), .Y(n_900) );
INVxp67_ASAP7_75t_SL g983 ( .A(n_137), .Y(n_983) );
INVx1_ASAP7_75t_L g810 ( .A(n_139), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_141), .A2(n_731), .B1(n_790), .B2(n_791), .Y(n_730) );
INVx1_ASAP7_75t_L g791 ( .A(n_141), .Y(n_791) );
OAI211xp5_ASAP7_75t_SL g986 ( .A1(n_142), .A2(n_414), .B(n_987), .C(n_992), .Y(n_986) );
INVx1_ASAP7_75t_L g1015 ( .A(n_142), .Y(n_1015) );
CKINVDCx5p33_ASAP7_75t_R g1487 ( .A(n_143), .Y(n_1487) );
XOR2x2_ASAP7_75t_L g606 ( .A(n_144), .B(n_607), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g1126 ( .A1(n_146), .A2(n_564), .B1(n_1127), .B2(n_1130), .Y(n_1126) );
INVx1_ASAP7_75t_L g1145 ( .A(n_146), .Y(n_1145) );
INVx1_ASAP7_75t_L g686 ( .A(n_147), .Y(n_686) );
AOI22xp33_ASAP7_75t_SL g757 ( .A1(n_148), .A2(n_208), .B1(n_684), .B2(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g575 ( .A(n_149), .Y(n_575) );
INVx1_ASAP7_75t_L g739 ( .A(n_150), .Y(n_739) );
OAI221xp5_ASAP7_75t_L g765 ( .A1(n_150), .A2(n_206), .B1(n_666), .B2(n_709), .C(n_766), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g1031 ( .A(n_151), .Y(n_1031) );
INVx1_ASAP7_75t_L g807 ( .A(n_152), .Y(n_807) );
INVx1_ASAP7_75t_L g1009 ( .A(n_153), .Y(n_1009) );
INVx1_ASAP7_75t_L g1075 ( .A(n_154), .Y(n_1075) );
CKINVDCx5p33_ASAP7_75t_R g1179 ( .A(n_155), .Y(n_1179) );
AOI22xp5_ASAP7_75t_L g1236 ( .A1(n_156), .A2(n_194), .B1(n_1220), .B2(n_1237), .Y(n_1236) );
OAI211xp5_ASAP7_75t_L g1502 ( .A1(n_157), .A2(n_1503), .B(n_1504), .C(n_1510), .Y(n_1502) );
BUFx3_ASAP7_75t_L g322 ( .A(n_158), .Y(n_322) );
INVx1_ASAP7_75t_L g978 ( .A(n_159), .Y(n_978) );
INVx1_ASAP7_75t_L g740 ( .A(n_160), .Y(n_740) );
INVx1_ASAP7_75t_L g674 ( .A(n_161), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g511 ( .A1(n_162), .A2(n_217), .B1(n_512), .B2(n_515), .C(n_518), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_163), .A2(n_207), .B1(n_666), .B2(n_709), .Y(n_708) );
XNOR2x1_ASAP7_75t_L g970 ( .A(n_164), .B(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g610 ( .A(n_165), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g1458 ( .A1(n_167), .A2(n_247), .B1(n_473), .B2(n_989), .C(n_1459), .Y(n_1458) );
AOI22xp33_ASAP7_75t_SL g954 ( .A1(n_168), .A2(n_242), .B1(n_955), .B2(n_956), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_169), .A2(n_173), .B1(n_357), .B2(n_1172), .Y(n_1171) );
AOI22xp33_ASAP7_75t_SL g1188 ( .A1(n_169), .A2(n_229), .B1(n_439), .B2(n_441), .Y(n_1188) );
INVx1_ASAP7_75t_L g1492 ( .A(n_170), .Y(n_1492) );
INVxp67_ASAP7_75t_SL g471 ( .A(n_172), .Y(n_471) );
OAI21xp5_ASAP7_75t_SL g1199 ( .A1(n_174), .A2(n_398), .B(n_1200), .Y(n_1199) );
AOI22xp5_ASAP7_75t_L g1231 ( .A1(n_175), .A2(n_227), .B1(n_1220), .B2(n_1227), .Y(n_1231) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_176), .Y(n_303) );
INVx1_ASAP7_75t_L g885 ( .A(n_177), .Y(n_885) );
OAI211xp5_ASAP7_75t_L g1143 ( .A1(n_178), .A2(n_817), .B(n_1144), .C(n_1147), .Y(n_1143) );
INVx1_ASAP7_75t_L g1146 ( .A(n_179), .Y(n_1146) );
CKINVDCx5p33_ASAP7_75t_R g1123 ( .A(n_180), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1438 ( .A1(n_181), .A2(n_183), .B1(n_692), .B2(n_1439), .Y(n_1438) );
INVx1_ASAP7_75t_L g1062 ( .A(n_182), .Y(n_1062) );
OAI222xp33_ASAP7_75t_L g386 ( .A1(n_184), .A2(n_225), .B1(n_243), .B2(n_387), .C1(n_398), .C2(n_408), .Y(n_386) );
OAI211xp5_ASAP7_75t_L g413 ( .A1(n_184), .A2(n_414), .B(n_421), .C(n_444), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_185), .A2(n_583), .B(n_617), .Y(n_616) );
INVxp67_ASAP7_75t_SL g647 ( .A(n_185), .Y(n_647) );
OAI21xp5_ASAP7_75t_L g996 ( .A1(n_186), .A2(n_997), .B(n_998), .Y(n_996) );
INVx1_ASAP7_75t_L g1044 ( .A(n_187), .Y(n_1044) );
INVx1_ASAP7_75t_L g928 ( .A(n_190), .Y(n_928) );
OAI221xp5_ASAP7_75t_L g957 ( .A1(n_190), .A2(n_707), .B1(n_958), .B2(n_961), .C(n_962), .Y(n_957) );
CKINVDCx5p33_ASAP7_75t_R g1085 ( .A(n_191), .Y(n_1085) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_192), .A2(n_221), .B1(n_492), .B2(n_664), .C(n_666), .Y(n_663) );
INVx1_ASAP7_75t_L g1133 ( .A(n_193), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_193), .A2(n_204), .B1(n_416), .B2(n_776), .Y(n_1153) );
CKINVDCx5p33_ASAP7_75t_R g1451 ( .A(n_195), .Y(n_1451) );
INVx1_ASAP7_75t_L g869 ( .A(n_197), .Y(n_869) );
OAI22xp33_ASAP7_75t_L g1499 ( .A1(n_199), .A2(n_259), .B1(n_1444), .B2(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1511 ( .A(n_199), .Y(n_1511) );
INVxp67_ASAP7_75t_SL g843 ( .A(n_201), .Y(n_843) );
INVx1_ASAP7_75t_L g635 ( .A(n_202), .Y(n_635) );
INVx1_ASAP7_75t_L g688 ( .A(n_203), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g1121 ( .A1(n_204), .A2(n_233), .B1(n_632), .B2(n_684), .C(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1434 ( .A(n_205), .Y(n_1434) );
INVx1_ASAP7_75t_L g761 ( .A(n_206), .Y(n_761) );
CKINVDCx5p33_ASAP7_75t_R g919 ( .A(n_209), .Y(n_919) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_210), .Y(n_302) );
INVx1_ASAP7_75t_L g619 ( .A(n_211), .Y(n_619) );
XNOR2x1_ASAP7_75t_L g670 ( .A(n_212), .B(n_671), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g1163 ( .A(n_213), .Y(n_1163) );
CKINVDCx5p33_ASAP7_75t_R g1128 ( .A(n_214), .Y(n_1128) );
CKINVDCx5p33_ASAP7_75t_R g1081 ( .A(n_215), .Y(n_1081) );
INVxp67_ASAP7_75t_SL g1093 ( .A(n_216), .Y(n_1093) );
OAI22xp5_ASAP7_75t_L g1108 ( .A1(n_216), .A2(n_564), .B1(n_1109), .B2(n_1111), .Y(n_1108) );
INVx1_ASAP7_75t_L g572 ( .A(n_217), .Y(n_572) );
INVx1_ASAP7_75t_L g534 ( .A(n_218), .Y(n_534) );
INVx1_ASAP7_75t_L g837 ( .A(n_219), .Y(n_837) );
INVx1_ASAP7_75t_L g840 ( .A(n_220), .Y(n_840) );
OAI221xp5_ASAP7_75t_L g611 ( .A1(n_221), .A2(n_239), .B1(n_552), .B2(n_554), .C(n_556), .Y(n_611) );
INVxp67_ASAP7_75t_SL g815 ( .A(n_224), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_226), .A2(n_250), .B1(n_376), .B2(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g1516 ( .A(n_228), .Y(n_1516) );
INVx1_ASAP7_75t_L g915 ( .A(n_230), .Y(n_915) );
INVxp67_ASAP7_75t_SL g920 ( .A(n_231), .Y(n_920) );
OAI221xp5_ASAP7_75t_L g934 ( .A1(n_231), .A2(n_556), .B1(n_560), .B2(n_935), .C(n_940), .Y(n_934) );
CKINVDCx5p33_ASAP7_75t_R g1076 ( .A(n_232), .Y(n_1076) );
BUFx3_ASAP7_75t_L g306 ( .A(n_235), .Y(n_306) );
INVx1_ASAP7_75t_L g420 ( .A(n_235), .Y(n_420) );
INVx1_ASAP7_75t_L g909 ( .A(n_236), .Y(n_909) );
INVxp67_ASAP7_75t_SL g701 ( .A(n_237), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g932 ( .A1(n_238), .A2(n_376), .B(n_629), .Y(n_932) );
INVx1_ASAP7_75t_L g953 ( .A(n_238), .Y(n_953) );
INVxp67_ASAP7_75t_SL g668 ( .A(n_239), .Y(n_668) );
XOR2xp5_ASAP7_75t_L g1156 ( .A(n_240), .B(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g736 ( .A(n_241), .Y(n_736) );
INVx1_ASAP7_75t_L g939 ( .A(n_242), .Y(n_939) );
CKINVDCx5p33_ASAP7_75t_R g925 ( .A(n_244), .Y(n_925) );
INVx1_ASAP7_75t_L g1097 ( .A(n_246), .Y(n_1097) );
AOI22xp33_ASAP7_75t_SL g1442 ( .A1(n_247), .A2(n_265), .B1(n_583), .B2(n_861), .Y(n_1442) );
INVx1_ASAP7_75t_L g325 ( .A(n_248), .Y(n_325) );
INVx1_ASAP7_75t_L g353 ( .A(n_248), .Y(n_353) );
INVx2_ASAP7_75t_L g365 ( .A(n_248), .Y(n_365) );
INVxp67_ASAP7_75t_SL g544 ( .A(n_249), .Y(n_544) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_250), .A2(n_253), .B1(n_473), .B2(n_474), .C(n_476), .Y(n_472) );
XNOR2xp5_ASAP7_75t_L g1483 ( .A(n_251), .B(n_1484), .Y(n_1483) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_252), .A2(n_263), .B1(n_374), .B2(n_632), .Y(n_631) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_252), .Y(n_660) );
INVx1_ASAP7_75t_L g808 ( .A(n_254), .Y(n_808) );
INVx1_ASAP7_75t_L g1030 ( .A(n_255), .Y(n_1030) );
INVx1_ASAP7_75t_L g340 ( .A(n_256), .Y(n_340) );
INVx1_ASAP7_75t_L g1117 ( .A(n_257), .Y(n_1117) );
AOI22xp5_ASAP7_75t_L g1249 ( .A1(n_257), .A2(n_272), .B1(n_1212), .B2(n_1217), .Y(n_1249) );
INVx1_ASAP7_75t_L g1512 ( .A(n_259), .Y(n_1512) );
INVx1_ASAP7_75t_L g1135 ( .A(n_260), .Y(n_1135) );
CKINVDCx5p33_ASAP7_75t_R g930 ( .A(n_261), .Y(n_930) );
INVx1_ASAP7_75t_L g614 ( .A(n_262), .Y(n_614) );
INVxp67_ASAP7_75t_SL g646 ( .A(n_263), .Y(n_646) );
INVx1_ASAP7_75t_L g1301 ( .A(n_264), .Y(n_1301) );
INVxp67_ASAP7_75t_SL g1470 ( .A(n_265), .Y(n_1470) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_266), .B(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g745 ( .A(n_268), .Y(n_745) );
AOI22xp33_ASAP7_75t_SL g1498 ( .A1(n_269), .A2(n_280), .B1(n_583), .B2(n_884), .Y(n_1498) );
INVx1_ASAP7_75t_L g317 ( .A(n_270), .Y(n_317) );
XNOR2xp5_ASAP7_75t_L g312 ( .A(n_271), .B(n_313), .Y(n_312) );
NAND2xp33_ASAP7_75t_SL g507 ( .A(n_273), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g585 ( .A(n_273), .Y(n_585) );
OAI221xp5_ASAP7_75t_L g875 ( .A1(n_275), .A2(n_278), .B1(n_876), .B2(n_877), .C(n_881), .Y(n_875) );
INVx1_ASAP7_75t_L g927 ( .A(n_276), .Y(n_927) );
INVx1_ASAP7_75t_L g994 ( .A(n_277), .Y(n_994) );
INVxp67_ASAP7_75t_SL g893 ( .A(n_278), .Y(n_893) );
INVx1_ASAP7_75t_L g504 ( .A(n_279), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_307), .B(n_1203), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx4f_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_292), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g1427 ( .A(n_286), .B(n_295), .Y(n_1427) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g1481 ( .A(n_288), .B(n_291), .Y(n_1481) );
INVx1_ASAP7_75t_L g1521 ( .A(n_288), .Y(n_1521) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g1523 ( .A(n_291), .B(n_1521), .Y(n_1523) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g437 ( .A(n_296), .B(n_306), .Y(n_437) );
AND2x4_ASAP7_75t_L g477 ( .A(n_296), .B(n_305), .Y(n_477) );
AND2x4_ASAP7_75t_SL g1426 ( .A(n_297), .B(n_1427), .Y(n_1426) );
INVx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x6_ASAP7_75t_L g298 ( .A(n_299), .B(n_304), .Y(n_298) );
INVxp67_ASAP7_75t_L g715 ( .A(n_299), .Y(n_715) );
BUFx4f_ASAP7_75t_L g720 ( .A(n_299), .Y(n_720) );
INVx1_ASAP7_75t_L g839 ( .A(n_299), .Y(n_839) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx4f_ASAP7_75t_L g464 ( .A(n_300), .Y(n_464) );
INVx3_ASAP7_75t_L g517 ( .A(n_300), .Y(n_517) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g396 ( .A(n_302), .Y(n_396) );
INVx1_ASAP7_75t_L g402 ( .A(n_302), .Y(n_402) );
INVx2_ASAP7_75t_L g418 ( .A(n_302), .Y(n_418) );
AND2x2_ASAP7_75t_L g428 ( .A(n_302), .B(n_303), .Y(n_428) );
AND2x2_ASAP7_75t_L g434 ( .A(n_302), .B(n_435), .Y(n_434) );
NAND2x1_ASAP7_75t_L g494 ( .A(n_302), .B(n_303), .Y(n_494) );
INVx1_ASAP7_75t_L g397 ( .A(n_303), .Y(n_397) );
AND2x2_ASAP7_75t_L g417 ( .A(n_303), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g435 ( .A(n_303), .Y(n_435) );
BUFx2_ASAP7_75t_L g459 ( .A(n_303), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_303), .B(n_418), .Y(n_470) );
OR2x2_ASAP7_75t_L g510 ( .A(n_303), .B(n_396), .Y(n_510) );
INVxp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI22xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_850), .B1(n_1201), .B2(n_1202), .Y(n_307) );
INVxp67_ASAP7_75t_SL g1201 ( .A(n_308), .Y(n_1201) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_603), .B1(n_848), .B2(n_849), .Y(n_308) );
INVxp67_ASAP7_75t_SL g848 ( .A(n_309), .Y(n_848) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_482), .B1(n_600), .B2(n_601), .Y(n_309) );
INVx1_ASAP7_75t_L g600 ( .A(n_310), .Y(n_600) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_412), .Y(n_313) );
NOR3xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_386), .C(n_411), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_339), .C(n_360), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B1(n_331), .B2(n_332), .Y(n_316) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_323), .Y(n_318) );
AND2x6_ASAP7_75t_L g553 ( .A(n_319), .B(n_326), .Y(n_553) );
NAND2x1_ASAP7_75t_L g1011 ( .A(n_319), .B(n_323), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_319), .B(n_323), .Y(n_1045) );
INVx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g374 ( .A(n_321), .B(n_336), .Y(n_374) );
NAND2x1p5_ASAP7_75t_L g406 ( .A(n_321), .B(n_407), .Y(n_406) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g345 ( .A(n_322), .Y(n_345) );
AND2x4_ASAP7_75t_L g370 ( .A(n_322), .B(n_337), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_322), .B(n_338), .Y(n_391) );
OR2x2_ASAP7_75t_L g579 ( .A(n_322), .B(n_347), .Y(n_579) );
AND2x4_ASAP7_75t_L g332 ( .A(n_323), .B(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g411 ( .A(n_323), .B(n_385), .Y(n_411) );
AND2x4_ASAP7_75t_SL g1013 ( .A(n_323), .B(n_333), .Y(n_1013) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
OR2x2_ASAP7_75t_L g392 ( .A(n_324), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g546 ( .A(n_324), .Y(n_546) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g381 ( .A(n_325), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_325), .B(n_419), .Y(n_537) );
NAND2x1p5_ASAP7_75t_L g409 ( .A(n_326), .B(n_344), .Y(n_409) );
AND2x2_ASAP7_75t_L g555 ( .A(n_326), .B(n_335), .Y(n_555) );
INVx1_ASAP7_75t_L g558 ( .A(n_326), .Y(n_558) );
AND2x4_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
NAND3x1_ASAP7_75t_L g380 ( .A(n_327), .B(n_381), .C(n_382), .Y(n_380) );
NAND2x1p5_ASAP7_75t_L g581 ( .A(n_327), .B(n_382), .Y(n_581) );
INVx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx3_ASAP7_75t_L g363 ( .A(n_328), .Y(n_363) );
NAND2xp33_ASAP7_75t_SL g630 ( .A(n_328), .B(n_330), .Y(n_630) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND3x4_ASAP7_75t_L g362 ( .A(n_330), .B(n_363), .C(n_364), .Y(n_362) );
AND2x2_ASAP7_75t_L g587 ( .A(n_330), .B(n_363), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_332), .A2(n_1044), .B1(n_1045), .B2(n_1046), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_332), .A2(n_1010), .B1(n_1163), .B2(n_1164), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g1433 ( .A1(n_332), .A2(n_1010), .B1(n_1434), .B2(n_1435), .Y(n_1433) );
AOI22xp33_ASAP7_75t_L g1491 ( .A1(n_332), .A2(n_1045), .B1(n_1492), .B2(n_1493), .Y(n_1491) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g407 ( .A(n_338), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_355), .B2(n_356), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_340), .A2(n_355), .B1(n_445), .B2(n_448), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_341), .A2(n_356), .B1(n_1179), .B2(n_1180), .Y(n_1200) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_349), .Y(n_341) );
AND2x4_ASAP7_75t_L g999 ( .A(n_342), .B(n_349), .Y(n_999) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g367 ( .A(n_343), .Y(n_367) );
INVx8_ASAP7_75t_L g583 ( .A(n_343), .Y(n_583) );
INVx8_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g590 ( .A(n_344), .B(n_591), .Y(n_590) );
BUFx3_ASAP7_75t_L g632 ( .A(n_344), .Y(n_632) );
BUFx3_ASAP7_75t_L g682 ( .A(n_344), .Y(n_682) );
HB1xp67_ASAP7_75t_L g1035 ( .A(n_344), .Y(n_1035) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
AND2x4_ASAP7_75t_L g358 ( .A(n_345), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVxp67_ASAP7_75t_L g359 ( .A(n_348), .Y(n_359) );
AND2x4_ASAP7_75t_L g356 ( .A(n_349), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g388 ( .A(n_350), .B(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g404 ( .A(n_350), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g1002 ( .A(n_350), .Y(n_1002) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_354), .Y(n_350) );
INVx1_ASAP7_75t_L g520 ( .A(n_351), .Y(n_520) );
AND2x2_ASAP7_75t_SL g662 ( .A(n_351), .B(n_437), .Y(n_662) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx2_ASAP7_75t_L g403 ( .A(n_352), .Y(n_403) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g562 ( .A(n_354), .Y(n_562) );
INVx1_ASAP7_75t_L g591 ( .A(n_354), .Y(n_591) );
INVx2_ASAP7_75t_L g1448 ( .A(n_356), .Y(n_1448) );
INVx2_ASAP7_75t_L g1500 ( .A(n_356), .Y(n_1500) );
INVx3_ASAP7_75t_L g377 ( .A(n_357), .Y(n_377) );
INVx2_ASAP7_75t_SL g586 ( .A(n_357), .Y(n_586) );
INVx2_ASAP7_75t_SL g687 ( .A(n_357), .Y(n_687) );
INVx3_ASAP7_75t_L g1022 ( .A(n_357), .Y(n_1022) );
BUFx8_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g563 ( .A(n_358), .Y(n_563) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_358), .Y(n_569) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_358), .Y(n_628) );
AOI33xp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_366), .A3(n_371), .B1(n_375), .B2(n_379), .B3(n_383), .Y(n_360) );
AOI33xp33_ASAP7_75t_L g1165 ( .A1(n_361), .A2(n_1166), .A3(n_1170), .B1(n_1171), .B2(n_1173), .B3(n_1174), .Y(n_1165) );
BUFx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AOI33xp33_ASAP7_75t_L g1017 ( .A1(n_362), .A2(n_1018), .A3(n_1019), .B1(n_1020), .B2(n_1023), .B3(n_1024), .Y(n_1017) );
AOI33xp33_ASAP7_75t_L g1033 ( .A1(n_362), .A2(n_1034), .A3(n_1037), .B1(n_1039), .B2(n_1040), .B3(n_1041), .Y(n_1033) );
AOI33xp33_ASAP7_75t_L g1436 ( .A1(n_362), .A2(n_1024), .A3(n_1437), .B1(n_1438), .B2(n_1441), .B3(n_1442), .Y(n_1436) );
AOI33xp33_ASAP7_75t_L g1494 ( .A1(n_362), .A2(n_1041), .A3(n_1495), .B1(n_1496), .B2(n_1497), .B3(n_1498), .Y(n_1494) );
INVx1_ASAP7_75t_L g481 ( .A(n_364), .Y(n_481) );
INVx2_ASAP7_75t_SL g1475 ( .A(n_364), .Y(n_1475) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_365), .B(n_394), .Y(n_497) );
BUFx2_ASAP7_75t_L g531 ( .A(n_365), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_367), .A2(n_882), .B1(n_883), .B2(n_884), .Y(n_881) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g1036 ( .A(n_369), .Y(n_1036) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g385 ( .A(n_370), .Y(n_385) );
AND2x2_ASAP7_75t_L g593 ( .A(n_370), .B(n_591), .Y(n_593) );
BUFx2_ASAP7_75t_L g750 ( .A(n_370), .Y(n_750) );
BUFx2_ASAP7_75t_L g861 ( .A(n_370), .Y(n_861) );
BUFx3_ASAP7_75t_L g867 ( .A(n_370), .Y(n_867) );
BUFx2_ASAP7_75t_L g884 ( .A(n_370), .Y(n_884) );
BUFx2_ASAP7_75t_L g1169 ( .A(n_370), .Y(n_1169) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g378 ( .A(n_373), .Y(n_378) );
INVx2_ASAP7_75t_R g692 ( .A(n_373), .Y(n_692) );
INVx5_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g565 ( .A(n_374), .B(n_562), .Y(n_565) );
BUFx2_ASAP7_75t_L g570 ( .A(n_374), .Y(n_570) );
BUFx12f_ASAP7_75t_L g684 ( .A(n_374), .Y(n_684) );
BUFx3_ASAP7_75t_L g798 ( .A(n_374), .Y(n_798) );
BUFx3_ASAP7_75t_L g1172 ( .A(n_374), .Y(n_1172) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g1111 ( .A1(n_377), .A2(n_1078), .B1(n_1089), .B2(n_1112), .Y(n_1111) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx3_ASAP7_75t_L g1025 ( .A(n_380), .Y(n_1025) );
BUFx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx8_ASAP7_75t_L g1005 ( .A(n_387), .Y(n_1005) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_392), .Y(n_387) );
INVx1_ASAP7_75t_L g621 ( .A(n_389), .Y(n_621) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_390), .Y(n_747) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx2_ASAP7_75t_L g880 ( .A(n_391), .Y(n_880) );
INVx1_ASAP7_75t_L g890 ( .A(n_392), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_392), .B(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g547 ( .A(n_393), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_394), .B(n_401), .Y(n_400) );
AND2x6_ASAP7_75t_L g442 ( .A(n_394), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g460 ( .A(n_394), .Y(n_460) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_394), .B(n_1056), .Y(n_1055) );
INVx3_ASAP7_75t_L g440 ( .A(n_395), .Y(n_440) );
AND2x2_ASAP7_75t_L g447 ( .A(n_395), .B(n_419), .Y(n_447) );
BUFx6f_ASAP7_75t_L g776 ( .A(n_395), .Y(n_776) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
AND2x4_ASAP7_75t_L g398 ( .A(n_399), .B(n_404), .Y(n_398) );
INVx2_ASAP7_75t_SL g822 ( .A(n_399), .Y(n_822) );
AND2x4_ASAP7_75t_L g997 ( .A(n_399), .B(n_404), .Y(n_997) );
OR2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_403), .Y(n_399) );
OR2x2_ASAP7_75t_L g666 ( .A(n_400), .B(n_403), .Y(n_666) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g410 ( .A(n_403), .Y(n_410) );
INVx1_ASAP7_75t_L g489 ( .A(n_403), .Y(n_489) );
INVx4_ASAP7_75t_L g574 ( .A(n_405), .Y(n_574) );
INVx3_ASAP7_75t_L g626 ( .A(n_405), .Y(n_626) );
OAI221xp5_ASAP7_75t_L g1122 ( .A1(n_405), .A2(n_587), .B1(n_1123), .B2(n_1124), .C(n_1125), .Y(n_1122) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx2_ASAP7_75t_L g557 ( .A(n_406), .Y(n_557) );
BUFx3_ASAP7_75t_L g800 ( .A(n_406), .Y(n_800) );
INVx3_ASAP7_75t_L g1016 ( .A(n_408), .Y(n_1016) );
OR2x6_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx2_ASAP7_75t_L g550 ( .A(n_409), .Y(n_550) );
OR2x2_ASAP7_75t_L g917 ( .A(n_409), .B(n_410), .Y(n_917) );
INVx3_ASAP7_75t_L g1026 ( .A(n_411), .Y(n_1026) );
INVx3_ASAP7_75t_L g1175 ( .A(n_411), .Y(n_1175) );
NOR3xp33_ASAP7_75t_L g1489 ( .A(n_411), .B(n_1490), .C(n_1499), .Y(n_1489) );
OAI21xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_451), .B(n_478), .Y(n_412) );
INVx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g1057 ( .A1(n_415), .A2(n_442), .B1(n_1030), .B2(n_1058), .C(n_1059), .Y(n_1057) );
AOI221xp5_ASAP7_75t_L g1182 ( .A1(n_415), .A2(n_442), .B1(n_1159), .B2(n_1183), .C(n_1188), .Y(n_1182) );
INVx2_ASAP7_75t_SL g1503 ( .A(n_415), .Y(n_1503) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_419), .Y(n_415) );
BUFx2_ASAP7_75t_L g956 ( .A(n_416), .Y(n_956) );
HB1xp67_ASAP7_75t_L g1509 ( .A(n_416), .Y(n_1509) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx3_ASAP7_75t_L g441 ( .A(n_417), .Y(n_441) );
INVx2_ASAP7_75t_L g539 ( .A(n_417), .Y(n_539) );
BUFx3_ASAP7_75t_L g777 ( .A(n_417), .Y(n_777) );
AND2x4_ASAP7_75t_L g450 ( .A(n_419), .B(n_433), .Y(n_450) );
AND2x4_ASAP7_75t_SL g455 ( .A(n_419), .B(n_443), .Y(n_455) );
AND2x2_ASAP7_75t_L g598 ( .A(n_419), .B(n_433), .Y(n_598) );
AOI21xp5_ASAP7_75t_SL g421 ( .A1(n_422), .A2(n_438), .B(n_442), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g771 ( .A(n_426), .Y(n_771) );
BUFx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g1186 ( .A(n_427), .Y(n_1186) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_428), .Y(n_443) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g1460 ( .A(n_432), .Y(n_1460) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_433), .Y(n_475) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx3_ASAP7_75t_L g770 ( .A(n_434), .Y(n_770) );
INVx2_ASAP7_75t_L g897 ( .A(n_434), .Y(n_897) );
INVx4_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_437), .B(n_519), .Y(n_518) );
AND2x4_ASAP7_75t_L g722 ( .A(n_437), .B(n_519), .Y(n_722) );
INVx4_ASAP7_75t_L g989 ( .A(n_437), .Y(n_989) );
INVx1_ASAP7_75t_SL g1507 ( .A(n_437), .Y(n_1507) );
INVx2_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g955 ( .A(n_440), .Y(n_955) );
INVx2_ASAP7_75t_L g1457 ( .A(n_440), .Y(n_1457) );
AOI21xp5_ASAP7_75t_L g987 ( .A1(n_442), .A2(n_988), .B(n_990), .Y(n_987) );
AOI21xp5_ASAP7_75t_L g1455 ( .A1(n_442), .A2(n_1456), .B(n_1458), .Y(n_1455) );
AOI21xp5_ASAP7_75t_L g1504 ( .A1(n_442), .A2(n_1505), .B(n_1508), .Y(n_1504) );
BUFx3_ASAP7_75t_L g473 ( .A(n_443), .Y(n_473) );
INVx1_ASAP7_75t_L g828 ( .A(n_443), .Y(n_828) );
BUFx3_ASAP7_75t_L g835 ( .A(n_443), .Y(n_835) );
BUFx3_ASAP7_75t_L g898 ( .A(n_443), .Y(n_898) );
BUFx6f_ASAP7_75t_L g1052 ( .A(n_443), .Y(n_1052) );
BUFx3_ASAP7_75t_L g1194 ( .A(n_443), .Y(n_1194) );
AOI22xp5_ASAP7_75t_L g1461 ( .A1(n_445), .A2(n_1181), .B1(n_1462), .B2(n_1463), .Y(n_1461) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g488 ( .A(n_447), .B(n_489), .Y(n_488) );
BUFx6f_ASAP7_75t_L g993 ( .A(n_447), .Y(n_993) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_450), .A2(n_993), .B1(n_994), .B2(n_995), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_450), .A2(n_993), .B1(n_1062), .B2(n_1063), .Y(n_1061) );
BUFx6f_ASAP7_75t_L g1181 ( .A(n_450), .Y(n_1181) );
AOI22xp33_ASAP7_75t_L g1510 ( .A1(n_450), .A2(n_993), .B1(n_1511), .B2(n_1512), .Y(n_1510) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g975 ( .A(n_453), .Y(n_975) );
INVx2_ASAP7_75t_L g1465 ( .A(n_453), .Y(n_1465) );
INVx4_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx3_ASAP7_75t_L g1050 ( .A(n_455), .Y(n_1050) );
BUFx2_ASAP7_75t_L g1514 ( .A(n_456), .Y(n_1514) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g1466 ( .A(n_457), .Y(n_1466) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g501 ( .A(n_459), .Y(n_501) );
BUFx2_ASAP7_75t_L g1056 ( .A(n_459), .Y(n_1056) );
OAI221xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_465), .B1(n_466), .B2(n_471), .C(n_472), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g982 ( .A(n_463), .Y(n_982) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx4_ASAP7_75t_L g833 ( .A(n_464), .Y(n_833) );
INVx3_ASAP7_75t_L g901 ( .A(n_464), .Y(n_901) );
OAI22xp33_ASAP7_75t_L g899 ( .A1(n_466), .A2(n_900), .B1(n_901), .B2(n_902), .Y(n_899) );
INVx6_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx4_ASAP7_75t_L g506 ( .A(n_468), .Y(n_506) );
INVx2_ASAP7_75t_L g528 ( .A(n_468), .Y(n_528) );
INVx2_ASAP7_75t_SL g841 ( .A(n_468), .Y(n_841) );
INVx1_ASAP7_75t_L g985 ( .A(n_468), .Y(n_985) );
INVx8_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx2_ASAP7_75t_L g648 ( .A(n_469), .Y(n_648) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OAI221xp5_ASAP7_75t_L g976 ( .A1(n_477), .A2(n_524), .B1(n_977), .B2(n_978), .C(n_979), .Y(n_976) );
INVx3_ASAP7_75t_L g1053 ( .A(n_477), .Y(n_1053) );
INVx1_ASAP7_75t_L g1195 ( .A(n_477), .Y(n_1195) );
INVx2_ASAP7_75t_L g1474 ( .A(n_477), .Y(n_1474) );
A2O1A1Ixp33_ASAP7_75t_SL g548 ( .A1(n_478), .A2(n_549), .B(n_566), .C(n_594), .Y(n_548) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_SL g608 ( .A1(n_480), .A2(n_609), .B(n_633), .C(n_638), .Y(n_608) );
INVx1_ASAP7_75t_L g944 ( .A(n_480), .Y(n_944) );
BUFx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
HB1xp67_ASAP7_75t_L g1141 ( .A(n_481), .Y(n_1141) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g602 ( .A(n_484), .Y(n_602) );
XOR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_599), .Y(n_484) );
NOR2x1_ASAP7_75t_SL g485 ( .A(n_486), .B(n_548), .Y(n_485) );
INVx1_ASAP7_75t_L g640 ( .A(n_487), .Y(n_640) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_488), .B(n_725), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_488), .A2(n_702), .B1(n_736), .B2(n_760), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_488), .B(n_843), .Y(n_842) );
AOI222xp33_ASAP7_75t_L g914 ( .A1(n_488), .A2(n_597), .B1(n_915), .B2(n_916), .C1(n_919), .C2(n_920), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_488), .B(n_1097), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_488), .B(n_1139), .Y(n_1142) );
AND2x4_ASAP7_75t_L g597 ( .A(n_489), .B(n_598), .Y(n_597) );
NOR3xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_498), .C(n_502), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g844 ( .A1(n_491), .A2(n_541), .B(n_845), .Y(n_844) );
NOR3xp33_ASAP7_75t_L g1147 ( .A(n_491), .B(n_1148), .C(n_1154), .Y(n_1147) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_492), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g778 ( .A1(n_492), .A2(n_779), .B(n_783), .Y(n_778) );
OAI21xp5_ASAP7_75t_L g903 ( .A1(n_492), .A2(n_781), .B(n_904), .Y(n_903) );
OAI21xp5_ASAP7_75t_SL g946 ( .A1(n_492), .A2(n_947), .B(n_950), .Y(n_946) );
OR2x6_ASAP7_75t_L g492 ( .A(n_493), .B(n_495), .Y(n_492) );
INVx4_ASAP7_75t_L g514 ( .A(n_493), .Y(n_514) );
BUFx4f_ASAP7_75t_L g522 ( .A(n_493), .Y(n_522) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_493), .Y(n_656) );
BUFx4f_ASAP7_75t_L g959 ( .A(n_493), .Y(n_959) );
BUFx4f_ASAP7_75t_L g977 ( .A(n_493), .Y(n_977) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx3_ASAP7_75t_L g543 ( .A(n_494), .Y(n_543) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2x2_ASAP7_75t_L g499 ( .A(n_496), .B(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_SL g665 ( .A(n_499), .Y(n_665) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_499), .Y(n_709) );
INVx1_ASAP7_75t_L g820 ( .A(n_499), .Y(n_820) );
INVx2_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_521), .Y(n_502) );
OAI211xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .B(n_507), .C(n_511), .Y(n_503) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_506), .A2(n_808), .B1(n_832), .B2(n_833), .Y(n_831) );
INVx3_ASAP7_75t_L g524 ( .A(n_508), .Y(n_524) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OAI221xp5_ASAP7_75t_L g1149 ( .A1(n_509), .A2(n_522), .B1(n_1124), .B2(n_1131), .C(n_1150), .Y(n_1149) );
BUFx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g652 ( .A(n_510), .Y(n_652) );
BUFx2_ASAP7_75t_L g655 ( .A(n_510), .Y(n_655) );
BUFx2_ASAP7_75t_L g786 ( .A(n_510), .Y(n_786) );
INVx2_ASAP7_75t_L g952 ( .A(n_510), .Y(n_952) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OAI221xp5_ASAP7_75t_L g783 ( .A1(n_513), .A2(n_745), .B1(n_784), .B2(n_787), .C(n_788), .Y(n_783) );
OAI221xp5_ASAP7_75t_L g904 ( .A1(n_513), .A2(n_524), .B1(n_905), .B2(n_906), .C(n_907), .Y(n_904) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g1079 ( .A(n_514), .Y(n_1079) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_516), .A2(n_646), .B1(n_647), .B2(n_648), .Y(n_645) );
OAI221xp5_ASAP7_75t_L g1467 ( .A1(n_516), .A2(n_1468), .B1(n_1469), .B2(n_1470), .C(n_1471), .Y(n_1467) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_SL g659 ( .A(n_517), .Y(n_659) );
INVx1_ASAP7_75t_L g772 ( .A(n_518), .Y(n_772) );
OAI22xp5_ASAP7_75t_SL g1148 ( .A1(n_518), .A2(n_644), .B1(n_1149), .B2(n_1151), .Y(n_1148) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OAI221xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_524), .B2(n_525), .C(n_526), .Y(n_521) );
OAI221xp5_ASAP7_75t_L g950 ( .A1(n_522), .A2(n_941), .B1(n_951), .B2(n_953), .C(n_954), .Y(n_950) );
OAI221xp5_ASAP7_75t_L g584 ( .A1(n_525), .A2(n_573), .B1(n_585), .B2(n_586), .C(n_587), .Y(n_584) );
INVxp33_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_SL g949 ( .A(n_529), .Y(n_949) );
INVx4_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g644 ( .A(n_530), .Y(n_644) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_530), .Y(n_716) );
INVx2_ASAP7_75t_L g782 ( .A(n_530), .Y(n_782) );
AOI222xp33_ASAP7_75t_L g824 ( .A1(n_530), .A2(n_545), .B1(n_722), .B2(n_825), .C1(n_826), .C2(n_834), .Y(n_824) );
AND2x4_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g699 ( .A(n_531), .Y(n_699) );
OR2x6_ASAP7_75t_L g1042 ( .A(n_531), .B(n_581), .Y(n_1042) );
AOI222xp33_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B1(n_540), .B2(n_541), .C1(n_544), .C2(n_545), .Y(n_533) );
AOI211xp5_ASAP7_75t_SL g549 ( .A1(n_534), .A2(n_550), .B(n_551), .C(n_559), .Y(n_549) );
AOI222xp33_ASAP7_75t_L g667 ( .A1(n_535), .A2(n_541), .B1(n_545), .B2(n_610), .C1(n_636), .C2(n_668), .Y(n_667) );
AOI211xp5_ASAP7_75t_L g705 ( .A1(n_535), .A2(n_674), .B(n_706), .C(n_708), .Y(n_705) );
AOI222xp33_ASAP7_75t_L g762 ( .A1(n_535), .A2(n_541), .B1(n_545), .B2(n_737), .C1(n_740), .C2(n_763), .Y(n_762) );
AOI222xp33_ASAP7_75t_L g819 ( .A1(n_535), .A2(n_810), .B1(n_820), .B2(n_821), .C1(n_822), .C2(n_823), .Y(n_819) );
INVxp67_ASAP7_75t_L g891 ( .A(n_535), .Y(n_891) );
INVx1_ASAP7_75t_L g918 ( .A(n_535), .Y(n_918) );
AOI222xp33_ASAP7_75t_L g1092 ( .A1(n_535), .A2(n_541), .B1(n_545), .B2(n_1093), .C1(n_1094), .C2(n_1095), .Y(n_1092) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
AOI332xp33_ASAP7_75t_L g1144 ( .A1(n_536), .A2(n_538), .A3(n_541), .B1(n_546), .B2(n_547), .B3(n_1135), .C1(n_1145), .C2(n_1146), .Y(n_1144) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g542 ( .A(n_537), .B(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g707 ( .A(n_537), .B(n_543), .Y(n_707) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx3_ASAP7_75t_L g653 ( .A(n_543), .Y(n_653) );
AOI222xp33_ASAP7_75t_L g710 ( .A1(n_545), .A2(n_711), .B1(n_716), .B2(n_717), .C1(n_722), .C2(n_723), .Y(n_710) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
AOI211xp5_ASAP7_75t_L g609 ( .A1(n_550), .A2(n_610), .B(n_611), .C(n_612), .Y(n_609) );
AOI211xp5_ASAP7_75t_L g673 ( .A1(n_550), .A2(n_674), .B(n_675), .C(n_676), .Y(n_673) );
INVx2_ASAP7_75t_L g734 ( .A(n_550), .Y(n_734) );
AOI211xp5_ASAP7_75t_SL g809 ( .A1(n_550), .A2(n_810), .B(n_811), .C(n_812), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_550), .A2(n_872), .B1(n_875), .B2(n_885), .Y(n_871) );
AOI221xp5_ASAP7_75t_L g1099 ( .A1(n_550), .A2(n_1094), .B1(n_1100), .B2(n_1102), .C(n_1103), .Y(n_1099) );
AOI221xp5_ASAP7_75t_L g1134 ( .A1(n_550), .A2(n_1102), .B1(n_1135), .B2(n_1136), .C(n_1140), .Y(n_1134) );
INVx4_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AOI221xp5_ASAP7_75t_L g738 ( .A1(n_553), .A2(n_555), .B1(n_739), .B2(n_740), .C(n_741), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g868 ( .A1(n_553), .A2(n_555), .B1(n_741), .B2(n_869), .C(n_870), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_553), .A2(n_555), .B1(n_927), .B2(n_928), .Y(n_926) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g741 ( .A(n_556), .Y(n_741) );
OR2x6_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
OAI221xp5_ASAP7_75t_L g1127 ( .A1(n_557), .A2(n_578), .B1(n_580), .B2(n_1128), .C(n_1129), .Y(n_1127) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_560), .Y(n_634) );
OR2x6_ASAP7_75t_SL g560 ( .A(n_561), .B(n_563), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_562), .Y(n_874) );
INVx3_ASAP7_75t_L g1001 ( .A(n_563), .Y(n_1001) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_565), .A2(n_634), .B1(n_635), .B2(n_636), .C(n_637), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_565), .A2(n_634), .B1(n_736), .B2(n_737), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_565), .B(n_699), .Y(n_966) );
NOR3xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_582), .C(n_588), .Y(n_566) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_569), .Y(n_691) );
INVx2_ASAP7_75t_L g1125 ( .A(n_569), .Y(n_1125) );
INVx2_ASAP7_75t_L g1440 ( .A(n_569), .Y(n_1440) );
OAI221xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B1(n_575), .B2(n_576), .C(n_580), .Y(n_571) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g615 ( .A(n_574), .Y(n_615) );
OAI221xp5_ASAP7_75t_L g935 ( .A1(n_576), .A2(n_580), .B1(n_936), .B2(n_938), .C(n_939), .Y(n_935) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI221xp5_ASAP7_75t_L g806 ( .A1(n_578), .A2(n_580), .B1(n_800), .B2(n_807), .C(n_808), .Y(n_806) );
BUFx4f_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx3_ASAP7_75t_L g695 ( .A(n_579), .Y(n_695) );
BUFx3_ASAP7_75t_L g1110 ( .A(n_579), .Y(n_1110) );
INVx2_ASAP7_75t_L g1446 ( .A(n_579), .Y(n_1446) );
INVx3_ASAP7_75t_L g617 ( .A(n_580), .Y(n_617) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_580), .A2(n_625), .B1(n_694), .B2(n_695), .C(n_696), .Y(n_693) );
OAI221xp5_ASAP7_75t_L g1109 ( .A1(n_580), .A2(n_800), .B1(n_1076), .B2(n_1086), .C(n_1110), .Y(n_1109) );
INVx3_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_583), .A2(n_861), .B1(n_919), .B2(n_925), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_586), .A2(n_619), .B1(n_620), .B2(n_622), .Y(n_618) );
INVx1_ASAP7_75t_L g805 ( .A(n_586), .Y(n_805) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_587), .A2(n_625), .B1(n_686), .B2(n_687), .C(n_688), .Y(n_685) );
OAI221xp5_ASAP7_75t_L g799 ( .A1(n_587), .A2(n_800), .B1(n_801), .B2(n_802), .C(n_803), .Y(n_799) );
OAI221xp5_ASAP7_75t_L g1106 ( .A1(n_587), .A2(n_800), .B1(n_1081), .B2(n_1085), .C(n_1107), .Y(n_1106) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_590), .A2(n_593), .B1(n_760), .B2(n_761), .Y(n_759) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_596), .B(n_893), .Y(n_892) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_597), .B(n_635), .Y(n_669) );
INVx1_ASAP7_75t_L g703 ( .A(n_597), .Y(n_703) );
INVx1_ASAP7_75t_L g817 ( .A(n_597), .Y(n_817) );
NAND2xp33_ASAP7_75t_SL g1113 ( .A(n_597), .B(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g849 ( .A(n_603), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_728), .B1(n_846), .B2(n_847), .Y(n_603) );
INVx1_ASAP7_75t_L g846 ( .A(n_604), .Y(n_846) );
OA22x2_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_670), .B1(n_726), .B2(n_727), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx2_ASAP7_75t_SL g727 ( .A(n_606), .Y(n_727) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_641), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_618), .B(n_623), .Y(n_612) );
OAI21xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B(n_616), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_614), .A2(n_624), .B1(n_655), .B2(n_656), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_619), .A2(n_650), .B1(n_651), .B2(n_653), .Y(n_649) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_622), .A2(n_648), .B1(n_658), .B2(n_660), .Y(n_657) );
OAI211xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B(n_627), .C(n_631), .Y(n_623) );
INVx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g755 ( .A(n_626), .Y(n_755) );
INVx2_ASAP7_75t_L g1101 ( .A(n_626), .Y(n_1101) );
INVx5_ASAP7_75t_L g744 ( .A(n_628), .Y(n_744) );
INVx2_ASAP7_75t_SL g802 ( .A(n_628), .Y(n_802) );
INVx2_ASAP7_75t_SL g865 ( .A(n_628), .Y(n_865) );
INVx3_ASAP7_75t_L g876 ( .A(n_628), .Y(n_876) );
BUFx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g752 ( .A(n_632), .Y(n_752) );
BUFx2_ASAP7_75t_L g758 ( .A(n_632), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_667), .C(n_669), .Y(n_641) );
NOR2xp33_ASAP7_75t_SL g642 ( .A(n_643), .B(n_663), .Y(n_642) );
OAI33xp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .A3(n_649), .B1(n_654), .B2(n_657), .B3(n_661), .Y(n_643) );
OAI33xp33_ASAP7_75t_L g1073 ( .A1(n_644), .A2(n_1074), .A3(n_1077), .B1(n_1082), .B2(n_1087), .B3(n_1090), .Y(n_1073) );
OAI22xp33_ASAP7_75t_L g712 ( .A1(n_648), .A2(n_696), .B1(n_713), .B2(n_714), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_648), .A2(n_719), .B1(n_720), .B2(n_721), .Y(n_718) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g1082 ( .A1(n_653), .A2(n_1083), .B1(n_1085), .B2(n_1086), .Y(n_1082) );
OAI221xp5_ASAP7_75t_L g1151 ( .A1(n_656), .A2(n_1123), .B1(n_1128), .B2(n_1152), .C(n_1153), .Y(n_1151) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g1090 ( .A(n_662), .Y(n_1090) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g726 ( .A(n_670), .Y(n_726) );
OR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_704), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_SL g672 ( .A1(n_673), .A2(n_677), .B(n_697), .C(n_700), .Y(n_672) );
NOR3xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_689), .C(n_690), .Y(n_677) );
BUFx2_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_682), .B(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g1168 ( .A(n_682), .Y(n_1168) );
BUFx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_687), .A2(n_941), .B1(n_942), .B2(n_943), .Y(n_940) );
O2A1O1Ixp33_ASAP7_75t_SL g973 ( .A1(n_697), .A2(n_974), .B(n_986), .C(n_996), .Y(n_973) );
AOI21xp5_ASAP7_75t_SL g1176 ( .A1(n_697), .A2(n_1177), .B(n_1199), .Y(n_1176) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OAI21xp5_ASAP7_75t_L g732 ( .A1(n_698), .A2(n_733), .B(n_742), .Y(n_732) );
INVx2_ASAP7_75t_L g813 ( .A(n_698), .Y(n_813) );
AOI21xp5_ASAP7_75t_L g856 ( .A1(n_698), .A2(n_857), .B(n_886), .Y(n_856) );
BUFx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_710), .C(n_724), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_714), .A2(n_841), .B1(n_1088), .B2(n_1089), .Y(n_1087) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g1074 ( .A1(n_720), .A2(n_841), .B1(n_1075), .B2(n_1076), .Y(n_1074) );
AOI211xp5_ASAP7_75t_L g894 ( .A1(n_722), .A2(n_895), .B(n_903), .C(n_908), .Y(n_894) );
CKINVDCx5p33_ASAP7_75t_R g961 ( .A(n_722), .Y(n_961) );
INVx1_ASAP7_75t_L g847 ( .A(n_728), .Y(n_847) );
XOR2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_792), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g790 ( .A(n_731), .Y(n_790) );
NAND4xp25_ASAP7_75t_L g731 ( .A(n_732), .B(n_762), .C(n_764), .D(n_789), .Y(n_731) );
NOR3xp33_ASAP7_75t_L g1104 ( .A(n_741), .B(n_1105), .C(n_1108), .Y(n_1104) );
NOR3xp33_ASAP7_75t_L g1120 ( .A(n_741), .B(n_1121), .C(n_1126), .Y(n_1120) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_753), .C(n_759), .Y(n_742) );
OAI221xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B1(n_746), .B2(n_748), .C(n_749), .Y(n_743) );
INVx8_ASAP7_75t_L g1038 ( .A(n_744), .Y(n_1038) );
INVx3_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
CKINVDCx8_ASAP7_75t_R g942 ( .A(n_747), .Y(n_942) );
INVx3_ASAP7_75t_L g1112 ( .A(n_747), .Y(n_1112) );
INVx3_ASAP7_75t_L g1132 ( .A(n_747), .Y(n_1132) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI211xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .B(n_756), .C(n_757), .Y(n_753) );
HB1xp67_ASAP7_75t_L g931 ( .A(n_755), .Y(n_931) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_765), .B(n_778), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_772), .C(n_773), .Y(n_766) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g830 ( .A(n_770), .Y(n_830) );
BUFx2_ASAP7_75t_L g1187 ( .A(n_770), .Y(n_1187) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g1060 ( .A(n_775), .Y(n_1060) );
INVx3_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
BUFx6f_ASAP7_75t_L g991 ( .A(n_776), .Y(n_991) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
OAI221xp5_ASAP7_75t_L g958 ( .A1(n_784), .A2(n_930), .B1(n_938), .B2(n_959), .C(n_960), .Y(n_958) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx4_ASAP7_75t_L g1080 ( .A(n_785), .Y(n_1080) );
INVx4_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
OAI221xp5_ASAP7_75t_L g1299 ( .A1(n_791), .A2(n_1300), .B1(n_1301), .B2(n_1302), .C(n_1303), .Y(n_1299) );
OR2x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_818), .Y(n_793) );
A2O1A1Ixp33_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_809), .B(n_813), .C(n_814), .Y(n_794) );
NOR3xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .C(n_804), .Y(n_795) );
INVx2_ASAP7_75t_L g937 ( .A(n_800), .Y(n_937) );
INVx2_ASAP7_75t_L g862 ( .A(n_802), .Y(n_862) );
A2O1A1Ixp33_ASAP7_75t_L g1098 ( .A1(n_813), .A2(n_1099), .B(n_1104), .C(n_1113), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
NAND4xp25_ASAP7_75t_L g818 ( .A(n_819), .B(n_824), .C(n_842), .D(n_844), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g962 ( .A1(n_820), .A2(n_822), .B1(n_925), .B2(n_927), .Y(n_962) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_838), .B1(n_840), .B2(n_841), .Y(n_836) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
HB1xp67_ASAP7_75t_L g1469 ( .A(n_841), .Y(n_1469) );
INVx1_ASAP7_75t_L g1202 ( .A(n_850), .Y(n_1202) );
HB1xp67_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
XNOR2x1_ASAP7_75t_L g851 ( .A(n_852), .B(n_1155), .Y(n_851) );
XNOR2x1_ASAP7_75t_L g852 ( .A(n_853), .B(n_968), .Y(n_852) );
XNOR2x2_ASAP7_75t_L g853 ( .A(n_854), .B(n_911), .Y(n_853) );
AOI21xp5_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_909), .B(n_910), .Y(n_854) );
AND3x1_ASAP7_75t_L g855 ( .A(n_856), .B(n_887), .C(n_894), .Y(n_855) );
AOI31xp33_ASAP7_75t_L g910 ( .A1(n_856), .A2(n_887), .A3(n_894), .B(n_909), .Y(n_910) );
NAND3xp33_ASAP7_75t_SL g857 ( .A(n_858), .B(n_868), .C(n_871), .Y(n_857) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_860), .B1(n_863), .B2(n_866), .Y(n_858) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVxp67_ASAP7_75t_L g923 ( .A(n_872), .Y(n_923) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_874), .Y(n_1102) );
OAI22xp5_ASAP7_75t_L g1130 ( .A1(n_876), .A2(n_1131), .B1(n_1132), .B2(n_1133), .Y(n_1130) );
INVx3_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
BUFx2_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
AND2x2_ASAP7_75t_L g887 ( .A(n_888), .B(n_892), .Y(n_887) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx2_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx2_ASAP7_75t_L g1193 ( .A(n_897), .Y(n_1193) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
NAND3xp33_ASAP7_75t_L g913 ( .A(n_914), .B(n_921), .C(n_945), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_917), .B(n_918), .Y(n_916) );
OAI21xp33_ASAP7_75t_L g921 ( .A1(n_922), .A2(n_934), .B(n_944), .Y(n_921) );
OAI211xp5_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_924), .B(n_926), .C(n_929), .Y(n_922) );
OAI211xp5_ASAP7_75t_L g929 ( .A1(n_930), .A2(n_931), .B(n_932), .C(n_933), .Y(n_929) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g1064 ( .A(n_944), .Y(n_1064) );
NOR3xp33_ASAP7_75t_L g945 ( .A(n_946), .B(n_957), .C(n_963), .Y(n_945) );
INVxp67_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx2_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
BUFx2_ASAP7_75t_L g1084 ( .A(n_952), .Y(n_1084) );
INVx2_ASAP7_75t_L g1152 ( .A(n_952), .Y(n_1152) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
XNOR2xp5_ASAP7_75t_L g968 ( .A(n_969), .B(n_1067), .Y(n_968) );
XNOR2xp5_ASAP7_75t_L g969 ( .A(n_970), .B(n_1027), .Y(n_969) );
NOR2x1p5_ASAP7_75t_L g971 ( .A(n_972), .B(n_1003), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_982), .B1(n_983), .B2(n_984), .Y(n_980) );
BUFx3_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_993), .A2(n_1179), .B1(n_1180), .B2(n_1181), .Y(n_1178) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_994), .A2(n_995), .B1(n_999), .B2(n_1000), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_999), .A2(n_1000), .B1(n_1062), .B2(n_1063), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1002), .Y(n_1000) );
INVx2_ASAP7_75t_L g1107 ( .A(n_1001), .Y(n_1107) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1001), .Y(n_1137) );
INVxp67_ASAP7_75t_L g1447 ( .A(n_1002), .Y(n_1447) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1007), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1006), .Y(n_1004) );
AOI221xp5_ASAP7_75t_L g1029 ( .A1(n_1005), .A2(n_1016), .B1(n_1030), .B2(n_1031), .C(n_1032), .Y(n_1029) );
AOI221xp5_ASAP7_75t_L g1158 ( .A1(n_1005), .A2(n_1016), .B1(n_1159), .B2(n_1160), .C(n_1161), .Y(n_1158) );
AOI21xp33_ASAP7_75t_SL g1450 ( .A1(n_1005), .A2(n_1451), .B(n_1452), .Y(n_1450) );
AOI21xp33_ASAP7_75t_L g1486 ( .A1(n_1005), .A2(n_1487), .B(n_1488), .Y(n_1486) );
AND4x1_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1014), .C(n_1017), .D(n_1026), .Y(n_1007) );
AOI22xp5_ASAP7_75t_L g1008 ( .A1(n_1009), .A2(n_1010), .B1(n_1012), .B2(n_1013), .Y(n_1008) );
INVx2_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1016), .Y(n_1014) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
BUFx2_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
BUFx2_ASAP7_75t_L g1173 ( .A(n_1025), .Y(n_1173) );
NAND3xp33_ASAP7_75t_L g1032 ( .A(n_1026), .B(n_1033), .C(n_1043), .Y(n_1032) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1026), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1047), .Y(n_1028) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
AOI222xp33_ASAP7_75t_L g1049 ( .A1(n_1044), .A2(n_1046), .B1(n_1050), .B2(n_1051), .C1(n_1054), .C2(n_1055), .Y(n_1049) );
AOI21xp5_ASAP7_75t_L g1047 ( .A1(n_1048), .A2(n_1064), .B(n_1065), .Y(n_1047) );
NAND3xp33_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1057), .C(n_1061), .Y(n_1048) );
AOI222xp33_ASAP7_75t_L g1189 ( .A1(n_1050), .A2(n_1163), .B1(n_1164), .B2(n_1190), .C1(n_1196), .C2(n_1197), .Y(n_1189) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1055), .Y(n_1198) );
OAI21xp5_ASAP7_75t_L g1501 ( .A1(n_1064), .A2(n_1502), .B(n_1513), .Y(n_1501) );
XNOR2x1_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1115), .Y(n_1067) );
XNOR2x1_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1070), .Y(n_1068) );
NOR2x1_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1098), .Y(n_1070) );
NAND3xp33_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1092), .C(n_1096), .Y(n_1071) );
NOR2xp33_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1091), .Y(n_1072) );
OAI22xp5_ASAP7_75t_L g1077 ( .A1(n_1078), .A2(n_1079), .B1(n_1080), .B2(n_1081), .Y(n_1077) );
OAI211xp5_ASAP7_75t_SL g1515 ( .A1(n_1079), .A2(n_1516), .B(n_1517), .C(n_1518), .Y(n_1515) );
INVx4_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
XNOR2x1_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1118), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1143), .Y(n_1118) );
A2O1A1Ixp33_ASAP7_75t_L g1119 ( .A1(n_1120), .A2(n_1134), .B(n_1141), .C(n_1142), .Y(n_1119) );
BUFx3_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1176), .Y(n_1157) );
NAND3xp33_ASAP7_75t_SL g1161 ( .A(n_1162), .B(n_1165), .C(n_1175), .Y(n_1161) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
NAND3xp33_ASAP7_75t_SL g1177 ( .A(n_1178), .B(n_1182), .C(n_1189), .Y(n_1177) );
INVx2_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
INVx2_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
INVx2_ASAP7_75t_L g1506 ( .A(n_1192), .Y(n_1506) );
INVx2_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1193), .Y(n_1473) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
OAI221xp5_ASAP7_75t_L g1203 ( .A1(n_1204), .A2(n_1422), .B1(n_1425), .B2(n_1428), .C(n_1476), .Y(n_1203) );
AND4x1_ASAP7_75t_L g1204 ( .A(n_1205), .B(n_1325), .C(n_1376), .D(n_1407), .Y(n_1204) );
O2A1O1Ixp33_ASAP7_75t_L g1205 ( .A1(n_1206), .A2(n_1262), .B(n_1296), .C(n_1304), .Y(n_1205) );
OAI221xp5_ASAP7_75t_L g1206 ( .A1(n_1207), .A2(n_1232), .B1(n_1242), .B2(n_1245), .C(n_1251), .Y(n_1206) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1207), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1400 ( .A(n_1207), .B(n_1401), .Y(n_1400) );
OR2x2_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1224), .Y(n_1207) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1208), .B(n_1368), .Y(n_1375) );
CKINVDCx5p33_ASAP7_75t_R g1208 ( .A(n_1209), .Y(n_1208) );
NOR2xp33_ASAP7_75t_L g1264 ( .A(n_1209), .B(n_1265), .Y(n_1264) );
O2A1O1Ixp33_ASAP7_75t_L g1285 ( .A1(n_1209), .A2(n_1286), .B(n_1287), .C(n_1291), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1209), .B(n_1282), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1209), .B(n_1267), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1209), .B(n_1318), .Y(n_1395) );
NAND2xp5_ASAP7_75t_L g1404 ( .A(n_1209), .B(n_1405), .Y(n_1404) );
INVx4_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
INVx4_ASAP7_75t_L g1272 ( .A(n_1210), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1210), .B(n_1307), .Y(n_1306) );
NAND2xp5_ASAP7_75t_SL g1316 ( .A(n_1210), .B(n_1229), .Y(n_1316) );
OR2x2_ASAP7_75t_L g1322 ( .A(n_1210), .B(n_1229), .Y(n_1322) );
NOR2xp33_ASAP7_75t_L g1335 ( .A(n_1210), .B(n_1336), .Y(n_1335) );
NOR2xp33_ASAP7_75t_L g1347 ( .A(n_1210), .B(n_1290), .Y(n_1347) );
NOR2xp33_ASAP7_75t_L g1392 ( .A(n_1210), .B(n_1359), .Y(n_1392) );
AND2x4_ASAP7_75t_SL g1210 ( .A(n_1211), .B(n_1219), .Y(n_1210) );
AND2x4_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1214), .Y(n_1212) );
AND2x6_ASAP7_75t_L g1217 ( .A(n_1213), .B(n_1218), .Y(n_1217) );
AND2x6_ASAP7_75t_L g1220 ( .A(n_1213), .B(n_1221), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1213), .B(n_1223), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1213), .B(n_1223), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1213), .B(n_1223), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_1213), .B(n_1214), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1216), .Y(n_1214) );
INVx2_ASAP7_75t_L g1302 ( .A(n_1217), .Y(n_1302) );
INVx2_ASAP7_75t_L g1424 ( .A(n_1220), .Y(n_1424) );
OAI21xp5_ASAP7_75t_L g1520 ( .A1(n_1221), .A2(n_1521), .B(n_1522), .Y(n_1520) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1224), .B(n_1273), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1229), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1225), .B(n_1248), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1225), .B(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1225), .Y(n_1276) );
OR2x2_ASAP7_75t_L g1284 ( .A(n_1225), .B(n_1274), .Y(n_1284) );
OR2x2_ASAP7_75t_L g1290 ( .A(n_1225), .B(n_1248), .Y(n_1290) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1225), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1228), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1229), .B(n_1247), .Y(n_1246) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1229), .Y(n_1268) );
OR2x2_ASAP7_75t_L g1286 ( .A(n_1229), .B(n_1248), .Y(n_1286) );
OR2x2_ASAP7_75t_L g1336 ( .A(n_1229), .B(n_1253), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_1229), .B(n_1253), .Y(n_1356) );
OR2x2_ASAP7_75t_L g1416 ( .A(n_1229), .B(n_1334), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1231), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1230), .B(n_1231), .Y(n_1274) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1234), .B(n_1238), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1234), .B(n_1244), .Y(n_1243) );
INVx3_ASAP7_75t_L g1256 ( .A(n_1234), .Y(n_1256) );
NOR2xp33_ASAP7_75t_SL g1324 ( .A(n_1234), .B(n_1298), .Y(n_1324) );
A2O1A1Ixp33_ASAP7_75t_L g1325 ( .A1(n_1234), .A2(n_1326), .B(n_1348), .C(n_1361), .Y(n_1325) );
OR2x2_ASAP7_75t_L g1339 ( .A(n_1234), .B(n_1238), .Y(n_1339) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1234), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1236), .Y(n_1234) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1238), .Y(n_1244) );
OR2x2_ASAP7_75t_L g1277 ( .A(n_1238), .B(n_1258), .Y(n_1277) );
INVx2_ASAP7_75t_L g1279 ( .A(n_1238), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1238), .B(n_1256), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1333 ( .A(n_1238), .B(n_1320), .Y(n_1333) );
OR2x2_ASAP7_75t_L g1359 ( .A(n_1238), .B(n_1259), .Y(n_1359) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
OR2x2_ASAP7_75t_L g1257 ( .A(n_1239), .B(n_1258), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1241), .Y(n_1239) );
OAI222xp33_ASAP7_75t_L g1353 ( .A1(n_1242), .A2(n_1291), .B1(n_1354), .B2(n_1355), .C1(n_1357), .C2(n_1360), .Y(n_1353) );
AOI21xp33_ASAP7_75t_SL g1419 ( .A1(n_1242), .A2(n_1420), .B(n_1421), .Y(n_1419) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
NOR2xp33_ASAP7_75t_L g1310 ( .A(n_1244), .B(n_1272), .Y(n_1310) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1244), .Y(n_1406) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
O2A1O1Ixp33_ASAP7_75t_L g1370 ( .A1(n_1246), .A2(n_1371), .B(n_1372), .C(n_1373), .Y(n_1370) );
NAND2x1_ASAP7_75t_L g1421 ( .A(n_1246), .B(n_1272), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1247), .B(n_1315), .Y(n_1314) );
OAI221xp5_ASAP7_75t_L g1340 ( .A1(n_1247), .A2(n_1316), .B1(n_1341), .B2(n_1342), .C(n_1344), .Y(n_1340) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1247), .B(n_1352), .Y(n_1351) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1247), .Y(n_1374) );
OAI21xp5_ASAP7_75t_L g1410 ( .A1(n_1247), .A2(n_1288), .B(n_1411), .Y(n_1410) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1248), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1275 ( .A(n_1248), .B(n_1276), .Y(n_1275) );
NAND2x1p5_ASAP7_75t_L g1248 ( .A(n_1249), .B(n_1250), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1254), .Y(n_1251) );
NAND3xp33_ASAP7_75t_L g1293 ( .A(n_1252), .B(n_1294), .C(n_1295), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1252), .B(n_1268), .Y(n_1307) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1252), .Y(n_1341) );
NOR2xp33_ASAP7_75t_L g1267 ( .A(n_1253), .B(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
OR2x2_ASAP7_75t_L g1255 ( .A(n_1256), .B(n_1257), .Y(n_1255) );
OR2x2_ASAP7_75t_L g1291 ( .A(n_1256), .B(n_1282), .Y(n_1291) );
CKINVDCx14_ASAP7_75t_R g1295 ( .A(n_1256), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_1256), .B(n_1320), .Y(n_1327) );
O2A1O1Ixp33_ASAP7_75t_L g1376 ( .A1(n_1256), .A2(n_1377), .B(n_1388), .C(n_1393), .Y(n_1376) );
CKINVDCx5p33_ASAP7_75t_R g1368 ( .A(n_1257), .Y(n_1368) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1258), .Y(n_1282) );
NOR2xp33_ASAP7_75t_L g1380 ( .A(n_1258), .B(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1259), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1259 ( .A(n_1260), .B(n_1261), .Y(n_1259) );
A2O1A1Ixp33_ASAP7_75t_L g1262 ( .A1(n_1263), .A2(n_1269), .B(n_1277), .C(n_1278), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
HB1xp67_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1268), .B(n_1289), .Y(n_1288) );
OR2x2_ASAP7_75t_L g1360 ( .A(n_1268), .B(n_1290), .Y(n_1360) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1268), .B(n_1385), .Y(n_1384) );
OR2x2_ASAP7_75t_L g1387 ( .A(n_1268), .B(n_1275), .Y(n_1387) );
OAI211xp5_ASAP7_75t_L g1388 ( .A1(n_1269), .A2(n_1308), .B(n_1389), .C(n_1391), .Y(n_1388) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
NOR2xp33_ASAP7_75t_L g1270 ( .A(n_1271), .B(n_1273), .Y(n_1270) );
NOR2xp33_ASAP7_75t_L g1331 ( .A(n_1271), .B(n_1332), .Y(n_1331) );
NAND2xp5_ASAP7_75t_L g1344 ( .A(n_1271), .B(n_1289), .Y(n_1344) );
CKINVDCx5p33_ASAP7_75t_R g1271 ( .A(n_1272), .Y(n_1271) );
NOR2xp33_ASAP7_75t_L g1283 ( .A(n_1272), .B(n_1284), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1272), .B(n_1320), .Y(n_1343) );
NOR2x1_ASAP7_75t_L g1385 ( .A(n_1272), .B(n_1374), .Y(n_1385) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1272), .B(n_1399), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1418 ( .A(n_1272), .B(n_1299), .Y(n_1418) );
NOR2xp33_ASAP7_75t_L g1390 ( .A(n_1273), .B(n_1342), .Y(n_1390) );
OR2x2_ASAP7_75t_L g1273 ( .A(n_1274), .B(n_1275), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1274), .B(n_1347), .Y(n_1346) );
OR2x2_ASAP7_75t_L g1354 ( .A(n_1275), .B(n_1316), .Y(n_1354) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1275), .Y(n_1399) );
CKINVDCx5p33_ASAP7_75t_R g1318 ( .A(n_1277), .Y(n_1318) );
AOI211xp5_ASAP7_75t_L g1278 ( .A1(n_1279), .A2(n_1280), .B(n_1285), .C(n_1292), .Y(n_1278) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1279), .Y(n_1308) );
A2O1A1Ixp33_ASAP7_75t_L g1377 ( .A1(n_1279), .A2(n_1378), .B(n_1379), .C(n_1383), .Y(n_1377) );
AOI32xp33_ASAP7_75t_L g1414 ( .A1(n_1279), .A2(n_1333), .A3(n_1345), .B1(n_1415), .B2(n_1417), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1283), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1281), .B(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
NOR2xp33_ASAP7_75t_L g1403 ( .A(n_1282), .B(n_1404), .Y(n_1403) );
INVxp67_ASAP7_75t_L g1405 ( .A(n_1284), .Y(n_1405) );
AOI21xp5_ASAP7_75t_L g1373 ( .A1(n_1286), .A2(n_1374), .B(n_1375), .Y(n_1373) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1289), .B(n_1315), .Y(n_1382) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_1289), .B(n_1395), .Y(n_1394) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
OR2x2_ASAP7_75t_L g1321 ( .A(n_1290), .B(n_1322), .Y(n_1321) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1295), .B(n_1298), .Y(n_1363) );
AOI22xp33_ASAP7_75t_L g1393 ( .A1(n_1296), .A2(n_1394), .B1(n_1396), .B2(n_1402), .Y(n_1393) );
AOI221xp5_ASAP7_75t_L g1396 ( .A1(n_1296), .A2(n_1368), .B1(n_1397), .B2(n_1398), .C(n_1400), .Y(n_1396) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1296), .Y(n_1408) );
INVx2_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
AOI211xp5_ASAP7_75t_SL g1337 ( .A1(n_1297), .A2(n_1338), .B(n_1340), .C(n_1345), .Y(n_1337) );
OAI21xp33_ASAP7_75t_L g1350 ( .A1(n_1297), .A2(n_1318), .B(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
O2A1O1Ixp33_ASAP7_75t_SL g1304 ( .A1(n_1305), .A2(n_1308), .B(n_1309), .C(n_1323), .Y(n_1304) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
OAI31xp33_ASAP7_75t_L g1402 ( .A1(n_1306), .A2(n_1380), .A3(n_1403), .B(n_1406), .Y(n_1402) );
NAND2xp5_ASAP7_75t_L g1317 ( .A(n_1307), .B(n_1318), .Y(n_1317) );
AOI211xp5_ASAP7_75t_L g1309 ( .A1(n_1310), .A2(n_1311), .B(n_1312), .C(n_1319), .Y(n_1309) );
NAND2xp33_ASAP7_75t_SL g1312 ( .A(n_1313), .B(n_1317), .Y(n_1312) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1314), .Y(n_1378) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
OAI21xp5_ASAP7_75t_SL g1383 ( .A1(n_1318), .A2(n_1384), .B(n_1386), .Y(n_1383) );
NOR2xp33_ASAP7_75t_L g1319 ( .A(n_1320), .B(n_1321), .Y(n_1319) );
INVx2_ASAP7_75t_L g1372 ( .A(n_1320), .Y(n_1372) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1322), .Y(n_1352) );
AOI21xp5_ASAP7_75t_L g1349 ( .A1(n_1323), .A2(n_1350), .B(n_1353), .Y(n_1349) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
A2O1A1Ixp33_ASAP7_75t_L g1326 ( .A1(n_1327), .A2(n_1328), .B(n_1330), .C(n_1337), .Y(n_1326) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
AOI21xp5_ASAP7_75t_L g1330 ( .A1(n_1331), .A2(n_1334), .B(n_1335), .Y(n_1330) );
NOR2xp33_ASAP7_75t_L g1369 ( .A(n_1332), .B(n_1354), .Y(n_1369) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
AOI221xp5_ASAP7_75t_SL g1364 ( .A1(n_1333), .A2(n_1365), .B1(n_1367), .B2(n_1368), .C(n_1369), .Y(n_1364) );
CKINVDCx14_ASAP7_75t_R g1338 ( .A(n_1339), .Y(n_1338) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1347), .Y(n_1366) );
INVxp67_ASAP7_75t_SL g1348 ( .A(n_1349), .Y(n_1348) );
OAI211xp5_ASAP7_75t_L g1361 ( .A1(n_1349), .A2(n_1362), .B(n_1364), .C(n_1370), .Y(n_1361) );
CKINVDCx14_ASAP7_75t_R g1355 ( .A(n_1356), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1356), .B(n_1392), .Y(n_1391) );
A2O1A1Ixp33_ASAP7_75t_L g1412 ( .A1(n_1357), .A2(n_1360), .B(n_1413), .C(n_1414), .Y(n_1412) );
OR2x2_ASAP7_75t_L g1357 ( .A(n_1358), .B(n_1359), .Y(n_1357) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1359), .Y(n_1397) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1367), .Y(n_1401) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1372), .Y(n_1420) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1375), .Y(n_1411) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1384), .Y(n_1413) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
INVxp67_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
AOI211xp5_ASAP7_75t_L g1407 ( .A1(n_1408), .A2(n_1409), .B(n_1412), .C(n_1419), .Y(n_1407) );
INVxp67_ASAP7_75t_SL g1409 ( .A(n_1410), .Y(n_1409) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
CKINVDCx20_ASAP7_75t_R g1422 ( .A(n_1423), .Y(n_1422) );
CKINVDCx20_ASAP7_75t_R g1423 ( .A(n_1424), .Y(n_1423) );
INVx3_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
NAND3xp33_ASAP7_75t_L g1430 ( .A(n_1431), .B(n_1450), .C(n_1453), .Y(n_1430) );
NOR3xp33_ASAP7_75t_L g1431 ( .A(n_1432), .B(n_1443), .C(n_1449), .Y(n_1431) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_1433), .B(n_1436), .Y(n_1432) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
OR2x2_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1447), .Y(n_1444) );
INVx2_ASAP7_75t_SL g1445 ( .A(n_1446), .Y(n_1445) );
OAI21xp5_ASAP7_75t_L g1453 ( .A1(n_1454), .A2(n_1464), .B(n_1475), .Y(n_1453) );
BUFx2_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
HB1xp67_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
BUFx3_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
INVxp33_ASAP7_75t_L g1482 ( .A(n_1483), .Y(n_1482) );
INVxp33_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
NAND3xp33_ASAP7_75t_SL g1485 ( .A(n_1486), .B(n_1489), .C(n_1501), .Y(n_1485) );
NAND2xp5_ASAP7_75t_L g1490 ( .A(n_1491), .B(n_1494), .Y(n_1490) );
HB1xp67_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
endmodule