module real_jpeg_16340_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_249;
wire n_78;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_244;
wire n_213;
wire n_202;
wire n_128;
wire n_179;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_0),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_51)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_0),
.A2(n_56),
.B1(n_221),
.B2(n_224),
.Y(n_220)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_1),
.Y(n_103)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_1),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_2),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_3),
.A2(n_72),
.B1(n_75),
.B2(n_76),
.Y(n_71)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_3),
.A2(n_75),
.B1(n_175),
.B2(n_178),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_4),
.A2(n_135),
.B1(n_139),
.B2(n_140),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_4),
.Y(n_139)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_5),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_6),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_6),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_7),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_7),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_8),
.B(n_94),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_8),
.A2(n_112),
.A3(n_118),
.B1(n_120),
.B2(n_124),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_8),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_8),
.A2(n_121),
.B1(n_159),
.B2(n_163),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_8),
.A2(n_63),
.B1(n_243),
.B2(n_249),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_9),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_9),
.A2(n_46),
.B1(n_167),
.B2(n_171),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_9),
.A2(n_46),
.B1(n_244),
.B2(n_248),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_10),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_10),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_11),
.Y(n_91)
);

BUFx4f_ASAP7_75t_L g210 ( 
.A(n_11),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_184),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_182),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_109),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_15),
.B(n_109),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_62),
.C(n_92),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_16),
.A2(n_17),
.B1(n_92),
.B2(n_93),
.Y(n_215)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_41),
.B1(n_49),
.B2(n_51),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_18),
.A2(n_49),
.B1(n_51),
.B2(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_18),
.A2(n_41),
.B1(n_49),
.B2(n_213),
.Y(n_212)
);

AND2x2_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_29),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_23),
.B2(n_25),
.Y(n_19)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_22),
.Y(n_138)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_22),
.Y(n_142)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_39),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_50),
.B(n_121),
.Y(n_255)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_61),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_62),
.B(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_71),
.B1(n_78),
.B2(n_81),
.Y(n_62)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_63),
.A2(n_220),
.B1(n_243),
.B2(n_252),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g133 ( 
.A(n_64),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_64),
.Y(n_241)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_64),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_70),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_71),
.Y(n_228)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_78),
.Y(n_227)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_82),
.A2(n_131),
.B1(n_132),
.B2(n_134),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_88),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_90),
.Y(n_247)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_91),
.Y(n_226)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_95),
.A2(n_148),
.B1(n_158),
.B2(n_166),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AO21x2_ASAP7_75t_L g148 ( 
.A1(n_97),
.A2(n_124),
.B(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B1(n_104),
.B2(n_106),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_105),
.Y(n_181)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_145),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_130),
.B1(n_143),
.B2(n_144),
.Y(n_110)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_SL g213 ( 
.A1(n_118),
.A2(n_121),
.B(n_201),
.Y(n_213)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_121),
.B(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_121),
.B(n_239),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_131),
.A2(n_219),
.B1(n_227),
.B2(n_228),
.Y(n_218)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_172),
.B2(n_173),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_216),
.B(n_258),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_214),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_186),
.B(n_214),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_211),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_187),
.A2(n_211),
.B1(n_212),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_193),
.A3(n_197),
.B1(n_201),
.B2(n_206),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_207),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_231),
.B(n_257),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_229),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_229),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_250),
.B(n_256),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_242),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_255),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_255),
.Y(n_256)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);


endmodule