module fake_ibex_1215_n_1069 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_195, n_163, n_26, n_188, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1069);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1069;

wire n_599;
wire n_778;
wire n_822;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_1031;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_510;
wire n_845;
wire n_972;
wire n_947;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_991;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1018;
wire n_1044;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_280;
wire n_375;
wire n_340;
wire n_317;
wire n_708;
wire n_901;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_326;
wire n_327;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_339;
wire n_470;
wire n_276;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_1053;
wire n_343;
wire n_310;
wire n_714;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_1055;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_1025;
wire n_590;
wire n_893;
wire n_465;
wire n_1057;
wire n_1068;
wire n_325;
wire n_496;
wire n_301;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_1052;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_490;
wire n_407;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_623;
wire n_585;
wire n_1030;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_980;
wire n_454;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_968;
wire n_625;
wire n_953;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_1064;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_1028;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_1038;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_1009;
wire n_910;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1062;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_837;
wire n_797;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_1063;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_553;
wire n_554;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_567;
wire n_516;
wire n_548;
wire n_943;
wire n_1049;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_200;
wire n_564;
wire n_562;
wire n_506;
wire n_444;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_520;
wire n_411;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_1033;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_499;
wire n_227;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_379;
wire n_320;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_385;
wire n_233;
wire n_342;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_1005;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_890;
wire n_921;
wire n_912;
wire n_874;
wire n_1058;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

INVx1_ASAP7_75t_L g197 ( 
.A(n_32),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_19),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_161),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_76),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_55),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_196),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_96),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_182),
.Y(n_204)
);

NOR2xp67_ASAP7_75t_L g205 ( 
.A(n_129),
.B(n_60),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_8),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_48),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_59),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_9),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_86),
.B(n_119),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_84),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

BUFx4f_ASAP7_75t_SL g213 ( 
.A(n_139),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_124),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_68),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_42),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_156),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_102),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_11),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_115),
.B(n_167),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_64),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_114),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_47),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_93),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_91),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_75),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_31),
.Y(n_228)
);

INVxp33_ASAP7_75t_SL g229 ( 
.A(n_66),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_85),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_108),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_132),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_126),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_160),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_95),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_125),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_140),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_62),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_54),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_87),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_136),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_14),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_141),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_169),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_154),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_100),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_145),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_120),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_131),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_135),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_118),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_153),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_44),
.Y(n_258)
);

BUFx8_ASAP7_75t_SL g259 ( 
.A(n_142),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_157),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_143),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_113),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_7),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_1),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_159),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_116),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_10),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_162),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_109),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_22),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_65),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_138),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_112),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_192),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_56),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_137),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_24),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_181),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_105),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_13),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_35),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_110),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_32),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_117),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_49),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_5),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_106),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_9),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_148),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g290 ( 
.A(n_25),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_53),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_74),
.Y(n_292)
);

BUFx8_ASAP7_75t_SL g293 ( 
.A(n_19),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_104),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_35),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_83),
.B(n_146),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_77),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_173),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_71),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_166),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_149),
.Y(n_301)
);

NOR2xp67_ASAP7_75t_L g302 ( 
.A(n_51),
.B(n_2),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_69),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_42),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_107),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_82),
.Y(n_306)
);

BUFx5_ASAP7_75t_L g307 ( 
.A(n_190),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_194),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_147),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_134),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_36),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_61),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_176),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_3),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_1),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_133),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_73),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_186),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_193),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_98),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_7),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_144),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_90),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_285),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_251),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_326)
);

OA21x2_ASAP7_75t_L g327 ( 
.A1(n_218),
.A2(n_79),
.B(n_195),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_226),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_307),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_197),
.B(n_4),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_263),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_263),
.B(n_4),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_207),
.Y(n_333)
);

AND2x4_ASAP7_75t_L g334 ( 
.A(n_201),
.B(n_5),
.Y(n_334)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_209),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_226),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_307),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_307),
.B(n_6),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_200),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_203),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_208),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_212),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_198),
.B(n_6),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_214),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_307),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_206),
.Y(n_346)
);

BUFx8_ASAP7_75t_L g347 ( 
.A(n_307),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_207),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_290),
.B(n_8),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_218),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_223),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_219),
.Y(n_354)
);

AND2x4_ASAP7_75t_L g355 ( 
.A(n_201),
.B(n_11),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_267),
.Y(n_356)
);

OAI21x1_ASAP7_75t_L g357 ( 
.A1(n_223),
.A2(n_81),
.B(n_189),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_224),
.B(n_12),
.Y(n_358)
);

BUFx8_ASAP7_75t_SL g359 ( 
.A(n_267),
.Y(n_359)
);

AND2x4_ASAP7_75t_L g360 ( 
.A(n_297),
.B(n_13),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_228),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_258),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_362)
);

XNOR2x1_ASAP7_75t_L g363 ( 
.A(n_216),
.B(n_17),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_207),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_290),
.Y(n_365)
);

AND2x6_ASAP7_75t_L g366 ( 
.A(n_297),
.B(n_50),
.Y(n_366)
);

AND2x4_ASAP7_75t_L g367 ( 
.A(n_303),
.B(n_18),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_259),
.Y(n_368)
);

INVxp33_ASAP7_75t_SL g369 ( 
.A(n_247),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_259),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_255),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_277),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_227),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_283),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_215),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_295),
.Y(n_376)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_303),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_217),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_226),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_304),
.Y(n_380)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_199),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_311),
.B(n_18),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_226),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_255),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_227),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_315),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_269),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_264),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_280),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_234),
.B(n_254),
.Y(n_390)
);

BUFx8_ASAP7_75t_SL g391 ( 
.A(n_280),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_321),
.B(n_23),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_221),
.Y(n_393)
);

INVx6_ASAP7_75t_L g394 ( 
.A(n_235),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g395 ( 
.A1(n_234),
.A2(n_94),
.B(n_187),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_222),
.Y(n_396)
);

OA21x2_ASAP7_75t_L g397 ( 
.A1(n_254),
.A2(n_92),
.B(n_185),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_262),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_262),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_325),
.B(n_273),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_329),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_332),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_329),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_381),
.B(n_286),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_288),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_328),
.Y(n_407)
);

BUFx4f_ASAP7_75t_L g408 ( 
.A(n_334),
.Y(n_408)
);

AND2x6_ASAP7_75t_L g409 ( 
.A(n_334),
.B(n_230),
.Y(n_409)
);

BUFx8_ASAP7_75t_SL g410 ( 
.A(n_359),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_337),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_368),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_R g415 ( 
.A(n_370),
.B(n_269),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_381),
.B(n_274),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_328),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_366),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_351),
.Y(n_419)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_366),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_347),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_388),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_388),
.B(n_202),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_351),
.Y(n_424)
);

INVxp33_ASAP7_75t_L g425 ( 
.A(n_324),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_352),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_332),
.A2(n_229),
.B1(n_281),
.B2(n_270),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_374),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_347),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_352),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_368),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_365),
.B(n_278),
.Y(n_432)
);

AO22x2_ASAP7_75t_L g433 ( 
.A1(n_363),
.A2(n_275),
.B1(n_322),
.B2(n_238),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_365),
.B(n_289),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_346),
.B(n_354),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_349),
.B(n_313),
.Y(n_436)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_366),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_328),
.Y(n_438)
);

AND2x6_ASAP7_75t_L g439 ( 
.A(n_334),
.B(n_231),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_353),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_L g441 ( 
.A1(n_339),
.A2(n_213),
.B1(n_250),
.B2(n_252),
.Y(n_441)
);

NAND3xp33_ASAP7_75t_L g442 ( 
.A(n_350),
.B(n_360),
.C(n_355),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_SL g443 ( 
.A1(n_335),
.A2(n_288),
.B1(n_323),
.B2(n_291),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_336),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_393),
.B(n_204),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_353),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_366),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_336),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_336),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_373),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_373),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_385),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_385),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_398),
.Y(n_454)
);

AO21x2_ASAP7_75t_L g455 ( 
.A1(n_357),
.A2(n_233),
.B(n_232),
.Y(n_455)
);

BUFx10_ASAP7_75t_L g456 ( 
.A(n_355),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_350),
.B(n_316),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_335),
.Y(n_458)
);

INVxp33_ASAP7_75t_L g459 ( 
.A(n_359),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_339),
.A2(n_213),
.B1(n_268),
.B2(n_236),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_398),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_379),
.Y(n_462)
);

INVx8_ASAP7_75t_L g463 ( 
.A(n_366),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_355),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_370),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_383),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_383),
.Y(n_467)
);

INVxp33_ASAP7_75t_SL g468 ( 
.A(n_371),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_R g469 ( 
.A(n_371),
.B(n_291),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_396),
.B(n_211),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_340),
.B(n_237),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_383),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_383),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_369),
.B(n_244),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_360),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_340),
.A2(n_342),
.B1(n_375),
.B2(n_341),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_360),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_399),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_399),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_367),
.B(n_390),
.Y(n_480)
);

NAND2xp33_ASAP7_75t_R g481 ( 
.A(n_367),
.B(n_248),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_394),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_341),
.B(n_239),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_367),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_326),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_390),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_333),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_394),
.Y(n_488)
);

AND2x6_ASAP7_75t_L g489 ( 
.A(n_390),
.B(n_240),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_374),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_389),
.B(n_24),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_374),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_342),
.B(n_253),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_344),
.A2(n_378),
.B1(n_375),
.B2(n_372),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_377),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_344),
.B(n_260),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_394),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_391),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_376),
.B(n_266),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_394),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_R g501 ( 
.A(n_356),
.B(n_310),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_L g502 ( 
.A(n_378),
.B(n_220),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_380),
.B(n_241),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_333),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_480),
.A2(n_386),
.B1(n_338),
.B2(n_392),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_499),
.B(n_377),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_377),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_490),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_429),
.B(n_330),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_502),
.A2(n_310),
.B1(n_323),
.B2(n_387),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_420),
.B(n_242),
.Y(n_511)
);

OAI22xp33_ASAP7_75t_L g512 ( 
.A1(n_485),
.A2(n_384),
.B1(n_491),
.B2(n_442),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_420),
.B(n_243),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_490),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_435),
.B(n_343),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_429),
.B(n_358),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_471),
.B(n_382),
.Y(n_517)
);

NAND3xp33_ASAP7_75t_L g518 ( 
.A(n_427),
.B(n_363),
.C(n_362),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_431),
.B(n_361),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_480),
.A2(n_331),
.B1(n_395),
.B2(n_327),
.Y(n_520)
);

A2O1A1Ixp33_ASAP7_75t_L g521 ( 
.A1(n_408),
.A2(n_357),
.B(n_331),
.C(n_246),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_422),
.B(n_331),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_493),
.B(n_271),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_484),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_496),
.B(n_300),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_458),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_457),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_405),
.B(n_245),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_490),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_476),
.B(n_306),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_420),
.B(n_320),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_492),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_492),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_492),
.Y(n_534)
);

NOR3xp33_ASAP7_75t_L g535 ( 
.A(n_443),
.B(n_312),
.C(n_249),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_445),
.B(n_298),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_421),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_423),
.B(n_256),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_470),
.B(n_305),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_502),
.A2(n_319),
.B1(n_225),
.B2(n_314),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_426),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_426),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_437),
.B(n_257),
.Y(n_543)
);

AND2x6_ASAP7_75t_SL g544 ( 
.A(n_410),
.B(n_391),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_408),
.B(n_261),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_494),
.B(n_457),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_456),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_480),
.B(n_272),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_430),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_418),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_480),
.A2(n_395),
.B1(n_327),
.B2(n_397),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_428),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_480),
.A2(n_294),
.B1(n_292),
.B2(n_287),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_480),
.B(n_276),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_486),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_447),
.B(n_279),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_486),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_430),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_416),
.B(n_284),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_447),
.Y(n_560)
);

NOR3xp33_ASAP7_75t_L g561 ( 
.A(n_491),
.B(n_301),
.C(n_318),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_401),
.A2(n_395),
.B1(n_327),
.B2(n_397),
.Y(n_562)
);

AND2x6_ASAP7_75t_SL g563 ( 
.A(n_410),
.B(n_296),
.Y(n_563)
);

OAI22xp33_ASAP7_75t_L g564 ( 
.A1(n_485),
.A2(n_302),
.B1(n_309),
.B2(n_308),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_477),
.B(n_265),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_401),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_401),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_463),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_477),
.B(n_308),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_465),
.B(n_397),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_440),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_400),
.B(n_333),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_463),
.Y(n_573)
);

NOR2xp67_ASAP7_75t_L g574 ( 
.A(n_413),
.B(n_210),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_456),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_403),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_456),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_446),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_432),
.B(n_235),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_446),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_463),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_464),
.A2(n_296),
.B(n_205),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_450),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_489),
.B(n_348),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_489),
.B(n_364),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_450),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_451),
.Y(n_587)
);

NOR2xp67_ASAP7_75t_L g588 ( 
.A(n_413),
.B(n_364),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_451),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_452),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_409),
.A2(n_317),
.B1(n_299),
.B2(n_282),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_409),
.A2(n_317),
.B1(n_299),
.B2(n_282),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_464),
.B(n_317),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_452),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_464),
.B(n_317),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_436),
.Y(n_596)
);

O2A1O1Ixp33_ASAP7_75t_L g597 ( 
.A1(n_474),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_597)
);

INVxp33_ASAP7_75t_L g598 ( 
.A(n_501),
.Y(n_598)
);

AO21x1_ASAP7_75t_L g599 ( 
.A1(n_582),
.A2(n_483),
.B(n_454),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_SL g600 ( 
.A(n_526),
.B(n_468),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_515),
.B(n_527),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_561),
.A2(n_439),
.B1(n_433),
.B2(n_481),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_575),
.B(n_475),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_517),
.B(n_439),
.Y(n_604)
);

AND2x6_ASAP7_75t_SL g605 ( 
.A(n_544),
.B(n_406),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_575),
.B(n_475),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_524),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_568),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_561),
.A2(n_596),
.B1(n_512),
.B2(n_535),
.Y(n_609)
);

NOR3xp33_ASAP7_75t_L g610 ( 
.A(n_518),
.B(n_498),
.C(n_465),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_546),
.A2(n_453),
.B1(n_454),
.B2(n_461),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_568),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_511),
.A2(n_513),
.B(n_521),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_511),
.A2(n_455),
.B(n_495),
.Y(n_614)
);

AOI33xp33_ASAP7_75t_L g615 ( 
.A1(n_564),
.A2(n_460),
.A3(n_441),
.B1(n_453),
.B2(n_461),
.B3(n_479),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_522),
.B(n_433),
.Y(n_616)
);

A2O1A1Ixp33_ASAP7_75t_L g617 ( 
.A1(n_538),
.A2(n_503),
.B(n_412),
.C(n_479),
.Y(n_617)
);

O2A1O1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_512),
.A2(n_436),
.B(n_434),
.C(n_478),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_513),
.A2(n_455),
.B(n_495),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_537),
.B(n_439),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_566),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_598),
.B(n_425),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_551),
.A2(n_455),
.B(n_495),
.Y(n_623)
);

CKINVDCx6p67_ASAP7_75t_R g624 ( 
.A(n_519),
.Y(n_624)
);

NOR3xp33_ASAP7_75t_L g625 ( 
.A(n_535),
.B(n_406),
.C(n_468),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_528),
.A2(n_433),
.B1(n_402),
.B2(n_404),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_520),
.A2(n_424),
.B(n_411),
.Y(n_627)
);

NOR2x1_ASAP7_75t_L g628 ( 
.A(n_588),
.B(n_411),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_509),
.B(n_459),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_520),
.A2(n_414),
.B(n_419),
.Y(n_630)
);

BUFx8_ASAP7_75t_SL g631 ( 
.A(n_570),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_562),
.A2(n_487),
.B(n_504),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_528),
.B(n_433),
.Y(n_633)
);

AO22x1_ASAP7_75t_L g634 ( 
.A1(n_540),
.A2(n_469),
.B1(n_415),
.B2(n_299),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_524),
.Y(n_635)
);

A2O1A1Ixp33_ASAP7_75t_L g636 ( 
.A1(n_567),
.A2(n_500),
.B(n_482),
.C(n_488),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_516),
.B(n_27),
.Y(n_637)
);

NOR2x1_ASAP7_75t_L g638 ( 
.A(n_564),
.B(n_482),
.Y(n_638)
);

BUFx12f_ASAP7_75t_L g639 ( 
.A(n_563),
.Y(n_639)
);

CKINVDCx10_ASAP7_75t_R g640 ( 
.A(n_574),
.Y(n_640)
);

O2A1O1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_597),
.A2(n_565),
.B(n_569),
.C(n_548),
.Y(n_641)
);

NAND3xp33_ASAP7_75t_L g642 ( 
.A(n_505),
.B(n_235),
.C(n_282),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_559),
.B(n_28),
.Y(n_643)
);

BUFx8_ASAP7_75t_L g644 ( 
.A(n_547),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_510),
.B(n_28),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_559),
.B(n_29),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_543),
.A2(n_449),
.B(n_473),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_576),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_541),
.B(n_29),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_536),
.B(n_30),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_577),
.B(n_30),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_555),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_553),
.A2(n_497),
.B1(n_472),
.B2(n_448),
.Y(n_653)
);

A2O1A1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_580),
.A2(n_462),
.B(n_438),
.C(n_466),
.Y(n_654)
);

OAI21xp33_ASAP7_75t_L g655 ( 
.A1(n_530),
.A2(n_462),
.B(n_466),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_573),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_539),
.B(n_31),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_556),
.A2(n_448),
.B(n_438),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_506),
.B(n_33),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_507),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_542),
.B(n_33),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_579),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_557),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_549),
.B(n_34),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_523),
.B(n_525),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_558),
.Y(n_666)
);

BUFx12f_ASAP7_75t_L g667 ( 
.A(n_573),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_505),
.A2(n_497),
.B1(n_444),
.B2(n_467),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_545),
.B(n_34),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_579),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_573),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_591),
.A2(n_444),
.B1(n_467),
.B2(n_417),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_552),
.A2(n_586),
.B1(n_594),
.B2(n_587),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_589),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_L g675 ( 
.A(n_572),
.B(n_36),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_581),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_571),
.B(n_37),
.Y(n_677)
);

O2A1O1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_554),
.A2(n_578),
.B(n_590),
.C(n_583),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_591),
.A2(n_407),
.B1(n_417),
.B2(n_39),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_508),
.A2(n_407),
.B(n_121),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_534),
.B(n_38),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_514),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_592),
.A2(n_122),
.B(n_184),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_529),
.B(n_40),
.Y(n_684)
);

A2O1A1Ixp33_ASAP7_75t_L g685 ( 
.A1(n_665),
.A2(n_533),
.B(n_532),
.C(n_592),
.Y(n_685)
);

AO21x2_ASAP7_75t_L g686 ( 
.A1(n_623),
.A2(n_593),
.B(n_595),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_601),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_609),
.B(n_633),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_626),
.B(n_531),
.Y(n_689)
);

AO21x1_ASAP7_75t_L g690 ( 
.A1(n_613),
.A2(n_585),
.B(n_584),
.Y(n_690)
);

CKINVDCx16_ASAP7_75t_R g691 ( 
.A(n_600),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_644),
.Y(n_692)
);

INVxp67_ASAP7_75t_SL g693 ( 
.A(n_667),
.Y(n_693)
);

OAI21x1_ASAP7_75t_SL g694 ( 
.A1(n_683),
.A2(n_581),
.B(n_43),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_644),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_674),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_641),
.A2(n_581),
.B(n_560),
.C(n_550),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_616),
.B(n_41),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_660),
.B(n_560),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_602),
.A2(n_550),
.B1(n_43),
.B2(n_44),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_618),
.B(n_550),
.Y(n_701)
);

OAI22x1_ASAP7_75t_L g702 ( 
.A1(n_645),
.A2(n_41),
.B1(n_45),
.B2(n_46),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_615),
.B(n_45),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_611),
.B(n_46),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_611),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_666),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_624),
.A2(n_57),
.B1(n_58),
.B2(n_63),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_625),
.B(n_67),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_614),
.A2(n_70),
.B(n_72),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_622),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_627),
.A2(n_78),
.B(n_80),
.Y(n_711)
);

NOR4xp25_ASAP7_75t_L g712 ( 
.A(n_617),
.B(n_88),
.C(n_89),
.D(n_97),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_619),
.A2(n_99),
.B(n_101),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_640),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_639),
.Y(n_715)
);

OR2x6_ASAP7_75t_L g716 ( 
.A(n_634),
.B(n_103),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_650),
.B(n_123),
.Y(n_717)
);

AOI211x1_ASAP7_75t_L g718 ( 
.A1(n_599),
.A2(n_127),
.B(n_128),
.C(n_130),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_649),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_673),
.B(n_150),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_637),
.B(n_151),
.Y(n_721)
);

INVxp67_ASAP7_75t_SL g722 ( 
.A(n_631),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_604),
.A2(n_152),
.B(n_155),
.Y(n_723)
);

NAND3xp33_ASAP7_75t_L g724 ( 
.A(n_642),
.B(n_163),
.C(n_164),
.Y(n_724)
);

INVx5_ASAP7_75t_L g725 ( 
.A(n_608),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_638),
.B(n_165),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_610),
.B(n_168),
.Y(n_727)
);

AOI221x1_ASAP7_75t_L g728 ( 
.A1(n_680),
.A2(n_171),
.B1(n_172),
.B2(n_174),
.C(n_175),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_612),
.Y(n_729)
);

AO31x2_ASAP7_75t_L g730 ( 
.A1(n_630),
.A2(n_177),
.A3(n_178),
.B(n_183),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_661),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_677),
.Y(n_732)
);

OAI21xp5_ASAP7_75t_L g733 ( 
.A1(n_632),
.A2(n_678),
.B(n_659),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_681),
.A2(n_669),
.B(n_657),
.C(n_684),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_SL g735 ( 
.A1(n_683),
.A2(n_679),
.B(n_656),
.Y(n_735)
);

AOI221xp5_ASAP7_75t_L g736 ( 
.A1(n_629),
.A2(n_643),
.B1(n_646),
.B2(n_652),
.C(n_663),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_621),
.B(n_648),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_670),
.B(n_662),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_651),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_682),
.B(n_620),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_675),
.B(n_607),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_603),
.A2(n_606),
.B(n_655),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_654),
.A2(n_647),
.B(n_658),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_605),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_635),
.B(n_664),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_628),
.B(n_671),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_L g747 ( 
.A1(n_636),
.A2(n_668),
.B(n_653),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_679),
.Y(n_748)
);

BUFx8_ASAP7_75t_L g749 ( 
.A(n_676),
.Y(n_749)
);

O2A1O1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_617),
.A2(n_564),
.B(n_633),
.C(n_618),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_601),
.B(n_537),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_601),
.Y(n_752)
);

NOR2xp67_ASAP7_75t_L g753 ( 
.A(n_667),
.B(n_429),
.Y(n_753)
);

HB1xp67_ASAP7_75t_L g754 ( 
.A(n_601),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_666),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_609),
.A2(n_633),
.B1(n_602),
.B2(n_626),
.Y(n_756)
);

AO31x2_ASAP7_75t_L g757 ( 
.A1(n_599),
.A2(n_521),
.A3(n_623),
.B(n_611),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_SL g758 ( 
.A1(n_611),
.A2(n_437),
.B(n_420),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_624),
.B(n_468),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_SL g760 ( 
.A(n_600),
.B(n_410),
.Y(n_760)
);

AOI221xp5_ASAP7_75t_SL g761 ( 
.A1(n_618),
.A2(n_564),
.B1(n_512),
.B2(n_626),
.C(n_617),
.Y(n_761)
);

XNOR2xp5_ASAP7_75t_L g762 ( 
.A(n_609),
.B(n_406),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_601),
.B(n_527),
.Y(n_763)
);

OA21x2_ASAP7_75t_L g764 ( 
.A1(n_623),
.A2(n_521),
.B(n_562),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_667),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_623),
.A2(n_619),
.B(n_614),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_623),
.A2(n_619),
.B(n_614),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_L g768 ( 
.A(n_642),
.B(n_609),
.C(n_561),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_601),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_601),
.B(n_609),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_601),
.Y(n_771)
);

NAND2xp33_ASAP7_75t_L g772 ( 
.A(n_608),
.B(n_568),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_667),
.B(n_526),
.Y(n_773)
);

AO32x2_ASAP7_75t_L g774 ( 
.A1(n_611),
.A2(n_672),
.A3(n_679),
.B1(n_653),
.B2(n_599),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_601),
.B(n_527),
.Y(n_775)
);

AO21x1_ASAP7_75t_L g776 ( 
.A1(n_623),
.A2(n_613),
.B(n_680),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_665),
.A2(n_641),
.B(n_650),
.C(n_604),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_602),
.A2(n_611),
.B1(n_408),
.B2(n_609),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_623),
.A2(n_619),
.B(n_614),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_601),
.B(n_609),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_766),
.A2(n_779),
.B(n_767),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_696),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_770),
.B(n_780),
.Y(n_783)
);

OAI21x1_ASAP7_75t_SL g784 ( 
.A1(n_694),
.A2(n_778),
.B(n_707),
.Y(n_784)
);

BUFx8_ASAP7_75t_L g785 ( 
.A(n_714),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_687),
.B(n_752),
.Y(n_786)
);

CKINVDCx8_ASAP7_75t_R g787 ( 
.A(n_715),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_692),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_754),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_769),
.Y(n_790)
);

OA21x2_ASAP7_75t_L g791 ( 
.A1(n_697),
.A2(n_776),
.B(n_733),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_777),
.A2(n_743),
.B(n_734),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_695),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_688),
.A2(n_736),
.B1(n_768),
.B2(n_756),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_749),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_771),
.B(n_763),
.Y(n_796)
);

AO21x2_ASAP7_75t_L g797 ( 
.A1(n_747),
.A2(n_711),
.B(n_701),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_765),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_737),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_761),
.B(n_756),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_775),
.Y(n_801)
);

OAI21x1_ASAP7_75t_SL g802 ( 
.A1(n_707),
.A2(n_750),
.B(n_705),
.Y(n_802)
);

NAND2x1p5_ASAP7_75t_L g803 ( 
.A(n_765),
.B(n_725),
.Y(n_803)
);

BUFx2_ASAP7_75t_R g804 ( 
.A(n_744),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_765),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_751),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_751),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_719),
.Y(n_808)
);

OAI21x1_ASAP7_75t_L g809 ( 
.A1(n_764),
.A2(n_709),
.B(n_713),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_749),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_698),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_731),
.B(n_732),
.Y(n_812)
);

AO21x2_ASAP7_75t_L g813 ( 
.A1(n_735),
.A2(n_748),
.B(n_712),
.Y(n_813)
);

CKINVDCx16_ASAP7_75t_R g814 ( 
.A(n_760),
.Y(n_814)
);

INVx4_ASAP7_75t_L g815 ( 
.A(n_773),
.Y(n_815)
);

CKINVDCx8_ASAP7_75t_R g816 ( 
.A(n_691),
.Y(n_816)
);

AO31x2_ASAP7_75t_L g817 ( 
.A1(n_728),
.A2(n_690),
.A3(n_700),
.B(n_726),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_703),
.A2(n_685),
.B(n_689),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_702),
.Y(n_819)
);

OA21x2_ASAP7_75t_L g820 ( 
.A1(n_724),
.A2(n_742),
.B(n_723),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_773),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_773),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_725),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_722),
.Y(n_824)
);

INVx1_ASAP7_75t_SL g825 ( 
.A(n_725),
.Y(n_825)
);

AO31x2_ASAP7_75t_L g826 ( 
.A1(n_757),
.A2(n_720),
.A3(n_727),
.B(n_774),
.Y(n_826)
);

OA21x2_ASAP7_75t_L g827 ( 
.A1(n_704),
.A2(n_717),
.B(n_745),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_699),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_758),
.A2(n_740),
.B(n_721),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_755),
.Y(n_830)
);

OAI21x1_ASAP7_75t_SL g831 ( 
.A1(n_746),
.A2(n_738),
.B(n_741),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_729),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_706),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_708),
.Y(n_834)
);

OAI21x1_ASAP7_75t_SL g835 ( 
.A1(n_716),
.A2(n_774),
.B(n_718),
.Y(n_835)
);

AO21x2_ASAP7_75t_L g836 ( 
.A1(n_686),
.A2(n_774),
.B(n_757),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_693),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_772),
.A2(n_716),
.B(n_739),
.Y(n_838)
);

NAND3xp33_ASAP7_75t_L g839 ( 
.A(n_716),
.B(n_762),
.C(n_729),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_710),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_759),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_753),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_757),
.B(n_753),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_730),
.B(n_687),
.Y(n_844)
);

AO31x2_ASAP7_75t_L g845 ( 
.A1(n_730),
.A2(n_776),
.A3(n_767),
.B(n_766),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_763),
.B(n_775),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_749),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_766),
.A2(n_779),
.B(n_767),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_754),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_754),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_770),
.B(n_780),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_749),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_766),
.A2(n_779),
.B(n_767),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_754),
.Y(n_854)
);

INVx4_ASAP7_75t_SL g855 ( 
.A(n_765),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_754),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_754),
.B(n_687),
.Y(n_857)
);

AND2x2_ASAP7_75t_SL g858 ( 
.A(n_691),
.B(n_760),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_696),
.Y(n_859)
);

OAI21x1_ASAP7_75t_SL g860 ( 
.A1(n_694),
.A2(n_778),
.B(n_707),
.Y(n_860)
);

OAI21x1_ASAP7_75t_SL g861 ( 
.A1(n_694),
.A2(n_778),
.B(n_707),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_687),
.B(n_771),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_750),
.A2(n_777),
.B(n_768),
.C(n_736),
.Y(n_863)
);

AO31x2_ASAP7_75t_L g864 ( 
.A1(n_776),
.A2(n_767),
.A3(n_766),
.B(n_779),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_754),
.Y(n_865)
);

AO21x2_ASAP7_75t_L g866 ( 
.A1(n_781),
.A2(n_848),
.B(n_853),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_796),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_799),
.B(n_789),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_790),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_857),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_803),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_801),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_782),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_859),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_846),
.B(n_794),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_803),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_812),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_810),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_864),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_794),
.B(n_783),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_798),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_844),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_844),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_828),
.Y(n_884)
);

CKINVDCx14_ASAP7_75t_R g885 ( 
.A(n_805),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_843),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_789),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_783),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_786),
.B(n_862),
.Y(n_889)
);

OR2x2_ASAP7_75t_L g890 ( 
.A(n_851),
.B(n_800),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_865),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_851),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_795),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_800),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_865),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_786),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_862),
.B(n_840),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_808),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_849),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_850),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_854),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_856),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_830),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_819),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_806),
.B(n_807),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_863),
.B(n_834),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_833),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_795),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_831),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_847),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_863),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_792),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_811),
.B(n_841),
.Y(n_913)
);

NAND2x1_ASAP7_75t_L g914 ( 
.A(n_784),
.B(n_861),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_836),
.B(n_818),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_855),
.Y(n_916)
);

NAND2xp33_ASAP7_75t_R g917 ( 
.A(n_847),
.B(n_852),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_855),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_839),
.B(n_825),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_832),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_823),
.B(n_792),
.Y(n_921)
);

AO21x2_ASAP7_75t_L g922 ( 
.A1(n_835),
.A2(n_860),
.B(n_802),
.Y(n_922)
);

OR2x2_ASAP7_75t_L g923 ( 
.A(n_839),
.B(n_826),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_852),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_837),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_855),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_813),
.B(n_827),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_841),
.B(n_821),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_921),
.B(n_791),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_886),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_868),
.B(n_845),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_867),
.B(n_821),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_920),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_875),
.B(n_815),
.Y(n_934)
);

OAI31xp33_ASAP7_75t_L g935 ( 
.A1(n_888),
.A2(n_838),
.A3(n_822),
.B(n_788),
.Y(n_935)
);

OAI321xp33_ASAP7_75t_L g936 ( 
.A1(n_911),
.A2(n_829),
.A3(n_842),
.B1(n_841),
.B2(n_858),
.C(n_814),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_882),
.B(n_845),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_875),
.B(n_815),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_921),
.B(n_906),
.Y(n_939)
);

CKINVDCx11_ASAP7_75t_R g940 ( 
.A(n_878),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_870),
.B(n_858),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_868),
.B(n_845),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_906),
.B(n_826),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_880),
.B(n_915),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_878),
.B(n_793),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_877),
.B(n_816),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_880),
.B(n_797),
.Y(n_947)
);

OAI33xp33_ASAP7_75t_L g948 ( 
.A1(n_904),
.A2(n_824),
.A3(n_804),
.B1(n_785),
.B2(n_787),
.B3(n_817),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_915),
.B(n_827),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_919),
.B(n_817),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_925),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_911),
.A2(n_809),
.B1(n_820),
.B2(n_785),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_883),
.B(n_922),
.Y(n_953)
);

INVxp33_ASAP7_75t_L g954 ( 
.A(n_881),
.Y(n_954)
);

OR2x6_ASAP7_75t_L g955 ( 
.A(n_914),
.B(n_804),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_920),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_892),
.B(n_872),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_887),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_919),
.B(n_890),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_894),
.B(n_884),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_866),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_869),
.B(n_902),
.Y(n_962)
);

CKINVDCx6p67_ASAP7_75t_R g963 ( 
.A(n_881),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_866),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_930),
.Y(n_965)
);

INVxp67_ASAP7_75t_SL g966 ( 
.A(n_951),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_960),
.B(n_900),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_937),
.B(n_879),
.Y(n_968)
);

INVxp67_ASAP7_75t_SL g969 ( 
.A(n_933),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_930),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_933),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_959),
.B(n_923),
.Y(n_972)
);

OAI222xp33_ASAP7_75t_L g973 ( 
.A1(n_955),
.A2(n_909),
.B1(n_914),
.B2(n_923),
.C1(n_889),
.C2(n_895),
.Y(n_973)
);

CKINVDCx14_ASAP7_75t_R g974 ( 
.A(n_940),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_939),
.B(n_912),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_939),
.B(n_944),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_960),
.B(n_899),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_944),
.B(n_912),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_959),
.B(n_866),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_957),
.B(n_932),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_943),
.B(n_927),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_962),
.B(n_901),
.Y(n_982)
);

INVxp67_ASAP7_75t_SL g983 ( 
.A(n_956),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_958),
.B(n_891),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_956),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_943),
.B(n_927),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_931),
.B(n_942),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_966),
.Y(n_988)
);

AND2x2_ASAP7_75t_SL g989 ( 
.A(n_987),
.B(n_976),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_972),
.B(n_942),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_976),
.B(n_947),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_965),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_972),
.B(n_950),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_984),
.A2(n_946),
.B(n_897),
.C(n_941),
.Y(n_994)
);

OR2x6_ASAP7_75t_L g995 ( 
.A(n_971),
.B(n_955),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_965),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_981),
.B(n_929),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_970),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_981),
.B(n_929),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_967),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_SL g1001 ( 
.A(n_974),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_986),
.B(n_947),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_986),
.B(n_949),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_968),
.B(n_953),
.Y(n_1004)
);

NOR2xp67_ASAP7_75t_L g1005 ( 
.A(n_985),
.B(n_936),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_987),
.B(n_950),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_989),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_989),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_1000),
.B(n_978),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_1001),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_1002),
.B(n_978),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_988),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_992),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_1005),
.A2(n_955),
.B1(n_938),
.B2(n_934),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_996),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_998),
.Y(n_1016)
);

OAI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_995),
.A2(n_955),
.B1(n_963),
.B2(n_954),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_994),
.B(n_935),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_1003),
.B(n_975),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1003),
.B(n_975),
.Y(n_1020)
);

OAI322xp33_ASAP7_75t_L g1021 ( 
.A1(n_1018),
.A2(n_993),
.A3(n_1006),
.B1(n_990),
.B2(n_991),
.C1(n_979),
.C2(n_980),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_1007),
.A2(n_948),
.B(n_973),
.C(n_945),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_1012),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1019),
.B(n_1002),
.Y(n_1024)
);

INVxp67_ASAP7_75t_SL g1025 ( 
.A(n_1007),
.Y(n_1025)
);

AOI222xp33_ASAP7_75t_L g1026 ( 
.A1(n_1010),
.A2(n_977),
.B1(n_982),
.B2(n_997),
.C1(n_999),
.C2(n_913),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_1009),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1013),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_1008),
.A2(n_995),
.B1(n_955),
.B2(n_1004),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_1019),
.B(n_997),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1015),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1020),
.B(n_999),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_1021),
.A2(n_1017),
.B(n_1008),
.Y(n_1033)
);

AOI21xp33_ASAP7_75t_SL g1034 ( 
.A1(n_1026),
.A2(n_1014),
.B(n_917),
.Y(n_1034)
);

AOI221xp5_ASAP7_75t_L g1035 ( 
.A1(n_1025),
.A2(n_1011),
.B1(n_1020),
.B2(n_1013),
.C(n_1016),
.Y(n_1035)
);

OAI221xp5_ASAP7_75t_L g1036 ( 
.A1(n_1029),
.A2(n_1014),
.B1(n_995),
.B2(n_1006),
.C(n_993),
.Y(n_1036)
);

OAI211xp5_ASAP7_75t_L g1037 ( 
.A1(n_1022),
.A2(n_885),
.B(n_910),
.C(n_979),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_1023),
.A2(n_910),
.B(n_926),
.C(n_1004),
.Y(n_1038)
);

AOI321xp33_ASAP7_75t_L g1039 ( 
.A1(n_1030),
.A2(n_983),
.A3(n_969),
.B1(n_1004),
.B2(n_990),
.C(n_1016),
.Y(n_1039)
);

NOR3xp33_ASAP7_75t_L g1040 ( 
.A(n_1037),
.B(n_924),
.C(n_908),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1033),
.A2(n_1036),
.B1(n_1035),
.B2(n_1027),
.Y(n_1041)
);

NAND4xp25_ASAP7_75t_L g1042 ( 
.A(n_1039),
.B(n_952),
.C(n_928),
.D(n_971),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1041),
.B(n_1034),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_1040),
.A2(n_1038),
.B(n_1030),
.Y(n_1044)
);

AND2x2_ASAP7_75t_SL g1045 ( 
.A(n_1043),
.B(n_963),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_1044),
.Y(n_1046)
);

NAND3xp33_ASAP7_75t_SL g1047 ( 
.A(n_1045),
.B(n_918),
.C(n_916),
.Y(n_1047)
);

NOR2x1_ASAP7_75t_L g1048 ( 
.A(n_1045),
.B(n_1042),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1048),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_1047),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_1049),
.B(n_1046),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_SL g1052 ( 
.A1(n_1050),
.A2(n_908),
.B1(n_924),
.B2(n_893),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_SL g1053 ( 
.A1(n_1049),
.A2(n_893),
.B1(n_995),
.B2(n_871),
.Y(n_1053)
);

AO22x2_ASAP7_75t_L g1054 ( 
.A1(n_1051),
.A2(n_1032),
.B1(n_871),
.B2(n_876),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_1052),
.A2(n_1024),
.B(n_1032),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1053),
.Y(n_1056)
);

AOI22x1_ASAP7_75t_L g1057 ( 
.A1(n_1051),
.A2(n_876),
.B1(n_1028),
.B2(n_903),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_1056),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_1057),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1054),
.B(n_1031),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1054),
.A2(n_873),
.B(n_874),
.Y(n_1061)
);

OAI21xp33_ASAP7_75t_L g1062 ( 
.A1(n_1055),
.A2(n_896),
.B(n_907),
.Y(n_1062)
);

AO21x1_ASAP7_75t_SL g1063 ( 
.A1(n_1056),
.A2(n_1031),
.B(n_898),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1058),
.A2(n_922),
.B1(n_905),
.B2(n_961),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1059),
.A2(n_964),
.B1(n_961),
.B2(n_1015),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1061),
.B(n_961),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_1066),
.B(n_1062),
.Y(n_1067)
);

OA21x2_ASAP7_75t_L g1068 ( 
.A1(n_1067),
.A2(n_1060),
.B(n_1064),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1068),
.A2(n_1065),
.B1(n_1063),
.B2(n_971),
.Y(n_1069)
);


endmodule