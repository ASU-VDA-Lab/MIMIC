module real_jpeg_23765_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_354, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_354;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_323;
wire n_176;
wire n_215;
wire n_166;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_1),
.A2(n_66),
.B1(n_69),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_1),
.A2(n_29),
.B1(n_32),
.B2(n_77),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_77),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_1),
.A2(n_77),
.B1(n_92),
.B2(n_93),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g90 ( 
.A(n_4),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_5),
.A2(n_29),
.B1(n_32),
.B2(n_49),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_5),
.A2(n_49),
.B1(n_66),
.B2(n_69),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_5),
.A2(n_49),
.B1(n_83),
.B2(n_93),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_6),
.A2(n_61),
.B1(n_66),
.B2(n_69),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_6),
.A2(n_29),
.B1(n_32),
.B2(n_61),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_6),
.A2(n_61),
.B1(n_83),
.B2(n_86),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_7),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_7),
.B(n_94),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_7),
.B(n_29),
.C(n_43),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_84),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_7),
.B(n_75),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_7),
.A2(n_28),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_10),
.A2(n_80),
.B1(n_92),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_10),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_10),
.A2(n_66),
.B1(n_69),
.B2(n_97),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_97),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_10),
.A2(n_29),
.B1(n_32),
.B2(n_97),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_11),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_11),
.A2(n_68),
.B1(n_83),
.B2(n_93),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_68),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_11),
.A2(n_29),
.B1(n_32),
.B2(n_68),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_13),
.A2(n_29),
.B1(n_32),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_13),
.A2(n_39),
.B1(n_46),
.B2(n_47),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_13),
.A2(n_39),
.B1(n_66),
.B2(n_69),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_L g285 ( 
.A1(n_13),
.A2(n_39),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_14),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_14),
.A2(n_33),
.B1(n_46),
.B2(n_47),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_14),
.A2(n_33),
.B1(n_66),
.B2(n_69),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_14),
.A2(n_33),
.B1(n_80),
.B2(n_324),
.Y(n_323)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_15),
.Y(n_114)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_15),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_346),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_333),
.B(n_345),
.Y(n_17)
);

OAI321xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_299),
.A3(n_326),
.B1(n_331),
.B2(n_332),
.C(n_354),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_272),
.B(n_298),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_248),
.B(n_271),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_134),
.B(n_222),
.C(n_247),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_118),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_23),
.B(n_118),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_98),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_55),
.B2(n_56),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_25),
.B(n_56),
.C(n_98),
.Y(n_223)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_40),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_27),
.B(n_40),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B(n_34),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_28),
.A2(n_31),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_28),
.B(n_38),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_28),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_28),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_28),
.A2(n_164),
.B1(n_171),
.B2(n_177),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_28),
.A2(n_36),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_32),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g132 ( 
.A(n_30),
.Y(n_132)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_30),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_32),
.B(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_35),
.A2(n_158),
.B(n_162),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_36),
.Y(n_157)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_45),
.B(n_50),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_41),
.A2(n_53),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_41),
.A2(n_53),
.B1(n_146),
.B2(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_41),
.B(n_84),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_41),
.A2(n_45),
.B1(n_53),
.B2(n_243),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_41),
.A2(n_53),
.B(n_59),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_54)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_47),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_46),
.B(n_66),
.C(n_73),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_47),
.B(n_142),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_47),
.A2(n_72),
.B(n_189),
.C(n_190),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_50),
.B(n_212),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_52),
.A2(n_63),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_59),
.B(n_62),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_53),
.A2(n_211),
.B(n_212),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_53),
.A2(n_62),
.B(n_243),
.Y(n_256)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_64),
.C(n_78),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_57),
.A2(n_58),
.B1(n_64),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_60),
.B(n_63),
.Y(n_212)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_65),
.Y(n_127)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_69),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_66),
.A2(n_85),
.B(n_89),
.C(n_116),
.Y(n_115)
);

HAxp5_ASAP7_75t_SL g189 ( 
.A(n_66),
.B(n_84),
.CON(n_189),
.SN(n_189)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_90),
.C(n_93),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_70),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_70),
.A2(n_75),
.B1(n_126),
.B2(n_189),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_70),
.B(n_236),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_70),
.A2(n_75),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_70),
.A2(n_75),
.B(n_109),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_71),
.A2(n_107),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_71),
.A2(n_266),
.B(n_267),
.Y(n_265)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_75),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_75),
.B(n_236),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_76),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_78),
.B(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_87),
.B1(n_94),
.B2(n_95),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_84),
.B(n_85),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_83),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_84),
.B(n_177),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_91)
);

INVx11_ASAP7_75t_L g324 ( 
.A(n_86),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_87),
.A2(n_94),
.B1(n_104),
.B2(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_87),
.B(n_285),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_87),
.A2(n_94),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_87),
.A2(n_323),
.B(n_340),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_96),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_88),
.A2(n_304),
.B(n_305),
.Y(n_303)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_94),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_94),
.B(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_110),
.B2(n_117),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_101),
.B(n_105),
.C(n_117),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_102),
.A2(n_262),
.B(n_263),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_102),
.A2(n_283),
.B(n_284),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B(n_108),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_107),
.A2(n_234),
.B(n_235),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_L g308 ( 
.A1(n_107),
.A2(n_235),
.B(n_295),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_108),
.B(n_267),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_109),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_110),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_115),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_123),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_119),
.B(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_122),
.B(n_123),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.C(n_130),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_124),
.B(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_206)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_162),
.B1(n_163),
.B2(n_165),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_133),
.B(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_221),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_216),
.B(n_220),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_201),
.B(n_215),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_185),
.B(n_200),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_159),
.B(n_184),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_147),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_147),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_143),
.B1(n_144),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_154),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_149),
.B(n_152),
.C(n_154),
.Y(n_199)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_155),
.Y(n_165)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_156),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_158),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_168),
.B(n_183),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_166),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_166),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_179),
.B(n_182),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_175),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_180),
.B(n_181),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_199),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_199),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_194),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_195),
.C(n_198),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_188),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_193),
.Y(n_209)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_191),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_197),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_202),
.B(n_203),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_210),
.C(n_213),
.Y(n_219)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_219),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_224),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_246),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_237),
.B1(n_244),
.B2(n_245),
.Y(n_225)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_227),
.B(n_230),
.C(n_232),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_231),
.Y(n_262)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_244),
.C(n_246),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_242),
.Y(n_268)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_249),
.B(n_250),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_270),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_258),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_258),
.C(n_270),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_254),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_253),
.A2(n_278),
.B(n_282),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_256),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_256),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_268),
.B2(n_269),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_265),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_265),
.C(n_269),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_263),
.B(n_305),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_264),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_266),
.Y(n_293)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_268),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_273),
.B(n_274),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_297),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_289),
.B2(n_290),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_277),
.B(n_289),
.C(n_297),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_288),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_284),
.Y(n_340)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_286),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B(n_296),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_292),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_296),
.A2(n_301),
.B1(n_312),
.B2(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_314),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_300),
.B(n_314),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_312),
.C(n_313),
.Y(n_300)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_301),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_306),
.B2(n_311),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_303),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_307),
.C(n_310),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_317),
.C(n_325),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_304),
.Y(n_322)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_306),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_309),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_309),
.A2(n_310),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_309),
.B(n_319),
.C(n_321),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_325),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_321),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_327),
.B(n_328),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_335),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_343),
.B2(n_344),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_341),
.B2(n_342),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_338),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_339),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_341),
.C(n_343),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_351),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_348),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_352),
.Y(n_351)
);


endmodule