module fake_netlist_5_1079_n_27 (n_8, n_4, n_5, n_7, n_0, n_9, n_2, n_3, n_6, n_1, n_27);

input n_8;
input n_4;
input n_5;
input n_7;
input n_0;
input n_9;
input n_2;
input n_3;
input n_6;
input n_1;

output n_27;

wire n_16;
wire n_12;
wire n_25;
wire n_18;
wire n_22;
wire n_10;
wire n_24;
wire n_21;
wire n_11;
wire n_17;
wire n_19;
wire n_15;
wire n_26;
wire n_14;
wire n_23;
wire n_13;
wire n_20;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_7),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_1),
.B(n_9),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

AO21x2_ASAP7_75t_L g13 ( 
.A1(n_0),
.A2(n_3),
.B(n_5),
.Y(n_13)
);

NAND2xp33_ASAP7_75t_R g14 ( 
.A(n_4),
.B(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_2),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_6),
.B(n_3),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_12),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_17),
.B(n_14),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_19),
.B1(n_18),
.B2(n_13),
.Y(n_24)
);

AOI211xp5_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_22),
.B(n_19),
.C(n_12),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_24),
.B1(n_19),
.B2(n_13),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_26),
.B(n_2),
.Y(n_27)
);


endmodule