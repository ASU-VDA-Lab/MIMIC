module fake_jpeg_13463_n_538 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_538);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_538;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_23),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_65),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_55),
.B(n_79),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

CKINVDCx6p67_ASAP7_75t_R g117 ( 
.A(n_57),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_20),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_58),
.B(n_73),
.Y(n_145)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_61),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_66),
.Y(n_138)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_23),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_71),
.B(n_72),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_19),
.B(n_0),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_31),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_31),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g158 ( 
.A(n_84),
.Y(n_158)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_31),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_92),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_31),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_27),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_95),
.B(n_52),
.Y(n_152)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_106),
.B(n_152),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_55),
.A2(n_42),
.B1(n_32),
.B2(n_53),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_111),
.A2(n_119),
.B1(n_122),
.B2(n_40),
.Y(n_181)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_118),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_59),
.A2(n_42),
.B1(n_32),
.B2(n_53),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_63),
.A2(n_42),
.B1(n_22),
.B2(n_44),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_84),
.A2(n_68),
.B1(n_82),
.B2(n_56),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_127),
.A2(n_134),
.B1(n_155),
.B2(n_36),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_61),
.A2(n_35),
.B1(n_45),
.B2(n_19),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_77),
.Y(n_146)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_76),
.B(n_35),
.C(n_45),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_148),
.B(n_34),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_70),
.A2(n_36),
.B1(n_24),
.B2(n_44),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_78),
.B(n_40),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_83),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_60),
.A2(n_52),
.B1(n_49),
.B2(n_38),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_162),
.A2(n_99),
.B1(n_66),
.B2(n_62),
.Y(n_164)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_163),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_164),
.Y(n_242)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_85),
.B1(n_64),
.B2(n_74),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g250 ( 
.A1(n_165),
.A2(n_125),
.B1(n_121),
.B2(n_29),
.Y(n_250)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_166),
.Y(n_241)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_129),
.A2(n_101),
.B1(n_94),
.B2(n_86),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_168),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_142),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_176),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_123),
.B(n_104),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_170),
.Y(n_262)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_171),
.Y(n_247)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_174),
.Y(n_267)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_175),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_157),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_177),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_144),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_178),
.B(n_182),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_75),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_208),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_180),
.A2(n_183),
.B1(n_205),
.B2(n_34),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_181),
.A2(n_198),
.B1(n_87),
.B2(n_128),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_155),
.A2(n_162),
.B1(n_102),
.B2(n_89),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

INVx4_ASAP7_75t_SL g265 ( 
.A(n_184),
.Y(n_265)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_185),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_124),
.B(n_96),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_186),
.B(n_214),
.C(n_37),
.Y(n_251)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_107),
.Y(n_188)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_193),
.Y(n_231)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_191),
.Y(n_238)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_108),
.Y(n_192)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_192),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_140),
.B(n_80),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g252 ( 
.A(n_194),
.Y(n_252)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_195),
.Y(n_255)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_141),
.Y(n_196)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_196),
.Y(n_256)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_197),
.B(n_201),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_138),
.A2(n_90),
.B1(n_98),
.B2(n_97),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_L g199 ( 
.A1(n_145),
.A2(n_22),
.B(n_24),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_SL g233 ( 
.A(n_199),
.B(n_170),
.C(n_182),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_109),
.B(n_29),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_202),
.Y(n_239)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_110),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_141),
.Y(n_202)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_203),
.B(n_204),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_116),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_131),
.A2(n_93),
.B1(n_88),
.B2(n_103),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_206),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_114),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_207),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_117),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_117),
.B(n_100),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_210),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_137),
.B(n_28),
.Y(n_210)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_147),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_212),
.Y(n_226)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_116),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_215),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_126),
.B(n_69),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_138),
.B(n_28),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_130),
.B(n_37),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_216),
.B(n_52),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_181),
.A2(n_131),
.B1(n_151),
.B2(n_135),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_220),
.A2(n_232),
.B1(n_234),
.B2(n_240),
.Y(n_268)
);

AOI32xp33_ASAP7_75t_L g229 ( 
.A1(n_179),
.A2(n_169),
.A3(n_176),
.B1(n_172),
.B2(n_216),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_229),
.A2(n_251),
.B(n_233),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_183),
.A2(n_135),
.B1(n_151),
.B2(n_132),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_233),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_180),
.A2(n_132),
.B1(n_150),
.B2(n_154),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_170),
.B(n_174),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_236),
.B(n_248),
.C(n_266),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_165),
.A2(n_161),
.B1(n_133),
.B2(n_105),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_260),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_165),
.A2(n_133),
.B1(n_113),
.B2(n_156),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_165),
.A2(n_113),
.B1(n_156),
.B2(n_128),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_186),
.B(n_121),
.C(n_69),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_250),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_178),
.B1(n_197),
.B2(n_167),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_259),
.B(n_208),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_192),
.A2(n_52),
.B1(n_49),
.B2(n_38),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_191),
.A2(n_52),
.B1(n_49),
.B2(n_38),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_264),
.A2(n_213),
.B1(n_204),
.B2(n_188),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_186),
.B(n_57),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_270),
.A2(n_286),
.B1(n_290),
.B2(n_291),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_218),
.B(n_166),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_271),
.B(n_276),
.Y(n_323)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_267),
.Y(n_272)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_272),
.Y(n_315)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_238),
.Y(n_273)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_273),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_274),
.B(n_292),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_163),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_258),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_277),
.B(n_281),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_259),
.B(n_200),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_278),
.B(n_279),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_219),
.B(n_184),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_225),
.Y(n_280)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_280),
.Y(n_326)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_226),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_219),
.B(n_171),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_282),
.B(n_284),
.Y(n_330)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_283),
.B(n_285),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_173),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_258),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_257),
.A2(n_173),
.B1(n_212),
.B2(n_206),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_207),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_289),
.Y(n_334)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_293),
.Y(n_324)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_242),
.A2(n_188),
.B1(n_177),
.B2(n_211),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_242),
.A2(n_254),
.B1(n_222),
.B2(n_234),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_228),
.B(n_214),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_228),
.B(n_214),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_301),
.Y(n_317)
);

AND2x2_ASAP7_75t_SL g295 ( 
.A(n_266),
.B(n_194),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_295),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_254),
.A2(n_177),
.B1(n_203),
.B2(n_175),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_296),
.A2(n_302),
.B1(n_5),
.B2(n_8),
.Y(n_351)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_298),
.Y(n_344)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

NAND2xp33_ASAP7_75t_SL g346 ( 
.A(n_300),
.B(n_303),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_239),
.B(n_224),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_232),
.A2(n_201),
.B1(n_190),
.B2(n_187),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_241),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_220),
.A2(n_185),
.B1(n_217),
.B2(n_196),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_304),
.A2(n_249),
.B1(n_235),
.B2(n_223),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_231),
.A2(n_202),
.B(n_217),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_305),
.A2(n_312),
.B(n_221),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_224),
.B(n_49),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_310),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_253),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_307),
.B(n_311),
.Y(n_339)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_247),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_308),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_250),
.B(n_49),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_250),
.B(n_38),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_248),
.C(n_256),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_313),
.B(n_295),
.C(n_269),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_246),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_314),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_309),
.A2(n_250),
.B(n_261),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_SL g363 ( 
.A1(n_318),
.A2(n_319),
.B(n_321),
.C(n_342),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_309),
.A2(n_245),
.B1(n_244),
.B2(n_252),
.Y(n_319)
);

OA21x2_ASAP7_75t_L g321 ( 
.A1(n_275),
.A2(n_264),
.B(n_263),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_322),
.B(n_16),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_282),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_352),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_329),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_299),
.A2(n_263),
.B(n_265),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_331),
.A2(n_338),
.B(n_341),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_275),
.A2(n_227),
.B1(n_230),
.B2(n_243),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_332),
.A2(n_336),
.B1(n_343),
.B2(n_353),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_268),
.A2(n_227),
.B1(n_230),
.B2(n_243),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_297),
.A2(n_255),
.B(n_265),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_311),
.A2(n_241),
.B(n_195),
.Y(n_341)
);

OAI22x1_ASAP7_75t_L g342 ( 
.A1(n_268),
.A2(n_252),
.B1(n_57),
.B2(n_3),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_281),
.A2(n_252),
.B1(n_1),
.B2(n_4),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_291),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_345),
.A2(n_292),
.B(n_293),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_287),
.A2(n_277),
.B(n_285),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_347),
.A2(n_349),
.B(n_350),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_279),
.A2(n_5),
.B(n_6),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_284),
.A2(n_5),
.B(n_8),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_351),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_271),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_283),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_352),
.B(n_307),
.Y(n_354)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_354),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_356),
.B(n_365),
.C(n_380),
.Y(n_394)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_315),
.Y(n_357)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_357),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_327),
.B(n_276),
.Y(n_361)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_361),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_314),
.A2(n_270),
.B1(n_274),
.B2(n_312),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_362),
.A2(n_366),
.B1(n_370),
.B2(n_374),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_321),
.A2(n_286),
.B1(n_296),
.B2(n_302),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_364),
.A2(n_379),
.B1(n_384),
.B2(n_351),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_313),
.B(n_295),
.C(n_294),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_314),
.A2(n_319),
.B1(n_337),
.B2(n_318),
.Y(n_366)
);

AOI21xp33_ASAP7_75t_SL g368 ( 
.A1(n_338),
.A2(n_295),
.B(n_305),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_368),
.B(n_372),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_337),
.A2(n_288),
.B1(n_301),
.B2(n_304),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_371),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_317),
.B(n_278),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_315),
.Y(n_373)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_373),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_333),
.A2(n_306),
.B1(n_272),
.B2(n_273),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_334),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_378),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_330),
.A2(n_290),
.B1(n_303),
.B2(n_300),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_376),
.A2(n_382),
.B1(n_383),
.B2(n_389),
.Y(n_392)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_316),
.Y(n_377)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_377),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_334),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_321),
.A2(n_298),
.B1(n_308),
.B2(n_289),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_313),
.B(n_9),
.C(n_10),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_381),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_330),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_333),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_321),
.A2(n_18),
.B1(n_14),
.B2(n_15),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_347),
.A2(n_13),
.B(n_15),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_386),
.B(n_387),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_328),
.B(n_16),
.Y(n_387)
);

NOR2x1_ASAP7_75t_L g388 ( 
.A(n_339),
.B(n_16),
.Y(n_388)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_388),
.Y(n_413)
);

OAI22x1_ASAP7_75t_SL g389 ( 
.A1(n_342),
.A2(n_18),
.B1(n_341),
.B2(n_339),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_365),
.B(n_317),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_393),
.B(n_395),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_356),
.B(n_322),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_359),
.B(n_354),
.C(n_361),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_396),
.B(n_407),
.C(n_408),
.Y(n_435)
);

XNOR2x1_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_328),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_325),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_366),
.A2(n_324),
.B1(n_340),
.B2(n_332),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_401),
.A2(n_364),
.B1(n_379),
.B2(n_360),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_357),
.Y(n_405)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_405),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_367),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_406),
.B(n_410),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_359),
.B(n_331),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_323),
.C(n_348),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_348),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_409),
.B(n_411),
.C(n_349),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_375),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_370),
.B(n_335),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_414),
.A2(n_418),
.B1(n_420),
.B2(n_343),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_355),
.A2(n_324),
.B1(n_336),
.B2(n_340),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_416),
.A2(n_417),
.B1(n_358),
.B2(n_384),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_355),
.A2(n_324),
.B1(n_323),
.B2(n_329),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_360),
.A2(n_345),
.B1(n_335),
.B2(n_324),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_360),
.A2(n_325),
.B1(n_342),
.B2(n_316),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_422),
.A2(n_427),
.B1(n_404),
.B2(n_363),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_423),
.B(n_426),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_402),
.A2(n_388),
.B(n_369),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_424),
.A2(n_415),
.B(n_388),
.Y(n_457)
);

FAx1_ASAP7_75t_SL g425 ( 
.A(n_396),
.B(n_369),
.CI(n_378),
.CON(n_425),
.SN(n_425)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_425),
.B(n_440),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_393),
.B(n_371),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_416),
.Y(n_429)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_429),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_391),
.A2(n_358),
.B1(n_387),
.B2(n_386),
.Y(n_430)
);

AOI322xp5_ASAP7_75t_L g460 ( 
.A1(n_430),
.A2(n_414),
.A3(n_418),
.B1(n_420),
.B2(n_419),
.C1(n_415),
.C2(n_413),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_390),
.B(n_326),
.Y(n_431)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_431),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_411),
.Y(n_432)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_432),
.Y(n_454)
);

A2O1A1Ixp33_ASAP7_75t_SL g433 ( 
.A1(n_401),
.A2(n_363),
.B(n_389),
.C(n_385),
.Y(n_433)
);

BUFx12_ASAP7_75t_L g468 ( 
.A(n_433),
.Y(n_468)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_434),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_395),
.B(n_346),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_436),
.B(n_437),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_346),
.Y(n_437)
);

XOR2x1_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_363),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_439),
.B(n_445),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_399),
.B(n_326),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_405),
.Y(n_441)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_441),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_403),
.Y(n_442)
);

INVx11_ASAP7_75t_L g461 ( 
.A(n_442),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_400),
.B(n_382),
.Y(n_443)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_443),
.Y(n_470)
);

NAND2xp33_ASAP7_75t_SL g445 ( 
.A(n_402),
.B(n_350),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_409),
.B(n_376),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_446),
.B(n_448),
.C(n_394),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_344),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_447),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_453),
.B(n_437),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_457),
.A2(n_424),
.B(n_452),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_394),
.C(n_408),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_458),
.B(n_460),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_428),
.Y(n_459)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_459),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_435),
.B(n_444),
.C(n_426),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_462),
.B(n_467),
.C(n_449),
.Y(n_472)
);

AOI322xp5_ASAP7_75t_L g463 ( 
.A1(n_429),
.A2(n_397),
.A3(n_391),
.B1(n_363),
.B2(n_417),
.C1(n_392),
.C2(n_403),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_463),
.B(n_434),
.Y(n_477)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_466),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_363),
.C(n_405),
.Y(n_467)
);

NOR2xp67_ASAP7_75t_SL g488 ( 
.A(n_472),
.B(n_478),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_458),
.B(n_446),
.C(n_439),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_474),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_436),
.C(n_448),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_461),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_475),
.B(n_476),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_461),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_477),
.A2(n_456),
.B1(n_466),
.B2(n_450),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_453),
.B(n_423),
.C(n_438),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_465),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_459),
.B(n_425),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_480),
.A2(n_481),
.B(n_468),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_449),
.B(n_433),
.C(n_425),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_482),
.B(n_454),
.C(n_456),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_469),
.A2(n_433),
.B(n_392),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_483),
.A2(n_485),
.B(n_452),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_450),
.A2(n_433),
.B(n_421),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_467),
.B(n_373),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_454),
.Y(n_497)
);

AOI21x1_ASAP7_75t_L g507 ( 
.A1(n_489),
.A2(n_491),
.B(n_473),
.Y(n_507)
);

NOR2xp67_ASAP7_75t_L g491 ( 
.A(n_478),
.B(n_455),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_492),
.B(n_498),
.Y(n_513)
);

INVx11_ASAP7_75t_L g493 ( 
.A(n_483),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_493),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_495),
.A2(n_493),
.B1(n_502),
.B2(n_503),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_487),
.B(n_465),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_502),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_470),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_459),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_472),
.B(n_451),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_499),
.B(n_501),
.Y(n_514)
);

OAI21xp33_ASAP7_75t_SL g506 ( 
.A1(n_500),
.A2(n_484),
.B(n_468),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_471),
.B(n_464),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_485),
.B(n_464),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_503),
.A2(n_481),
.B(n_482),
.Y(n_504)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_504),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_479),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_505),
.B(n_509),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_507),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_488),
.A2(n_474),
.B(n_457),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_508),
.A2(n_500),
.B(n_496),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_495),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_451),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_510),
.B(n_377),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_511),
.B(n_515),
.Y(n_522)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_518),
.Y(n_526)
);

INVx6_ASAP7_75t_L g519 ( 
.A(n_513),
.Y(n_519)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_519),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_516),
.A2(n_501),
.B(n_497),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_521),
.B(n_524),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_509),
.A2(n_468),
.B1(n_470),
.B2(n_404),
.Y(n_524)
);

NOR2xp67_ASAP7_75t_SL g528 ( 
.A(n_525),
.B(n_514),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_528),
.B(n_529),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_520),
.B(n_516),
.C(n_512),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_526),
.B(n_517),
.C(n_523),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_531),
.Y(n_535)
);

AOI321xp33_ASAP7_75t_L g533 ( 
.A1(n_530),
.A2(n_522),
.A3(n_519),
.B1(n_527),
.B2(n_506),
.C(n_468),
.Y(n_533)
);

OAI321xp33_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_522),
.A3(n_320),
.B1(n_383),
.B2(n_353),
.C(n_18),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_534),
.B(n_532),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_535),
.B(n_320),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_18),
.Y(n_538)
);


endmodule