module fake_netlist_6_2887_n_2124 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2124);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2124;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_1094;
wire n_953;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_SL g211 ( 
.A(n_84),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_165),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_40),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_48),
.Y(n_214)
);

CKINVDCx11_ASAP7_75t_R g215 ( 
.A(n_154),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_78),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g217 ( 
.A(n_140),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_23),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_147),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_34),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_14),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_69),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_35),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_26),
.Y(n_226)
);

BUFx2_ASAP7_75t_SL g227 ( 
.A(n_124),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_91),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_131),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_39),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_158),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_27),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_8),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_16),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_62),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_203),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_178),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_81),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_126),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_51),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_208),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_51),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_49),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_105),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_89),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_92),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_37),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_188),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_152),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_73),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_111),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_200),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_78),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_31),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_189),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_160),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_72),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_0),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_88),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_85),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_162),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_157),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_142),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_101),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_29),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_77),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_167),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_50),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_172),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_103),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_132),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_113),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_185),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_37),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_79),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_148),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_117),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_45),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_195),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_18),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_125),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_2),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_7),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_151),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_38),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_41),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_11),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_25),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_55),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_53),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_74),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_10),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_41),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_204),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_76),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_79),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_8),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_71),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_64),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_170),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_179),
.Y(n_302)
);

BUFx2_ASAP7_75t_SL g303 ( 
.A(n_12),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_61),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_55),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_66),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_9),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_95),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_168),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_82),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_197),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_97),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_169),
.Y(n_313)
);

BUFx8_ASAP7_75t_SL g314 ( 
.A(n_199),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_138),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_50),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_128),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_133),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_1),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_59),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_164),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_16),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_7),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_29),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_210),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_144),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_52),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_191),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_67),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_61),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_54),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_0),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_80),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_98),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_4),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_119),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_100),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_75),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_32),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_28),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_171),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_36),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_43),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_77),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g345 ( 
.A(n_86),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_10),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_42),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_127),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_122),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_143),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_110),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_175),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_68),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_130),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_107),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_74),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_161),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_104),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_68),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_129),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_99),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_4),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_35),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_166),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_12),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_202),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_19),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_6),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_75),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_181),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_66),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_27),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_60),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_123),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_65),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_6),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_156),
.Y(n_377)
);

BUFx8_ASAP7_75t_SL g378 ( 
.A(n_205),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_54),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_53),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_2),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_108),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_187),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_15),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_116),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_72),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_137),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_136),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_139),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_52),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_135),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_57),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_38),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_94),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_149),
.Y(n_395)
);

BUFx5_ASAP7_75t_L g396 ( 
.A(n_150),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_141),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_121),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_62),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_201),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_23),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_87),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_14),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_36),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_186),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_11),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_42),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_20),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_18),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_159),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_109),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_20),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_32),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_71),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_26),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_114),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_49),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_184),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_90),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_341),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_292),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_221),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_212),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_268),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_341),
.B(n_1),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_347),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_221),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_239),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_239),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_218),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_278),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_317),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_347),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_259),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_398),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_314),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_292),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_378),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_292),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_292),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_213),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_259),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_211),
.B(n_3),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_292),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_215),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_292),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_376),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_237),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_376),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_214),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_237),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_251),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_R g453 ( 
.A(n_244),
.B(n_83),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_251),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_255),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_255),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_216),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_222),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_376),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_261),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_261),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_226),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_218),
.B(n_3),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_264),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_264),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_389),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_302),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_302),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_276),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_376),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_211),
.B(n_231),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_308),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_230),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_R g474 ( 
.A(n_419),
.B(n_5),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_308),
.Y(n_475)
);

INVxp33_ASAP7_75t_SL g476 ( 
.A(n_303),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_312),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_312),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_318),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_233),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_242),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_318),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_389),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_303),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_326),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_376),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_219),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_220),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_326),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_228),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_334),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_334),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_337),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_243),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_229),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_236),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_247),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_337),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_349),
.B(n_5),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_412),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g501 ( 
.A(n_348),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_238),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_217),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_245),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_348),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_250),
.Y(n_506)
);

CKINVDCx14_ASAP7_75t_R g507 ( 
.A(n_217),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_246),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_349),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_253),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_248),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_257),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_258),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_266),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_412),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_350),
.B(n_355),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_412),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_412),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_252),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_260),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_350),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_355),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_364),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_267),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_262),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_364),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_265),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_234),
.B(n_9),
.Y(n_528)
);

OR2x6_ASAP7_75t_L g529 ( 
.A(n_425),
.B(n_227),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_516),
.B(n_412),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_449),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_449),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_459),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_459),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_486),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_447),
.Y(n_536)
);

NOR2x1_ASAP7_75t_L g537 ( 
.A(n_471),
.B(n_227),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_486),
.Y(n_538)
);

AND2x6_ASAP7_75t_L g539 ( 
.A(n_463),
.B(n_357),
.Y(n_539)
);

CKINVDCx8_ASAP7_75t_R g540 ( 
.A(n_503),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_434),
.B(n_270),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_442),
.B(n_418),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_500),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_447),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_500),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_501),
.B(n_366),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_515),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_470),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_515),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_505),
.B(n_366),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_517),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_517),
.Y(n_552)
);

OA21x2_ASAP7_75t_L g553 ( 
.A1(n_421),
.A2(n_383),
.B(n_374),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_443),
.B(n_271),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_470),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_421),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_437),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_518),
.B(n_273),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_518),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_437),
.B(n_231),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_439),
.B(n_274),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_439),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_440),
.B(n_277),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_440),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_444),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_444),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_446),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_446),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_422),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_427),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_428),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_429),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_452),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_454),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_455),
.Y(n_575)
);

BUFx8_ASAP7_75t_L g576 ( 
.A(n_463),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_448),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_456),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_430),
.A2(n_223),
.B1(n_281),
.B2(n_235),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_460),
.B(n_280),
.Y(n_580)
);

CKINVDCx14_ASAP7_75t_R g581 ( 
.A(n_507),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_461),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_464),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_465),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_467),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_473),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_468),
.B(n_282),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_472),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_475),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_477),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_478),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_479),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_482),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_485),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_489),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_484),
.B(n_234),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_491),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_528),
.B(n_374),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_492),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_493),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_498),
.B(n_285),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_509),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_521),
.B(n_301),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_522),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_523),
.B(n_526),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_528),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_499),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_469),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_420),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_476),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_441),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_441),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_476),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_450),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_453),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_562),
.Y(n_616)
);

NAND2xp33_ASAP7_75t_L g617 ( 
.A(n_607),
.B(n_450),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_568),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_536),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_613),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_581),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_568),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_599),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_606),
.B(n_457),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_599),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_615),
.B(n_457),
.Y(n_626)
);

AO21x2_ASAP7_75t_L g627 ( 
.A1(n_554),
.A2(n_387),
.B(n_383),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_568),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_536),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_615),
.B(n_487),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_612),
.B(n_614),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_599),
.Y(n_632)
);

AND2x6_ASAP7_75t_L g633 ( 
.A(n_598),
.B(n_249),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_574),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_607),
.A2(n_550),
.B1(n_546),
.B2(n_598),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_536),
.Y(n_636)
);

NAND3xp33_ASAP7_75t_L g637 ( 
.A(n_607),
.B(n_395),
.C(n_387),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_607),
.A2(n_353),
.B1(n_283),
.B2(n_294),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_606),
.B(n_458),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_599),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_606),
.B(n_458),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_599),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_608),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_612),
.B(n_462),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_544),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_562),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_607),
.A2(n_490),
.B1(n_495),
.B2(n_488),
.Y(n_647)
);

INVxp67_ASAP7_75t_SL g648 ( 
.A(n_558),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_571),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_602),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_612),
.B(n_462),
.Y(n_651)
);

AOI22x1_ASAP7_75t_L g652 ( 
.A1(n_598),
.A2(n_353),
.B1(n_481),
.B2(n_480),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_571),
.B(n_395),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_602),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_612),
.B(n_614),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_602),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_607),
.B(n_480),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_541),
.B(n_496),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_568),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_607),
.B(n_481),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_546),
.B(n_494),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_568),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_568),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_571),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_541),
.B(n_494),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_544),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_544),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_542),
.B(n_502),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_556),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_612),
.B(n_497),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_556),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_613),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_546),
.A2(n_283),
.B1(n_294),
.B2(n_232),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_542),
.B(n_497),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_568),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_550),
.A2(n_381),
.B1(n_414),
.B2(n_232),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_555),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_602),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_602),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_555),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_613),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_612),
.B(n_506),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_612),
.B(n_506),
.Y(n_683)
);

BUFx4f_ASAP7_75t_L g684 ( 
.A(n_553),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_571),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_L g686 ( 
.A(n_550),
.B(n_263),
.C(n_249),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_574),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_613),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_611),
.B(n_504),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_614),
.B(n_510),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_555),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_555),
.Y(n_692)
);

INVx5_ASAP7_75t_L g693 ( 
.A(n_539),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_555),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_556),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_555),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_572),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_572),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_557),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_L g700 ( 
.A(n_539),
.B(n_510),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_554),
.B(n_537),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_R g702 ( 
.A(n_581),
.B(n_508),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_572),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_596),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_537),
.B(n_512),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_SL g706 ( 
.A(n_610),
.B(n_451),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_555),
.Y(n_707)
);

NAND2xp33_ASAP7_75t_SL g708 ( 
.A(n_610),
.B(n_466),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_572),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_557),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_600),
.Y(n_711)
);

OAI21xp33_ASAP7_75t_SL g712 ( 
.A1(n_529),
.A2(n_225),
.B(n_224),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_600),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_614),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_557),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_561),
.B(n_512),
.Y(n_716)
);

AND2x6_ASAP7_75t_L g717 ( 
.A(n_611),
.B(n_263),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_614),
.B(n_513),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_611),
.B(n_511),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_574),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_540),
.Y(n_721)
);

AND2x2_ASAP7_75t_SL g722 ( 
.A(n_553),
.B(n_295),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_596),
.Y(n_723)
);

NOR3xp33_ASAP7_75t_L g724 ( 
.A(n_579),
.B(n_586),
.C(n_433),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_605),
.B(n_513),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_562),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_600),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_539),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_562),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_609),
.B(n_519),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_609),
.B(n_520),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_600),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_529),
.A2(n_539),
.B1(n_576),
.B2(n_530),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_564),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_561),
.B(n_514),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_564),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_586),
.Y(n_737)
);

BUFx4f_ASAP7_75t_L g738 ( 
.A(n_553),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_564),
.Y(n_739)
);

NOR2x1p5_ASAP7_75t_L g740 ( 
.A(n_614),
.B(n_426),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_567),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_565),
.Y(n_742)
);

INVx5_ASAP7_75t_L g743 ( 
.A(n_539),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_565),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_566),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_605),
.B(n_295),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_605),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_567),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_563),
.B(n_514),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_567),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_605),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_566),
.Y(n_752)
);

INVx4_ASAP7_75t_L g753 ( 
.A(n_539),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_563),
.B(n_524),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_570),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_614),
.B(n_524),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_531),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_531),
.Y(n_758)
);

AND2x2_ASAP7_75t_SL g759 ( 
.A(n_553),
.B(n_315),
.Y(n_759)
);

OR2x6_ASAP7_75t_L g760 ( 
.A(n_529),
.B(n_315),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_577),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_570),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_L g763 ( 
.A(n_530),
.B(n_474),
.C(n_414),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_558),
.B(n_241),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_580),
.B(n_525),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_580),
.B(n_256),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_548),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_587),
.B(n_527),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_755),
.Y(n_769)
);

INVxp33_ASAP7_75t_L g770 ( 
.A(n_661),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_755),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_648),
.B(n_576),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_635),
.B(n_576),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_657),
.B(n_576),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_762),
.Y(n_775)
);

O2A1O1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_639),
.A2(n_601),
.B(n_603),
.C(n_587),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_762),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_660),
.B(n_576),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_701),
.B(n_601),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_764),
.B(n_603),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_766),
.B(n_539),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_747),
.Y(n_782)
);

OAI22xp33_ASAP7_75t_L g783 ( 
.A1(n_665),
.A2(n_529),
.B1(n_540),
.B2(n_433),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_685),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_685),
.B(n_539),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_684),
.A2(n_560),
.B(n_605),
.Y(n_786)
);

NAND3xp33_ASAP7_75t_L g787 ( 
.A(n_763),
.B(n_652),
.C(n_641),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_728),
.B(n_540),
.Y(n_788)
);

BUFx6f_ASAP7_75t_SL g789 ( 
.A(n_704),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_697),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_624),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_681),
.Y(n_792)
);

NOR2xp67_ASAP7_75t_SL g793 ( 
.A(n_693),
.B(n_357),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_643),
.B(n_608),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_757),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_697),
.B(n_539),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_698),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_704),
.B(n_608),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_633),
.B(n_539),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_723),
.B(n_596),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_698),
.B(n_529),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_716),
.B(n_529),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_723),
.B(n_426),
.Y(n_803)
);

NOR2xp67_ASAP7_75t_L g804 ( 
.A(n_647),
.B(n_575),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_735),
.B(n_483),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_728),
.B(n_753),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_749),
.B(n_575),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_703),
.B(n_574),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_754),
.B(n_582),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_703),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_747),
.B(n_582),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_757),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_722),
.A2(n_759),
.B1(n_627),
.B2(n_633),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_709),
.B(n_574),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_709),
.B(n_574),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_713),
.B(n_574),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_713),
.B(n_578),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_674),
.B(n_584),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_758),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_L g820 ( 
.A(n_633),
.B(n_396),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_681),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_761),
.B(n_577),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_624),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_727),
.B(n_578),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_617),
.A2(n_668),
.B1(n_658),
.B2(n_765),
.Y(n_825)
);

AOI221xp5_ASAP7_75t_L g826 ( 
.A1(n_724),
.A2(n_579),
.B1(n_363),
.B2(n_322),
.C(n_286),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_661),
.B(n_423),
.Y(n_827)
);

NOR3xp33_ASAP7_75t_L g828 ( 
.A(n_730),
.B(n_585),
.C(n_584),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_727),
.Y(n_829)
);

NAND2xp33_ASAP7_75t_L g830 ( 
.A(n_633),
.B(n_396),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_732),
.B(n_578),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_728),
.B(n_357),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_732),
.B(n_578),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_747),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_728),
.B(n_357),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_751),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_751),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_746),
.B(n_578),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_737),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_742),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_768),
.A2(n_431),
.B1(n_432),
.B2(n_424),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_746),
.B(n_578),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_751),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_742),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_620),
.B(n_585),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_744),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_649),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_649),
.Y(n_848)
);

BUFx6f_ASAP7_75t_SL g849 ( 
.A(n_653),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_746),
.B(n_578),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_620),
.B(n_589),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_746),
.B(n_590),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_722),
.B(n_590),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_744),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_722),
.B(n_590),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_759),
.B(n_590),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_672),
.B(n_589),
.Y(n_857)
);

BUFx8_ASAP7_75t_L g858 ( 
.A(n_725),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_702),
.Y(n_859)
);

O2A1O1Ixp5_ASAP7_75t_L g860 ( 
.A1(n_684),
.A2(n_560),
.B(n_591),
.C(n_588),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_745),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_745),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_649),
.B(n_592),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_753),
.B(n_357),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_664),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_753),
.B(n_396),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_753),
.B(n_396),
.Y(n_867)
);

AND2x6_ASAP7_75t_SL g868 ( 
.A(n_630),
.B(n_224),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_759),
.B(n_590),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_664),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_752),
.B(n_590),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_641),
.Y(n_872)
);

NOR3xp33_ASAP7_75t_L g873 ( 
.A(n_731),
.B(n_593),
.C(n_592),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_752),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_693),
.B(n_396),
.Y(n_875)
);

OAI21xp33_ASAP7_75t_L g876 ( 
.A1(n_673),
.A2(n_594),
.B(n_593),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_627),
.A2(n_553),
.B1(n_381),
.B2(n_225),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_664),
.B(n_590),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_672),
.B(n_594),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_711),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_689),
.B(n_435),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_712),
.A2(n_604),
.B(n_597),
.C(n_583),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_619),
.Y(n_883)
);

NOR2xp67_ASAP7_75t_L g884 ( 
.A(n_621),
.B(n_569),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_725),
.Y(n_885)
);

OAI22xp33_ASAP7_75t_L g886 ( 
.A1(n_760),
.A2(n_333),
.B1(n_400),
.B2(n_445),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_733),
.A2(n_688),
.B1(n_631),
.B2(n_655),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_619),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_688),
.B(n_595),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_711),
.B(n_595),
.Y(n_890)
);

BUFx6f_ASAP7_75t_SL g891 ( 
.A(n_653),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_693),
.B(n_396),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_711),
.B(n_595),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_629),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_629),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_653),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_721),
.Y(n_897)
);

NAND3xp33_ASAP7_75t_SL g898 ( 
.A(n_719),
.B(n_438),
.C(n_436),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_626),
.B(n_275),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_705),
.B(n_595),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_627),
.B(n_595),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_636),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_636),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_633),
.A2(n_356),
.B1(n_240),
.B2(n_254),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_717),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_623),
.B(n_595),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_645),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_645),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_740),
.B(n_569),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_763),
.B(n_595),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_693),
.B(n_396),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_666),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_623),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_712),
.A2(n_403),
.B(n_254),
.C(n_269),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_625),
.B(n_588),
.Y(n_915)
);

OR2x6_ASAP7_75t_L g916 ( 
.A(n_760),
.B(n_240),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_625),
.B(n_588),
.Y(n_917)
);

NAND2xp33_ASAP7_75t_L g918 ( 
.A(n_633),
.B(n_396),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_666),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_632),
.B(n_588),
.Y(n_920)
);

AND2x6_ASAP7_75t_SL g921 ( 
.A(n_760),
.B(n_269),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_SL g922 ( 
.A1(n_652),
.A2(n_306),
.B1(n_316),
.B2(n_359),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_632),
.B(n_591),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_693),
.B(n_396),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_653),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_740),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_693),
.B(n_560),
.Y(n_927)
);

NAND2x1_ASAP7_75t_L g928 ( 
.A(n_633),
.B(n_677),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_640),
.Y(n_929)
);

NAND3xp33_ASAP7_75t_L g930 ( 
.A(n_676),
.B(n_284),
.C(n_279),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_640),
.B(n_591),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_642),
.B(n_591),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_642),
.Y(n_933)
);

BUFx5_ASAP7_75t_L g934 ( 
.A(n_714),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_650),
.B(n_560),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_650),
.B(n_560),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_644),
.B(n_287),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_654),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_654),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_656),
.B(n_532),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_840),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_825),
.A2(n_738),
.B(n_684),
.C(n_686),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_802),
.A2(n_738),
.B(n_684),
.C(n_686),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_860),
.A2(n_738),
.B(n_637),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_780),
.B(n_651),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_840),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_802),
.A2(n_738),
.B(n_682),
.C(n_683),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_853),
.A2(n_637),
.B(n_700),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_779),
.B(n_714),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_846),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_846),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_776),
.A2(n_670),
.B(n_718),
.C(n_690),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_854),
.Y(n_953)
);

INVx4_ASAP7_75t_L g954 ( 
.A(n_847),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_791),
.B(n_714),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_806),
.A2(n_743),
.B(n_622),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_818),
.B(n_714),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_818),
.B(n_756),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_855),
.A2(n_743),
.B(n_622),
.Y(n_959)
);

AOI222xp33_ASAP7_75t_L g960 ( 
.A1(n_826),
.A2(n_407),
.B1(n_706),
.B2(n_708),
.C1(n_379),
.C2(n_289),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_807),
.B(n_809),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_807),
.A2(n_678),
.B(n_679),
.C(n_656),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_856),
.A2(n_869),
.B(n_786),
.Y(n_963)
);

OAI321xp33_ASAP7_75t_L g964 ( 
.A1(n_937),
.A2(n_393),
.A3(n_403),
.B1(n_384),
.B2(n_406),
.C(n_380),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_889),
.A2(n_743),
.B(n_622),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_823),
.B(n_743),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_770),
.B(n_760),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_889),
.A2(n_842),
.B(n_838),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_858),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_850),
.A2(n_743),
.B(n_659),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_852),
.A2(n_659),
.B(n_618),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_870),
.A2(n_659),
.B(n_618),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_809),
.B(n_678),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_845),
.B(n_679),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_870),
.A2(n_659),
.B(n_618),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_878),
.A2(n_662),
.B(n_618),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_787),
.A2(n_760),
.B1(n_717),
.B2(n_638),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_854),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_890),
.A2(n_675),
.B(n_662),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_893),
.A2(n_675),
.B(n_662),
.Y(n_980)
);

OR2x6_ASAP7_75t_L g981 ( 
.A(n_822),
.B(n_916),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_798),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_872),
.B(n_634),
.Y(n_983)
);

NOR2xp67_ASAP7_75t_L g984 ( 
.A(n_839),
.B(n_767),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_845),
.B(n_717),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_851),
.B(n_717),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_910),
.A2(n_646),
.B(n_616),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_914),
.A2(n_573),
.B(n_583),
.C(n_569),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_910),
.A2(n_646),
.B(n_616),
.Y(n_989)
);

OAI321xp33_ASAP7_75t_L g990 ( 
.A1(n_937),
.A2(n_342),
.A3(n_330),
.B1(n_324),
.B2(n_323),
.C(n_304),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_770),
.B(n_290),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_934),
.A2(n_675),
.B(n_662),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_934),
.A2(n_675),
.B(n_634),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_800),
.B(n_573),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_934),
.A2(n_687),
.B(n_634),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_934),
.A2(n_687),
.B(n_634),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_792),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_934),
.B(n_634),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_861),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_934),
.A2(n_687),
.B(n_634),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_900),
.A2(n_720),
.B(n_687),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_900),
.A2(n_720),
.B(n_687),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_794),
.B(n_573),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_803),
.B(n_583),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_896),
.A2(n_720),
.B(n_687),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_885),
.B(n_720),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_861),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_913),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_821),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_925),
.A2(n_720),
.B(n_680),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_851),
.B(n_857),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_857),
.B(n_717),
.Y(n_1012)
);

AO21x2_ASAP7_75t_L g1013 ( 
.A1(n_901),
.A2(n_671),
.B(n_669),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_914),
.A2(n_604),
.B(n_597),
.C(n_533),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_827),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_804),
.A2(n_879),
.B(n_813),
.C(n_805),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_781),
.A2(n_720),
.B(n_680),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_879),
.B(n_717),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_929),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_773),
.A2(n_604),
.B(n_597),
.C(n_543),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_811),
.B(n_309),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_847),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_887),
.A2(n_680),
.B(n_677),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_811),
.Y(n_1024)
);

CKINVDCx10_ASAP7_75t_R g1025 ( 
.A(n_789),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_813),
.A2(n_767),
.B1(n_677),
.B2(n_680),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_785),
.A2(n_691),
.B(n_677),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_805),
.B(n_291),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_769),
.B(n_717),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_771),
.B(n_628),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_847),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_796),
.A2(n_692),
.B(n_691),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_799),
.A2(n_692),
.B(n_691),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_775),
.B(n_777),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_844),
.B(n_628),
.Y(n_1035)
);

AOI21x1_ASAP7_75t_L g1036 ( 
.A1(n_866),
.A2(n_867),
.B(n_835),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_862),
.B(n_628),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_874),
.B(n_628),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_935),
.A2(n_692),
.B(n_691),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_811),
.B(n_663),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_847),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_795),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_863),
.B(n_663),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_936),
.A2(n_801),
.B(n_832),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_881),
.B(n_293),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_933),
.Y(n_1046)
);

BUFx4f_ASAP7_75t_L g1047 ( 
.A(n_916),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_772),
.B(n_310),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_863),
.B(n_663),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_832),
.A2(n_646),
.B(n_616),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_835),
.A2(n_694),
.B(n_692),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_863),
.B(n_663),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_828),
.B(n_873),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_864),
.A2(n_729),
.B(n_726),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_782),
.B(n_909),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_782),
.B(n_784),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_864),
.A2(n_696),
.B(n_694),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_790),
.B(n_767),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_783),
.B(n_311),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_876),
.A2(n_767),
.B(n_694),
.C(n_696),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_927),
.A2(n_696),
.B(n_694),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_938),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_858),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_797),
.B(n_734),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_812),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_810),
.B(n_734),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_897),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_882),
.A2(n_538),
.B(n_532),
.C(n_533),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_939),
.Y(n_1069)
);

NOR2x1_ASAP7_75t_L g1070 ( 
.A(n_788),
.B(n_898),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_774),
.A2(n_696),
.B1(n_707),
.B2(n_325),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_877),
.A2(n_729),
.B(n_726),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_778),
.A2(n_788),
.B(n_829),
.C(n_834),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_812),
.Y(n_1074)
);

NOR2xp67_ASAP7_75t_L g1075 ( 
.A(n_841),
.B(n_707),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_836),
.B(n_734),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_837),
.A2(n_707),
.B(n_748),
.C(n_710),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_778),
.A2(n_534),
.B(n_535),
.C(n_559),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_927),
.A2(n_707),
.B(n_671),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_843),
.B(n_734),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_848),
.B(n_741),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_899),
.B(n_789),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_928),
.A2(n_695),
.B(n_669),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_866),
.A2(n_699),
.B(n_695),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_886),
.B(n_296),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_848),
.B(n_741),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_819),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_820),
.A2(n_534),
.B(n_535),
.C(n_538),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_916),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_926),
.B(n_313),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_830),
.A2(n_547),
.B(n_549),
.C(n_543),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_884),
.B(n_288),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_877),
.A2(n_410),
.B1(n_328),
.B2(n_336),
.Y(n_1093)
);

INVxp67_ASAP7_75t_L g1094 ( 
.A(n_930),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_849),
.A2(n_385),
.B1(n_321),
.B2(n_416),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_867),
.A2(n_710),
.B(n_699),
.Y(n_1096)
);

INVxp67_ASAP7_75t_L g1097 ( 
.A(n_849),
.Y(n_1097)
);

NOR2xp67_ASAP7_75t_L g1098 ( 
.A(n_871),
.B(n_351),
.Y(n_1098)
);

OR2x6_ASAP7_75t_L g1099 ( 
.A(n_865),
.B(n_288),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_808),
.A2(n_748),
.B(n_715),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_918),
.A2(n_940),
.B(n_932),
.C(n_931),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_865),
.Y(n_1102)
);

INVx4_ASAP7_75t_L g1103 ( 
.A(n_865),
.Y(n_1103)
);

NOR2xp67_ASAP7_75t_L g1104 ( 
.A(n_883),
.B(n_352),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_859),
.B(n_297),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_915),
.A2(n_549),
.B(n_545),
.C(n_547),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_922),
.B(n_299),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_865),
.B(n_354),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_880),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_814),
.A2(n_729),
.B(n_726),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_880),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_880),
.B(n_741),
.Y(n_1112)
);

NAND2xp33_ASAP7_75t_L g1113 ( 
.A(n_880),
.B(n_358),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_891),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_904),
.A2(n_405),
.B1(n_361),
.B2(n_370),
.Y(n_1115)
);

BUFx8_ASAP7_75t_L g1116 ( 
.A(n_891),
.Y(n_1116)
);

INVxp67_ASAP7_75t_SL g1117 ( 
.A(n_904),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_905),
.A2(n_411),
.B1(n_402),
.B2(n_360),
.Y(n_1118)
);

OAI321xp33_ASAP7_75t_L g1119 ( 
.A1(n_868),
.A2(n_298),
.A3(n_379),
.B1(n_380),
.B2(n_384),
.C(n_369),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_883),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_888),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_888),
.B(n_741),
.Y(n_1122)
);

NAND2x1p5_ASAP7_75t_L g1123 ( 
.A(n_905),
.B(n_715),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_921),
.B(n_300),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_917),
.A2(n_377),
.B1(n_394),
.B2(n_391),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_894),
.B(n_289),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_894),
.B(n_750),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_895),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_815),
.A2(n_750),
.B(n_739),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_SL g1130 ( 
.A1(n_961),
.A2(n_320),
.B1(n_305),
.B2(n_307),
.Y(n_1130)
);

AOI222xp33_ASAP7_75t_L g1131 ( 
.A1(n_1085),
.A2(n_324),
.B1(n_298),
.B2(n_304),
.C1(n_323),
.C2(n_330),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1011),
.B(n_895),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1004),
.B(n_319),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_R g1134 ( 
.A(n_1067),
.B(n_920),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1016),
.A2(n_923),
.B1(n_816),
.B2(n_831),
.Y(n_1135)
);

BUFx8_ASAP7_75t_L g1136 ( 
.A(n_969),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_992),
.A2(n_833),
.B(n_817),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_1022),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_945),
.B(n_902),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_958),
.B(n_902),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_994),
.B(n_903),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1028),
.A2(n_824),
.B(n_906),
.C(n_912),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_952),
.A2(n_908),
.B(n_919),
.C(n_912),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_1015),
.B(n_903),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_982),
.B(n_1003),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_957),
.A2(n_907),
.B1(n_919),
.B2(n_908),
.Y(n_1146)
);

OA21x2_ASAP7_75t_L g1147 ( 
.A1(n_944),
.A2(n_907),
.B(n_911),
.Y(n_1147)
);

AOI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_1045),
.A2(n_327),
.B(n_329),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_991),
.B(n_1053),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_947),
.A2(n_924),
.B1(n_911),
.B2(n_892),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_942),
.A2(n_924),
.B(n_892),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_949),
.A2(n_875),
.B(n_739),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1128),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_963),
.A2(n_875),
.B(n_342),
.C(n_343),
.Y(n_1154)
);

INVxp67_ASAP7_75t_SL g1155 ( 
.A(n_1022),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_967),
.A2(n_397),
.B1(n_388),
.B2(n_382),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1116),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1117),
.A2(n_356),
.B1(n_393),
.B2(n_343),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_948),
.A2(n_739),
.B(n_736),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1117),
.A2(n_736),
.B1(n_375),
.B2(n_386),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_941),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_997),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1024),
.B(n_217),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_943),
.A2(n_736),
.B1(n_373),
.B2(n_390),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_973),
.B(n_667),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1092),
.B(n_331),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_997),
.B(n_332),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1024),
.B(n_1075),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_984),
.B(n_1047),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_1009),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_951),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1047),
.B(n_217),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_960),
.A2(n_346),
.B1(n_368),
.B2(n_369),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_L g1174 ( 
.A(n_1105),
.B(n_399),
.C(n_335),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1009),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1022),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1070),
.A2(n_1094),
.B1(n_1059),
.B2(n_1107),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_978),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_985),
.A2(n_401),
.B1(n_340),
.B2(n_344),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1034),
.B(n_272),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_1099),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_968),
.A2(n_667),
.B(n_793),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_993),
.A2(n_1044),
.B(n_1002),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_1116),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1094),
.B(n_338),
.Y(n_1185)
);

O2A1O1Ixp5_ASAP7_75t_L g1186 ( 
.A1(n_1023),
.A2(n_559),
.B(n_552),
.C(n_551),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1097),
.B(n_1114),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_981),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_946),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1022),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1008),
.B(n_545),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1120),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1019),
.B(n_551),
.Y(n_1193)
);

CKINVDCx8_ASAP7_75t_R g1194 ( 
.A(n_1025),
.Y(n_1194)
);

INVxp33_ASAP7_75t_SL g1195 ( 
.A(n_1082),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1031),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_981),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1092),
.B(n_339),
.Y(n_1198)
);

CKINVDCx14_ASAP7_75t_R g1199 ( 
.A(n_1063),
.Y(n_1199)
);

BUFx4f_ASAP7_75t_L g1200 ( 
.A(n_981),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1089),
.B(n_362),
.Y(n_1201)
);

OAI22x1_ASAP7_75t_L g1202 ( 
.A1(n_1089),
.A2(n_404),
.B1(n_365),
.B2(n_367),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1031),
.B(n_272),
.Y(n_1203)
);

CKINVDCx8_ASAP7_75t_R g1204 ( 
.A(n_1031),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_964),
.A2(n_406),
.B(n_346),
.C(n_368),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1046),
.B(n_552),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1062),
.B(n_371),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1069),
.B(n_372),
.Y(n_1208)
);

O2A1O1Ixp5_ASAP7_75t_L g1209 ( 
.A1(n_962),
.A2(n_548),
.B(n_345),
.C(n_272),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_974),
.B(n_392),
.Y(n_1210)
);

O2A1O1Ixp5_ASAP7_75t_L g1211 ( 
.A1(n_986),
.A2(n_548),
.B(n_345),
.C(n_272),
.Y(n_1211)
);

O2A1O1Ixp5_ASAP7_75t_L g1212 ( 
.A1(n_1012),
.A2(n_548),
.B(n_345),
.C(n_96),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1001),
.A2(n_93),
.B(n_207),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_995),
.A2(n_174),
.B(n_102),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1031),
.B(n_345),
.Y(n_1215)
);

AO21x1_ASAP7_75t_L g1216 ( 
.A1(n_1073),
.A2(n_1020),
.B(n_1018),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1042),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_996),
.A2(n_176),
.B(n_106),
.Y(n_1218)
);

OAI22x1_ASAP7_75t_L g1219 ( 
.A1(n_1124),
.A2(n_417),
.B1(n_415),
.B2(n_413),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1073),
.A2(n_409),
.B(n_408),
.C(n_17),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1000),
.A2(n_196),
.B(n_194),
.Y(n_1221)
);

INVxp67_ASAP7_75t_L g1222 ( 
.A(n_1099),
.Y(n_1222)
);

INVx4_ASAP7_75t_L g1223 ( 
.A(n_1041),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1099),
.Y(n_1224)
);

NOR3xp33_ASAP7_75t_SL g1225 ( 
.A(n_1119),
.B(n_13),
.C(n_15),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1055),
.B(n_13),
.Y(n_1226)
);

INVxp67_ASAP7_75t_L g1227 ( 
.A(n_1126),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_950),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_953),
.B(n_17),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_999),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1041),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1007),
.Y(n_1232)
);

AOI21x1_ASAP7_75t_L g1233 ( 
.A1(n_998),
.A2(n_193),
.B(n_192),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1041),
.B(n_190),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1126),
.B(n_19),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1101),
.A2(n_183),
.B(n_182),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1097),
.B(n_1114),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1087),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1121),
.B(n_1056),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1041),
.B(n_180),
.Y(n_1240)
);

INVx4_ASAP7_75t_L g1241 ( 
.A(n_1102),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1101),
.A2(n_975),
.B(n_972),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_977),
.A2(n_1020),
.B(n_990),
.C(n_1029),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1102),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1102),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1065),
.B(n_21),
.Y(n_1246)
);

OAI21xp33_ASAP7_75t_L g1247 ( 
.A1(n_1095),
.A2(n_21),
.B(n_22),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_1021),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1074),
.B(n_22),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1090),
.B(n_24),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_959),
.A2(n_177),
.B(n_173),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1104),
.A2(n_163),
.B1(n_155),
.B2(n_153),
.Y(n_1252)
);

INVxp33_ASAP7_75t_SL g1253 ( 
.A(n_1118),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1078),
.A2(n_1039),
.B(n_1040),
.C(n_1072),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1102),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1109),
.B(n_24),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1111),
.Y(n_1257)
);

INVxp67_ASAP7_75t_L g1258 ( 
.A(n_1111),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1093),
.A2(n_25),
.B(n_28),
.C(n_30),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1111),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1122),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1048),
.A2(n_146),
.B1(n_145),
.B2(n_134),
.Y(n_1262)
);

BUFx8_ASAP7_75t_SL g1263 ( 
.A(n_1111),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1109),
.B(n_30),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1030),
.B(n_31),
.Y(n_1265)
);

CKINVDCx16_ASAP7_75t_R g1266 ( 
.A(n_954),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1078),
.A2(n_33),
.B(n_34),
.C(n_39),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1035),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_SL g1269 ( 
.A(n_1103),
.B(n_120),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1103),
.B(n_118),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1043),
.B(n_112),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1125),
.B(n_33),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1049),
.B(n_40),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1115),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1052),
.B(n_44),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1127),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1098),
.B(n_46),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_R g1278 ( 
.A(n_1113),
.B(n_115),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1079),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1037),
.B(n_47),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1058),
.B(n_1081),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1123),
.B(n_1086),
.Y(n_1282)
);

O2A1O1Ixp5_ASAP7_75t_SL g1283 ( 
.A1(n_1071),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1123),
.B(n_56),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1038),
.B(n_58),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1013),
.B(n_59),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_956),
.A2(n_76),
.B(n_63),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_971),
.A2(n_60),
.B(n_63),
.Y(n_1288)
);

INVx6_ASAP7_75t_L g1289 ( 
.A(n_1108),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1112),
.A2(n_64),
.B(n_65),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1183),
.A2(n_1242),
.B(n_1137),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1159),
.A2(n_1017),
.B(n_980),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1149),
.B(n_1064),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1138),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1210),
.B(n_1066),
.Y(n_1295)
);

BUFx2_ASAP7_75t_R g1296 ( 
.A(n_1194),
.Y(n_1296)
);

AO21x2_ASAP7_75t_L g1297 ( 
.A1(n_1216),
.A2(n_987),
.B(n_989),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1170),
.Y(n_1298)
);

INVx1_ASAP7_75t_SL g1299 ( 
.A(n_1175),
.Y(n_1299)
);

AO31x2_ASAP7_75t_L g1300 ( 
.A1(n_1254),
.A2(n_1077),
.A3(n_1026),
.B(n_1060),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1144),
.B(n_1145),
.Y(n_1301)
);

CKINVDCx11_ASAP7_75t_R g1302 ( 
.A(n_1184),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1238),
.Y(n_1303)
);

AO31x2_ASAP7_75t_L g1304 ( 
.A1(n_1243),
.A2(n_979),
.A3(n_976),
.B(n_1129),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1135),
.A2(n_1100),
.B(n_1096),
.Y(n_1305)
);

CKINVDCx11_ASAP7_75t_R g1306 ( 
.A(n_1157),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1148),
.A2(n_1220),
.B(n_1272),
.C(n_1259),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1263),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1253),
.B(n_983),
.Y(n_1309)
);

A2O1A1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1177),
.A2(n_988),
.B(n_1068),
.C(n_1014),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1138),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1139),
.A2(n_955),
.B(n_965),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1192),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1143),
.A2(n_1084),
.B(n_1054),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1132),
.A2(n_1033),
.B(n_970),
.Y(n_1315)
);

INVx2_ASAP7_75t_SL g1316 ( 
.A(n_1175),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1162),
.Y(n_1317)
);

AOI221x1_ASAP7_75t_L g1318 ( 
.A1(n_1267),
.A2(n_1032),
.B1(n_1027),
.B2(n_1110),
.C(n_1057),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1161),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1142),
.A2(n_1212),
.B(n_1151),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1144),
.B(n_1080),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1154),
.A2(n_1005),
.A3(n_1010),
.B(n_1083),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1281),
.A2(n_1013),
.B(n_1051),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1165),
.A2(n_1061),
.B(n_966),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1187),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1212),
.A2(n_1050),
.B(n_1068),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1134),
.B(n_1006),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1227),
.A2(n_1036),
.B1(n_1076),
.B2(n_1088),
.Y(n_1328)
);

OR2x6_ASAP7_75t_L g1329 ( 
.A(n_1188),
.B(n_1197),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1155),
.A2(n_1091),
.B(n_1088),
.Y(n_1330)
);

AO31x2_ASAP7_75t_L g1331 ( 
.A1(n_1236),
.A2(n_1106),
.A3(n_1014),
.B(n_988),
.Y(n_1331)
);

CKINVDCx11_ASAP7_75t_R g1332 ( 
.A(n_1187),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1152),
.A2(n_1091),
.B(n_1106),
.Y(n_1333)
);

AOI221x1_ASAP7_75t_L g1334 ( 
.A1(n_1247),
.A2(n_1288),
.B1(n_1279),
.B2(n_1287),
.C(n_1286),
.Y(n_1334)
);

NAND3xp33_ASAP7_75t_L g1335 ( 
.A(n_1185),
.B(n_67),
.C(n_69),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1195),
.B(n_70),
.Y(n_1336)
);

AND2x2_ASAP7_75t_SL g1337 ( 
.A(n_1269),
.B(n_70),
.Y(n_1337)
);

BUFx4f_ASAP7_75t_SL g1338 ( 
.A(n_1136),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1150),
.A2(n_73),
.B(n_1182),
.Y(n_1339)
);

AOI221x1_ASAP7_75t_L g1340 ( 
.A1(n_1290),
.A2(n_1213),
.B1(n_1250),
.B2(n_1265),
.C(n_1280),
.Y(n_1340)
);

AOI221x1_ASAP7_75t_L g1341 ( 
.A1(n_1250),
.A2(n_1280),
.B1(n_1265),
.B2(n_1226),
.C(n_1202),
.Y(n_1341)
);

AOI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1282),
.A2(n_1140),
.B(n_1146),
.Y(n_1342)
);

AO32x2_ASAP7_75t_L g1343 ( 
.A1(n_1164),
.A2(n_1160),
.A3(n_1179),
.B1(n_1130),
.B2(n_1283),
.Y(n_1343)
);

NAND3x1_ASAP7_75t_L g1344 ( 
.A(n_1167),
.B(n_1201),
.C(n_1166),
.Y(n_1344)
);

CKINVDCx8_ASAP7_75t_R g1345 ( 
.A(n_1237),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1224),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1181),
.Y(n_1347)
);

NOR4xp25_ASAP7_75t_L g1348 ( 
.A(n_1274),
.B(n_1173),
.C(n_1205),
.D(n_1158),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1237),
.Y(n_1349)
);

INVxp67_ASAP7_75t_L g1350 ( 
.A(n_1167),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1248),
.B(n_1222),
.Y(n_1351)
);

BUFx5_ASAP7_75t_L g1352 ( 
.A(n_1271),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1227),
.B(n_1222),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1189),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1133),
.B(n_1208),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1141),
.A2(n_1168),
.B(n_1268),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1266),
.B(n_1248),
.Y(n_1357)
);

AO31x2_ASAP7_75t_L g1358 ( 
.A1(n_1226),
.A2(n_1285),
.A3(n_1229),
.B(n_1251),
.Y(n_1358)
);

AOI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1173),
.A2(n_1207),
.B1(n_1235),
.B2(n_1225),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1186),
.A2(n_1221),
.B(n_1233),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1228),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1276),
.B(n_1207),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1174),
.B(n_1200),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1204),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1158),
.B(n_1239),
.Y(n_1365)
);

AOI21xp33_ASAP7_75t_L g1366 ( 
.A1(n_1156),
.A2(n_1198),
.B(n_1180),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1155),
.A2(n_1261),
.B(n_1147),
.Y(n_1367)
);

AO32x2_ASAP7_75t_L g1368 ( 
.A1(n_1223),
.A2(n_1241),
.A3(n_1209),
.B1(n_1211),
.B2(n_1225),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1230),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1181),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1209),
.A2(n_1186),
.B(n_1211),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1200),
.B(n_1219),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1289),
.B(n_1172),
.Y(n_1373)
);

AO21x2_ASAP7_75t_L g1374 ( 
.A1(n_1273),
.A2(n_1275),
.B(n_1256),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1232),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1191),
.B(n_1193),
.Y(n_1376)
);

O2A1O1Ixp33_ASAP7_75t_L g1377 ( 
.A1(n_1163),
.A2(n_1277),
.B(n_1215),
.C(n_1203),
.Y(n_1377)
);

CKINVDCx11_ASAP7_75t_R g1378 ( 
.A(n_1199),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1271),
.A2(n_1262),
.B(n_1252),
.C(n_1169),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1264),
.A2(n_1246),
.A3(n_1249),
.B(n_1214),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1217),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1289),
.A2(n_1178),
.B1(n_1171),
.B2(n_1258),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_1289),
.Y(n_1383)
);

AO21x1_ASAP7_75t_L g1384 ( 
.A1(n_1284),
.A2(n_1240),
.B(n_1234),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1218),
.A2(n_1206),
.B(n_1270),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1258),
.A2(n_1231),
.B(n_1244),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1244),
.A2(n_1257),
.B(n_1131),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1138),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1257),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1255),
.A2(n_1260),
.B(n_1245),
.C(n_1190),
.Y(n_1390)
);

NAND3xp33_ASAP7_75t_SL g1391 ( 
.A(n_1278),
.B(n_1223),
.C(n_1241),
.Y(n_1391)
);

AO31x2_ASAP7_75t_L g1392 ( 
.A1(n_1138),
.A2(n_1176),
.A3(n_1190),
.B(n_1196),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1176),
.A2(n_1190),
.B(n_1196),
.Y(n_1393)
);

AO31x2_ASAP7_75t_L g1394 ( 
.A1(n_1176),
.A2(n_1216),
.A3(n_1254),
.B(n_1242),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1176),
.A2(n_1190),
.B(n_1196),
.Y(n_1395)
);

CKINVDCx8_ASAP7_75t_R g1396 ( 
.A(n_1196),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1177),
.A2(n_961),
.B(n_825),
.C(n_945),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1153),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1183),
.A2(n_992),
.B(n_963),
.Y(n_1399)
);

OA21x2_ASAP7_75t_L g1400 ( 
.A1(n_1212),
.A2(n_1254),
.B(n_1216),
.Y(n_1400)
);

CKINVDCx11_ASAP7_75t_R g1401 ( 
.A(n_1194),
.Y(n_1401)
);

INVx6_ASAP7_75t_SL g1402 ( 
.A(n_1187),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1149),
.B(n_961),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1183),
.A2(n_992),
.B(n_963),
.Y(n_1404)
);

AO31x2_ASAP7_75t_L g1405 ( 
.A1(n_1216),
.A2(n_1254),
.A3(n_1242),
.B(n_1243),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1153),
.Y(n_1406)
);

AO31x2_ASAP7_75t_L g1407 ( 
.A1(n_1216),
.A2(n_1254),
.A3(n_1242),
.B(n_1243),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1177),
.A2(n_961),
.B(n_825),
.C(n_945),
.Y(n_1408)
);

AO21x2_ASAP7_75t_L g1409 ( 
.A1(n_1242),
.A2(n_1183),
.B(n_1216),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1253),
.A2(n_1028),
.B1(n_1272),
.B2(n_1149),
.Y(n_1410)
);

NAND3xp33_ASAP7_75t_L g1411 ( 
.A(n_1272),
.B(n_825),
.C(n_961),
.Y(n_1411)
);

AOI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1242),
.A2(n_1159),
.B(n_1183),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1149),
.B(n_423),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1177),
.A2(n_961),
.B(n_825),
.C(n_945),
.Y(n_1414)
);

AO31x2_ASAP7_75t_L g1415 ( 
.A1(n_1216),
.A2(n_1254),
.A3(n_1242),
.B(n_1243),
.Y(n_1415)
);

INVx3_ASAP7_75t_SL g1416 ( 
.A(n_1187),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1153),
.Y(n_1417)
);

AO31x2_ASAP7_75t_L g1418 ( 
.A1(n_1216),
.A2(n_1254),
.A3(n_1242),
.B(n_1243),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1170),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1170),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_SL g1421 ( 
.A1(n_1220),
.A2(n_961),
.B(n_1016),
.C(n_952),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1149),
.B(n_961),
.Y(n_1422)
);

OA21x2_ASAP7_75t_L g1423 ( 
.A1(n_1212),
.A2(n_1254),
.B(n_1216),
.Y(n_1423)
);

AOI31xp67_ASAP7_75t_L g1424 ( 
.A1(n_1286),
.A2(n_778),
.A3(n_655),
.B(n_631),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1183),
.A2(n_992),
.B(n_963),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1153),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1149),
.B(n_1015),
.Y(n_1427)
);

AO31x2_ASAP7_75t_L g1428 ( 
.A1(n_1216),
.A2(n_1254),
.A3(n_1242),
.B(n_1243),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_SL g1429 ( 
.A(n_1269),
.B(n_961),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1212),
.A2(n_1254),
.B(n_1216),
.Y(n_1430)
);

AOI221x1_ASAP7_75t_L g1431 ( 
.A1(n_1220),
.A2(n_961),
.B1(n_1267),
.B2(n_1236),
.C(n_1242),
.Y(n_1431)
);

AO32x2_ASAP7_75t_L g1432 ( 
.A1(n_1135),
.A2(n_1164),
.A3(n_1150),
.B1(n_1160),
.B2(n_1146),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1149),
.B(n_770),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1149),
.B(n_1015),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1183),
.A2(n_992),
.B(n_963),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1183),
.A2(n_1023),
.B(n_1242),
.Y(n_1436)
);

AOI221xp5_ASAP7_75t_SL g1437 ( 
.A1(n_1173),
.A2(n_961),
.B1(n_1247),
.B2(n_1158),
.C(n_1259),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1183),
.A2(n_992),
.B(n_963),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1149),
.B(n_961),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1183),
.A2(n_992),
.B(n_963),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1153),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1149),
.B(n_1015),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1183),
.A2(n_1023),
.B(n_1242),
.Y(n_1443)
);

BUFx3_ASAP7_75t_L g1444 ( 
.A(n_1170),
.Y(n_1444)
);

CKINVDCx14_ASAP7_75t_R g1445 ( 
.A(n_1199),
.Y(n_1445)
);

OAI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1254),
.A2(n_1016),
.B(n_942),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1149),
.B(n_770),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_SL g1448 ( 
.A(n_1157),
.Y(n_1448)
);

O2A1O1Ixp33_ASAP7_75t_SL g1449 ( 
.A1(n_1220),
.A2(n_961),
.B(n_1016),
.C(n_952),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1254),
.A2(n_1016),
.B(n_942),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1183),
.A2(n_992),
.B(n_963),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1183),
.A2(n_992),
.B(n_963),
.Y(n_1452)
);

A2O1A1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1177),
.A2(n_961),
.B(n_825),
.C(n_945),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1401),
.Y(n_1454)
);

OAI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1359),
.A2(n_1429),
.B1(n_1335),
.B2(n_1411),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1313),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1410),
.A2(n_1350),
.B1(n_1359),
.B2(n_1309),
.Y(n_1457)
);

INVx6_ASAP7_75t_L g1458 ( 
.A(n_1364),
.Y(n_1458)
);

BUFx12f_ASAP7_75t_L g1459 ( 
.A(n_1378),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1403),
.B(n_1422),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1349),
.Y(n_1461)
);

INVx8_ASAP7_75t_L g1462 ( 
.A(n_1364),
.Y(n_1462)
);

INVx6_ASAP7_75t_L g1463 ( 
.A(n_1364),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1319),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1354),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1411),
.A2(n_1335),
.B1(n_1337),
.B2(n_1439),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1361),
.Y(n_1467)
);

INVx2_ASAP7_75t_SL g1468 ( 
.A(n_1420),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1362),
.A2(n_1427),
.B1(n_1442),
.B2(n_1434),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1444),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1341),
.A2(n_1307),
.B(n_1366),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1302),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_SL g1473 ( 
.A1(n_1429),
.A2(n_1336),
.B1(n_1450),
.B2(n_1446),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1298),
.Y(n_1474)
);

OAI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1301),
.A2(n_1376),
.B1(n_1355),
.B2(n_1293),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_1338),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1369),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1353),
.B(n_1325),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1446),
.A2(n_1450),
.B1(n_1447),
.B2(n_1433),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1419),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1413),
.A2(n_1365),
.B1(n_1373),
.B2(n_1295),
.Y(n_1481)
);

BUFx4f_ASAP7_75t_L g1482 ( 
.A(n_1308),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1397),
.B(n_1408),
.Y(n_1483)
);

BUFx8_ASAP7_75t_L g1484 ( 
.A(n_1448),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1414),
.A2(n_1453),
.B1(n_1351),
.B2(n_1344),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1372),
.A2(n_1363),
.B1(n_1384),
.B2(n_1353),
.Y(n_1486)
);

BUFx8_ASAP7_75t_L g1487 ( 
.A(n_1448),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1375),
.Y(n_1488)
);

OAI21xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1320),
.A2(n_1348),
.B(n_1327),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1383),
.A2(n_1437),
.B1(n_1357),
.B2(n_1329),
.Y(n_1490)
);

CKINVDCx11_ASAP7_75t_R g1491 ( 
.A(n_1306),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1387),
.A2(n_1352),
.B1(n_1347),
.B2(n_1329),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_SL g1493 ( 
.A1(n_1379),
.A2(n_1340),
.B(n_1377),
.Y(n_1493)
);

INVx4_ASAP7_75t_L g1494 ( 
.A(n_1308),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1387),
.A2(n_1320),
.B1(n_1339),
.B2(n_1423),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1400),
.A2(n_1423),
.B1(n_1430),
.B2(n_1297),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1400),
.A2(n_1430),
.B1(n_1297),
.B2(n_1406),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1299),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1381),
.Y(n_1499)
);

CKINVDCx20_ASAP7_75t_R g1500 ( 
.A(n_1445),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1402),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1394),
.Y(n_1502)
);

OAI21xp33_ASAP7_75t_L g1503 ( 
.A1(n_1348),
.A2(n_1321),
.B(n_1310),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1370),
.A2(n_1345),
.B1(n_1390),
.B2(n_1316),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1398),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1417),
.A2(n_1441),
.B1(n_1426),
.B2(n_1437),
.Y(n_1506)
);

INVx11_ASAP7_75t_L g1507 ( 
.A(n_1402),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1374),
.A2(n_1333),
.B1(n_1356),
.B2(n_1326),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1374),
.A2(n_1333),
.B1(n_1326),
.B2(n_1352),
.Y(n_1509)
);

BUFx4_ASAP7_75t_R g1510 ( 
.A(n_1296),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1352),
.A2(n_1409),
.B1(n_1389),
.B2(n_1371),
.Y(n_1511)
);

CKINVDCx11_ASAP7_75t_R g1512 ( 
.A(n_1416),
.Y(n_1512)
);

INVx1_ASAP7_75t_SL g1513 ( 
.A(n_1317),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1346),
.A2(n_1382),
.B1(n_1396),
.B2(n_1330),
.Y(n_1514)
);

BUFx8_ASAP7_75t_L g1515 ( 
.A(n_1388),
.Y(n_1515)
);

BUFx5_ASAP7_75t_L g1516 ( 
.A(n_1412),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1352),
.A2(n_1409),
.B1(n_1371),
.B2(n_1332),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1352),
.A2(n_1328),
.B1(n_1305),
.B2(n_1391),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1392),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_SL g1520 ( 
.A1(n_1388),
.A2(n_1294),
.B1(n_1311),
.B2(n_1343),
.Y(n_1520)
);

INVx6_ASAP7_75t_L g1521 ( 
.A(n_1294),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1311),
.B(n_1343),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1386),
.A2(n_1385),
.B1(n_1312),
.B2(n_1305),
.Y(n_1523)
);

NAND2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1393),
.B(n_1395),
.Y(n_1524)
);

CKINVDCx11_ASAP7_75t_R g1525 ( 
.A(n_1421),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1392),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1314),
.A2(n_1449),
.B1(n_1324),
.B2(n_1367),
.Y(n_1527)
);

CKINVDCx6p67_ASAP7_75t_R g1528 ( 
.A(n_1343),
.Y(n_1528)
);

BUFx4f_ASAP7_75t_SL g1529 ( 
.A(n_1334),
.Y(n_1529)
);

BUFx8_ASAP7_75t_L g1530 ( 
.A(n_1368),
.Y(n_1530)
);

BUFx2_ASAP7_75t_R g1531 ( 
.A(n_1368),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1358),
.B(n_1428),
.Y(n_1532)
);

BUFx10_ASAP7_75t_L g1533 ( 
.A(n_1358),
.Y(n_1533)
);

BUFx12f_ASAP7_75t_L g1534 ( 
.A(n_1424),
.Y(n_1534)
);

BUFx10_ASAP7_75t_L g1535 ( 
.A(n_1431),
.Y(n_1535)
);

BUFx10_ASAP7_75t_L g1536 ( 
.A(n_1368),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1394),
.Y(n_1537)
);

INVx4_ASAP7_75t_L g1538 ( 
.A(n_1342),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1405),
.Y(n_1539)
);

BUFx12f_ASAP7_75t_L g1540 ( 
.A(n_1380),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1314),
.A2(n_1323),
.B1(n_1315),
.B2(n_1399),
.Y(n_1541)
);

INVx4_ASAP7_75t_L g1542 ( 
.A(n_1380),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_SL g1543 ( 
.A1(n_1432),
.A2(n_1415),
.B1(n_1428),
.B2(n_1418),
.Y(n_1543)
);

BUFx2_ASAP7_75t_SL g1544 ( 
.A(n_1404),
.Y(n_1544)
);

INVx1_ASAP7_75t_SL g1545 ( 
.A(n_1425),
.Y(n_1545)
);

NAND2x1p5_ASAP7_75t_L g1546 ( 
.A(n_1436),
.B(n_1443),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1435),
.A2(n_1452),
.B1(n_1451),
.B2(n_1440),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1438),
.A2(n_1291),
.B1(n_1432),
.B2(n_1292),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1407),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_SL g1550 ( 
.A1(n_1432),
.A2(n_1428),
.B1(n_1418),
.B2(n_1415),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1407),
.A2(n_1418),
.B1(n_1415),
.B2(n_1300),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1318),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1360),
.A2(n_1300),
.B1(n_1331),
.B2(n_1304),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1300),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1304),
.A2(n_1410),
.B1(n_1411),
.B2(n_1272),
.Y(n_1555)
);

NAND2x1p5_ASAP7_75t_L g1556 ( 
.A(n_1322),
.B(n_1304),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1331),
.A2(n_1411),
.B1(n_961),
.B2(n_1410),
.Y(n_1557)
);

OAI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1331),
.A2(n_961),
.B1(n_1359),
.B2(n_1429),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1322),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1313),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1364),
.Y(n_1561)
);

INVx2_ASAP7_75t_SL g1562 ( 
.A(n_1349),
.Y(n_1562)
);

INVx2_ASAP7_75t_SL g1563 ( 
.A(n_1349),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1411),
.A2(n_961),
.B1(n_1410),
.B2(n_1335),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1298),
.Y(n_1565)
);

INVx6_ASAP7_75t_L g1566 ( 
.A(n_1364),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1303),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1411),
.A2(n_961),
.B1(n_1410),
.B2(n_1335),
.Y(n_1568)
);

BUFx12f_ASAP7_75t_L g1569 ( 
.A(n_1378),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1303),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1420),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_SL g1572 ( 
.A1(n_1337),
.A2(n_1429),
.B1(n_961),
.B2(n_1335),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1303),
.Y(n_1573)
);

BUFx10_ASAP7_75t_L g1574 ( 
.A(n_1308),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1401),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1303),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1411),
.A2(n_961),
.B1(n_1410),
.B2(n_1335),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1410),
.A2(n_961),
.B1(n_825),
.B2(n_1350),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1411),
.A2(n_961),
.B1(n_1410),
.B2(n_1335),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1364),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1364),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1396),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1401),
.Y(n_1583)
);

CKINVDCx20_ASAP7_75t_R g1584 ( 
.A(n_1401),
.Y(n_1584)
);

INVx6_ASAP7_75t_L g1585 ( 
.A(n_1364),
.Y(n_1585)
);

CKINVDCx20_ASAP7_75t_R g1586 ( 
.A(n_1401),
.Y(n_1586)
);

INVx4_ASAP7_75t_L g1587 ( 
.A(n_1364),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1337),
.A2(n_1429),
.B1(n_961),
.B2(n_1335),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1411),
.A2(n_961),
.B1(n_1410),
.B2(n_1335),
.Y(n_1589)
);

AOI21xp33_ASAP7_75t_L g1590 ( 
.A1(n_1307),
.A2(n_1028),
.B(n_825),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1364),
.Y(n_1591)
);

INVx6_ASAP7_75t_L g1592 ( 
.A(n_1364),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1411),
.A2(n_961),
.B1(n_1410),
.B2(n_1335),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1337),
.A2(n_1429),
.B1(n_961),
.B2(n_1335),
.Y(n_1594)
);

BUFx4f_ASAP7_75t_L g1595 ( 
.A(n_1364),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1313),
.Y(n_1596)
);

BUFx8_ASAP7_75t_L g1597 ( 
.A(n_1448),
.Y(n_1597)
);

BUFx10_ASAP7_75t_L g1598 ( 
.A(n_1308),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_SL g1599 ( 
.A1(n_1410),
.A2(n_825),
.B(n_960),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1298),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1410),
.A2(n_1411),
.B1(n_1272),
.B2(n_1028),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1411),
.A2(n_961),
.B1(n_1410),
.B2(n_1335),
.Y(n_1602)
);

CKINVDCx6p67_ASAP7_75t_R g1603 ( 
.A(n_1401),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1411),
.A2(n_961),
.B1(n_1410),
.B2(n_1335),
.Y(n_1604)
);

INVx6_ASAP7_75t_L g1605 ( 
.A(n_1364),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1475),
.B(n_1601),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1457),
.B(n_1460),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1519),
.Y(n_1608)
);

OAI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1590),
.A2(n_1471),
.B(n_1599),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1477),
.Y(n_1610)
);

OR2x6_ASAP7_75t_L g1611 ( 
.A(n_1544),
.B(n_1540),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1526),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1539),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1522),
.B(n_1532),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1549),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1479),
.B(n_1528),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1488),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1537),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1554),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1502),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1502),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1524),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1479),
.B(n_1531),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1464),
.Y(n_1624)
);

OAI21x1_ASAP7_75t_L g1625 ( 
.A1(n_1546),
.A2(n_1523),
.B(n_1547),
.Y(n_1625)
);

AOI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1485),
.A2(n_1483),
.B(n_1559),
.Y(n_1626)
);

CKINVDCx11_ASAP7_75t_R g1627 ( 
.A(n_1584),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1465),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1498),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1531),
.B(n_1473),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1545),
.A2(n_1547),
.B(n_1541),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1515),
.Y(n_1632)
);

INVxp67_ASAP7_75t_L g1633 ( 
.A(n_1513),
.Y(n_1633)
);

NAND2x1p5_ASAP7_75t_L g1634 ( 
.A(n_1542),
.B(n_1538),
.Y(n_1634)
);

INVx6_ASAP7_75t_L g1635 ( 
.A(n_1515),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1467),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1552),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1567),
.Y(n_1638)
);

INVx6_ASAP7_75t_L g1639 ( 
.A(n_1462),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1570),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1573),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1576),
.Y(n_1642)
);

AO21x2_ASAP7_75t_L g1643 ( 
.A1(n_1455),
.A2(n_1558),
.B(n_1493),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1551),
.Y(n_1644)
);

AOI21xp33_ASAP7_75t_L g1645 ( 
.A1(n_1455),
.A2(n_1589),
.B(n_1568),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1565),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1504),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1533),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1541),
.A2(n_1558),
.B(n_1508),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1533),
.Y(n_1650)
);

AO21x2_ASAP7_75t_L g1651 ( 
.A1(n_1503),
.A2(n_1475),
.B(n_1514),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1530),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1556),
.Y(n_1653)
);

OA21x2_ASAP7_75t_L g1654 ( 
.A1(n_1495),
.A2(n_1496),
.B(n_1548),
.Y(n_1654)
);

NAND2x1p5_ASAP7_75t_L g1655 ( 
.A(n_1542),
.B(n_1538),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1530),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1572),
.A2(n_1594),
.B1(n_1588),
.B2(n_1604),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1546),
.A2(n_1548),
.B(n_1527),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1578),
.A2(n_1572),
.B1(n_1588),
.B2(n_1594),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1527),
.A2(n_1524),
.B(n_1496),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1536),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1534),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1543),
.Y(n_1663)
);

AND2x2_ASAP7_75t_SL g1664 ( 
.A(n_1517),
.B(n_1509),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1543),
.Y(n_1665)
);

AOI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1505),
.A2(n_1499),
.B(n_1456),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1517),
.B(n_1509),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1557),
.B(n_1550),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1469),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1550),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1557),
.B(n_1497),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1489),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1535),
.Y(n_1673)
);

AO21x1_ASAP7_75t_L g1674 ( 
.A1(n_1490),
.A2(n_1529),
.B(n_1604),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1535),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1470),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_1529),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1571),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1497),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1520),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1564),
.A2(n_1593),
.B1(n_1579),
.B2(n_1568),
.Y(n_1681)
);

CKINVDCx14_ASAP7_75t_R g1682 ( 
.A(n_1586),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1555),
.B(n_1508),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1481),
.B(n_1564),
.Y(n_1684)
);

INVx2_ASAP7_75t_SL g1685 ( 
.A(n_1521),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1516),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1481),
.B(n_1511),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1553),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1553),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1511),
.Y(n_1690)
);

INVx4_ASAP7_75t_L g1691 ( 
.A(n_1462),
.Y(n_1691)
);

AO21x2_ASAP7_75t_L g1692 ( 
.A1(n_1495),
.A2(n_1518),
.B(n_1560),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1577),
.A2(n_1579),
.B1(n_1593),
.B2(n_1589),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1600),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1510),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1525),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1474),
.Y(n_1697)
);

OR2x6_ASAP7_75t_L g1698 ( 
.A(n_1462),
.B(n_1587),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1577),
.B(n_1602),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1454),
.Y(n_1700)
);

AO21x2_ASAP7_75t_L g1701 ( 
.A1(n_1518),
.A2(n_1596),
.B(n_1602),
.Y(n_1701)
);

BUFx12f_ASAP7_75t_L g1702 ( 
.A(n_1491),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1506),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1480),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1506),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1492),
.Y(n_1706)
);

OA21x2_ASAP7_75t_L g1707 ( 
.A1(n_1466),
.A2(n_1486),
.B(n_1478),
.Y(n_1707)
);

O2A1O1Ixp33_ASAP7_75t_L g1708 ( 
.A1(n_1466),
.A2(n_1582),
.B(n_1468),
.C(n_1562),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1563),
.A2(n_1461),
.B1(n_1501),
.B2(n_1587),
.C(n_1591),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1561),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1575),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1583),
.B(n_1458),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1582),
.Y(n_1713)
);

OA21x2_ASAP7_75t_L g1714 ( 
.A1(n_1472),
.A2(n_1458),
.B(n_1592),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1561),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1580),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1580),
.B(n_1591),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1580),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1581),
.B(n_1595),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1581),
.Y(n_1720)
);

OA21x2_ASAP7_75t_L g1721 ( 
.A1(n_1458),
.A2(n_1605),
.B(n_1463),
.Y(n_1721)
);

OAI21x1_ASAP7_75t_L g1722 ( 
.A1(n_1605),
.A2(n_1585),
.B(n_1463),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1581),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1566),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1566),
.Y(n_1725)
);

OAI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1609),
.A2(n_1595),
.B(n_1482),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1694),
.Y(n_1727)
);

OAI21x1_ASAP7_75t_SL g1728 ( 
.A1(n_1674),
.A2(n_1626),
.B(n_1659),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1607),
.B(n_1603),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1614),
.B(n_1690),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1690),
.B(n_1494),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1619),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1657),
.A2(n_1482),
.B1(n_1500),
.B2(n_1507),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1669),
.B(n_1597),
.Y(n_1734)
);

NOR2x1_ASAP7_75t_SL g1735 ( 
.A(n_1611),
.B(n_1459),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1613),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1668),
.B(n_1598),
.Y(n_1737)
);

BUFx3_ASAP7_75t_L g1738 ( 
.A(n_1721),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1697),
.B(n_1512),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1663),
.B(n_1574),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1693),
.A2(n_1476),
.B(n_1484),
.Y(n_1741)
);

OR2x6_ASAP7_75t_L g1742 ( 
.A(n_1611),
.B(n_1569),
.Y(n_1742)
);

BUFx3_ASAP7_75t_L g1743 ( 
.A(n_1721),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1699),
.B(n_1484),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1699),
.B(n_1487),
.Y(n_1745)
);

OA21x2_ASAP7_75t_L g1746 ( 
.A1(n_1658),
.A2(n_1597),
.B(n_1574),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1663),
.B(n_1598),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_SL g1748 ( 
.A1(n_1696),
.A2(n_1681),
.B1(n_1695),
.B2(n_1637),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1721),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1646),
.B(n_1695),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1665),
.B(n_1670),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1633),
.B(n_1704),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1613),
.Y(n_1753)
);

CKINVDCx6p67_ASAP7_75t_R g1754 ( 
.A(n_1702),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_1721),
.Y(n_1755)
);

AOI211xp5_ASAP7_75t_L g1756 ( 
.A1(n_1645),
.A2(n_1674),
.B(n_1606),
.C(n_1684),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1629),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1665),
.B(n_1670),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1671),
.B(n_1616),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_1714),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1671),
.B(n_1616),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1637),
.B(n_1700),
.Y(n_1762)
);

OA21x2_ASAP7_75t_L g1763 ( 
.A1(n_1658),
.A2(n_1660),
.B(n_1649),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1688),
.B(n_1689),
.Y(n_1764)
);

AO21x2_ASAP7_75t_L g1765 ( 
.A1(n_1631),
.A2(n_1625),
.B(n_1686),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1679),
.B(n_1644),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1688),
.B(n_1689),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1683),
.B(n_1679),
.Y(n_1768)
);

AOI221xp5_ASAP7_75t_L g1769 ( 
.A1(n_1672),
.A2(n_1630),
.B1(n_1623),
.B2(n_1687),
.C(n_1683),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1651),
.A2(n_1611),
.B(n_1643),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1651),
.A2(n_1611),
.B(n_1643),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1610),
.B(n_1617),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1664),
.B(n_1624),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1628),
.B(n_1636),
.Y(n_1774)
);

AOI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1643),
.A2(n_1651),
.B1(n_1706),
.B2(n_1647),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1628),
.B(n_1636),
.Y(n_1776)
);

OAI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1708),
.A2(n_1687),
.B(n_1626),
.Y(n_1777)
);

A2O1A1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1672),
.A2(n_1623),
.B(n_1677),
.C(n_1667),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1696),
.A2(n_1635),
.B1(n_1677),
.B2(n_1713),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1714),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1610),
.B(n_1617),
.Y(n_1781)
);

OAI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1706),
.A2(n_1713),
.B(n_1678),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1714),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1638),
.B(n_1640),
.Y(n_1784)
);

OA21x2_ASAP7_75t_L g1785 ( 
.A1(n_1644),
.A2(n_1615),
.B(n_1618),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1714),
.Y(n_1786)
);

AO21x2_ASAP7_75t_L g1787 ( 
.A1(n_1648),
.A2(n_1650),
.B(n_1673),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1638),
.B(n_1640),
.Y(n_1788)
);

INVxp67_ASAP7_75t_L g1789 ( 
.A(n_1723),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1707),
.A2(n_1709),
.B1(n_1696),
.B2(n_1701),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1641),
.B(n_1642),
.Y(n_1791)
);

OA21x2_ASAP7_75t_L g1792 ( 
.A1(n_1618),
.A2(n_1608),
.B(n_1612),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1611),
.A2(n_1692),
.B(n_1701),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1700),
.B(n_1711),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_SL g1795 ( 
.A1(n_1682),
.A2(n_1635),
.B1(n_1632),
.B2(n_1702),
.Y(n_1795)
);

AOI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1692),
.A2(n_1701),
.B(n_1677),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1722),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1676),
.A2(n_1675),
.B(n_1673),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1711),
.B(n_1627),
.Y(n_1799)
);

OAI21x1_ASAP7_75t_L g1800 ( 
.A1(n_1634),
.A2(n_1655),
.B(n_1666),
.Y(n_1800)
);

OAI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1635),
.A2(n_1680),
.B1(n_1652),
.B2(n_1656),
.Y(n_1801)
);

AO32x2_ASAP7_75t_L g1802 ( 
.A1(n_1685),
.A2(n_1620),
.A3(n_1621),
.B1(n_1632),
.B2(n_1654),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1730),
.B(n_1661),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1792),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1749),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1759),
.B(n_1761),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1732),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1748),
.A2(n_1667),
.B1(n_1707),
.B2(n_1680),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1802),
.B(n_1654),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1738),
.B(n_1622),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1785),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1768),
.B(n_1764),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1733),
.A2(n_1707),
.B1(n_1652),
.B2(n_1656),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1768),
.B(n_1764),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1760),
.B(n_1620),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1785),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_1738),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1802),
.B(n_1654),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1767),
.B(n_1675),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1802),
.B(n_1654),
.Y(n_1820)
);

OAI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1775),
.A2(n_1707),
.B1(n_1705),
.B2(n_1703),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1736),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1753),
.Y(n_1823)
);

INVx2_ASAP7_75t_SL g1824 ( 
.A(n_1743),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1743),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1760),
.B(n_1621),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1802),
.B(n_1653),
.Y(n_1827)
);

NOR2x1_ASAP7_75t_L g1828 ( 
.A(n_1787),
.B(n_1662),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1755),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1802),
.B(n_1763),
.Y(n_1830)
);

AND2x4_ASAP7_75t_SL g1831 ( 
.A(n_1742),
.B(n_1622),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1774),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1776),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1766),
.B(n_1692),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1729),
.B(n_1712),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1784),
.Y(n_1836)
);

OAI21xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1741),
.A2(n_1719),
.B(n_1705),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1751),
.B(n_1703),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1788),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1817),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1821),
.A2(n_1796),
.B(n_1793),
.Y(n_1841)
);

NAND4xp25_ASAP7_75t_L g1842 ( 
.A(n_1808),
.B(n_1756),
.C(n_1769),
.D(n_1777),
.Y(n_1842)
);

AOI221xp5_ASAP7_75t_L g1843 ( 
.A1(n_1821),
.A2(n_1728),
.B1(n_1778),
.B2(n_1727),
.C(n_1771),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1824),
.B(n_1797),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1827),
.B(n_1780),
.Y(n_1845)
);

OAI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1837),
.A2(n_1790),
.B1(n_1726),
.B2(n_1770),
.C(n_1744),
.Y(n_1846)
);

NAND3xp33_ASAP7_75t_L g1847 ( 
.A(n_1837),
.B(n_1782),
.C(n_1798),
.Y(n_1847)
);

O2A1O1Ixp33_ASAP7_75t_L g1848 ( 
.A1(n_1813),
.A2(n_1728),
.B(n_1745),
.C(n_1734),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1827),
.B(n_1780),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1809),
.B(n_1780),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1822),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1805),
.B(n_1765),
.Y(n_1852)
);

HB1xp67_ASAP7_75t_L g1853 ( 
.A(n_1805),
.Y(n_1853)
);

BUFx2_ASAP7_75t_L g1854 ( 
.A(n_1817),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1804),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1815),
.Y(n_1856)
);

INVx1_ASAP7_75t_SL g1857 ( 
.A(n_1825),
.Y(n_1857)
);

INVx3_ASAP7_75t_L g1858 ( 
.A(n_1810),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1809),
.B(n_1780),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1834),
.B(n_1791),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1815),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1804),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1834),
.B(n_1783),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1822),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1822),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1818),
.B(n_1786),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1826),
.B(n_1765),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1826),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1823),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1816),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1820),
.B(n_1786),
.Y(n_1871)
);

OAI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1812),
.A2(n_1742),
.B1(n_1801),
.B2(n_1779),
.Y(n_1872)
);

INVx3_ASAP7_75t_L g1873 ( 
.A(n_1810),
.Y(n_1873)
);

NAND3xp33_ASAP7_75t_L g1874 ( 
.A(n_1820),
.B(n_1731),
.C(n_1757),
.Y(n_1874)
);

INVx2_ASAP7_75t_SL g1875 ( 
.A(n_1824),
.Y(n_1875)
);

AOI222xp33_ASAP7_75t_L g1876 ( 
.A1(n_1835),
.A2(n_1795),
.B1(n_1762),
.B2(n_1773),
.C1(n_1758),
.C2(n_1751),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1830),
.B(n_1746),
.Y(n_1877)
);

AND2x4_ASAP7_75t_L g1878 ( 
.A(n_1824),
.B(n_1797),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1807),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1830),
.B(n_1746),
.Y(n_1880)
);

OAI21xp33_ASAP7_75t_L g1881 ( 
.A1(n_1838),
.A2(n_1742),
.B(n_1731),
.Y(n_1881)
);

OAI33xp33_ASAP7_75t_L g1882 ( 
.A1(n_1838),
.A2(n_1789),
.A3(n_1781),
.B1(n_1772),
.B2(n_1715),
.B3(n_1720),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1811),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1842),
.A2(n_1742),
.B1(n_1662),
.B2(n_1737),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1863),
.B(n_1812),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1863),
.B(n_1814),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1845),
.B(n_1806),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1845),
.B(n_1806),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1874),
.B(n_1814),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1879),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1856),
.B(n_1832),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1874),
.B(n_1819),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1860),
.B(n_1819),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1855),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1856),
.B(n_1832),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1858),
.B(n_1828),
.Y(n_1896)
);

AOI21xp33_ASAP7_75t_L g1897 ( 
.A1(n_1847),
.A2(n_1752),
.B(n_1747),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1845),
.B(n_1836),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1855),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1879),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1849),
.B(n_1850),
.Y(n_1901)
);

OR2x2_ASAP7_75t_L g1902 ( 
.A(n_1860),
.B(n_1803),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1858),
.B(n_1828),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1861),
.B(n_1868),
.Y(n_1904)
);

HB1xp67_ASAP7_75t_L g1905 ( 
.A(n_1853),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1853),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1851),
.Y(n_1907)
);

INVxp67_ASAP7_75t_L g1908 ( 
.A(n_1840),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1851),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1849),
.B(n_1839),
.Y(n_1910)
);

NAND2x1p5_ASAP7_75t_L g1911 ( 
.A(n_1841),
.B(n_1800),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1864),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1864),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1865),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1865),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1883),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1861),
.B(n_1803),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1868),
.B(n_1833),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1859),
.B(n_1825),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1870),
.B(n_1857),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1869),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1859),
.B(n_1829),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1901),
.B(n_1858),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1889),
.B(n_1867),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1889),
.B(n_1904),
.Y(n_1925)
);

AO21x2_ASAP7_75t_L g1926 ( 
.A1(n_1897),
.A2(n_1841),
.B(n_1870),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1901),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1890),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1890),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1901),
.B(n_1858),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1904),
.B(n_1867),
.Y(n_1931)
);

OAI21xp5_ASAP7_75t_SL g1932 ( 
.A1(n_1897),
.A2(n_1842),
.B(n_1847),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1908),
.B(n_1873),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1887),
.B(n_1873),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1892),
.B(n_1885),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1884),
.B(n_1843),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1894),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1887),
.B(n_1873),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1900),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1900),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1887),
.B(n_1873),
.Y(n_1941)
);

INVx2_ASAP7_75t_SL g1942 ( 
.A(n_1905),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1905),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1906),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_L g1945 ( 
.A(n_1885),
.B(n_1754),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1892),
.B(n_1843),
.Y(n_1946)
);

AO22x1_ASAP7_75t_L g1947 ( 
.A1(n_1906),
.A2(n_1799),
.B1(n_1794),
.B2(n_1750),
.Y(n_1947)
);

NAND4xp25_ASAP7_75t_L g1948 ( 
.A(n_1908),
.B(n_1848),
.C(n_1876),
.D(n_1846),
.Y(n_1948)
);

INVxp67_ASAP7_75t_SL g1949 ( 
.A(n_1920),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1886),
.B(n_1867),
.Y(n_1950)
);

NAND2x1p5_ASAP7_75t_L g1951 ( 
.A(n_1896),
.B(n_1857),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1888),
.B(n_1866),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1888),
.B(n_1866),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1907),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1907),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1893),
.B(n_1881),
.Y(n_1956)
);

INVxp67_ASAP7_75t_L g1957 ( 
.A(n_1920),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1909),
.Y(n_1958)
);

NAND2x1_ASAP7_75t_L g1959 ( 
.A(n_1896),
.B(n_1840),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1909),
.Y(n_1960)
);

AOI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1911),
.A2(n_1848),
.B(n_1872),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1894),
.Y(n_1962)
);

NAND2x1p5_ASAP7_75t_L g1963 ( 
.A(n_1896),
.B(n_1854),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1894),
.Y(n_1964)
);

INVxp67_ASAP7_75t_L g1965 ( 
.A(n_1917),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1886),
.B(n_1917),
.Y(n_1966)
);

INVx3_ASAP7_75t_L g1967 ( 
.A(n_1896),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1927),
.B(n_1919),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1942),
.B(n_1903),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1927),
.B(n_1919),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1952),
.B(n_1919),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1942),
.B(n_1903),
.Y(n_1972)
);

NAND4xp25_ASAP7_75t_L g1973 ( 
.A(n_1932),
.B(n_1876),
.C(n_1846),
.D(n_1881),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1952),
.B(n_1922),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_L g1975 ( 
.A(n_1936),
.B(n_1754),
.Y(n_1975)
);

INVx1_ASAP7_75t_SL g1976 ( 
.A(n_1947),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1953),
.B(n_1922),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1953),
.B(n_1922),
.Y(n_1978)
);

AND2x4_ASAP7_75t_SL g1979 ( 
.A(n_1933),
.B(n_1923),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1946),
.B(n_1893),
.Y(n_1980)
);

HB1xp67_ASAP7_75t_L g1981 ( 
.A(n_1943),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1923),
.B(n_1877),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1947),
.B(n_1902),
.Y(n_1983)
);

NAND4xp25_ASAP7_75t_SL g1984 ( 
.A(n_1961),
.B(n_1880),
.C(n_1877),
.D(n_1737),
.Y(n_1984)
);

NOR2x1_ASAP7_75t_L g1985 ( 
.A(n_1948),
.B(n_1903),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1928),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1925),
.B(n_1935),
.Y(n_1987)
);

BUFx2_ASAP7_75t_L g1988 ( 
.A(n_1963),
.Y(n_1988)
);

NOR2x1_ASAP7_75t_L g1989 ( 
.A(n_1926),
.B(n_1903),
.Y(n_1989)
);

OR2x2_ASAP7_75t_L g1990 ( 
.A(n_1925),
.B(n_1902),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1930),
.B(n_1877),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1935),
.B(n_1891),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1934),
.Y(n_1993)
);

INVx2_ASAP7_75t_SL g1994 ( 
.A(n_1959),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1929),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_L g1996 ( 
.A(n_1945),
.B(n_1739),
.Y(n_1996)
);

INVxp67_ASAP7_75t_SL g1997 ( 
.A(n_1959),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1957),
.B(n_1910),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1930),
.B(n_1899),
.Y(n_1999)
);

BUFx3_ASAP7_75t_L g2000 ( 
.A(n_1944),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1934),
.B(n_1880),
.Y(n_2001)
);

AND2x4_ASAP7_75t_L g2002 ( 
.A(n_1933),
.B(n_1899),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1939),
.Y(n_2003)
);

NAND2xp33_ASAP7_75t_L g2004 ( 
.A(n_1951),
.B(n_1911),
.Y(n_2004)
);

NAND2x1p5_ASAP7_75t_L g2005 ( 
.A(n_1967),
.B(n_1854),
.Y(n_2005)
);

NAND2xp33_ASAP7_75t_SL g2006 ( 
.A(n_1926),
.B(n_1875),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1986),
.Y(n_2007)
);

AOI322xp5_ASAP7_75t_L g2008 ( 
.A1(n_1985),
.A2(n_1976),
.A3(n_1975),
.B1(n_1983),
.B2(n_2006),
.C1(n_1980),
.C2(n_1949),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1985),
.B(n_1965),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_L g2010 ( 
.A(n_1996),
.B(n_1956),
.Y(n_2010)
);

AOI22xp33_ASAP7_75t_SL g2011 ( 
.A1(n_1997),
.A2(n_1926),
.B1(n_1911),
.B2(n_1735),
.Y(n_2011)
);

AOI21xp33_ASAP7_75t_L g2012 ( 
.A1(n_1987),
.A2(n_1911),
.B(n_1924),
.Y(n_2012)
);

OAI21xp33_ASAP7_75t_SL g2013 ( 
.A1(n_1989),
.A2(n_1973),
.B(n_1994),
.Y(n_2013)
);

OAI31xp33_ASAP7_75t_L g2014 ( 
.A1(n_1984),
.A2(n_1951),
.A3(n_1963),
.B(n_1933),
.Y(n_2014)
);

AOI21xp33_ASAP7_75t_L g2015 ( 
.A1(n_1987),
.A2(n_1924),
.B(n_1931),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1986),
.Y(n_2016)
);

OAI21xp5_ASAP7_75t_SL g2017 ( 
.A1(n_1979),
.A2(n_1951),
.B(n_1963),
.Y(n_2017)
);

AOI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1979),
.A2(n_1882),
.B1(n_1941),
.B2(n_1938),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1995),
.Y(n_2019)
);

AOI222xp33_ASAP7_75t_L g2020 ( 
.A1(n_2000),
.A2(n_1981),
.B1(n_2004),
.B2(n_1998),
.C1(n_1988),
.C2(n_1989),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1995),
.Y(n_2021)
);

OAI221xp5_ASAP7_75t_L g2022 ( 
.A1(n_2000),
.A2(n_1966),
.B1(n_1931),
.B2(n_1967),
.C(n_1950),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_2005),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_1990),
.B(n_1966),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1971),
.B(n_1938),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_2003),
.Y(n_2026)
);

OAI21xp5_ASAP7_75t_SL g2027 ( 
.A1(n_1988),
.A2(n_1831),
.B(n_1941),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1971),
.B(n_1940),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_2003),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1968),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1974),
.B(n_1954),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1974),
.B(n_1955),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1968),
.Y(n_2033)
);

OAI31xp33_ASAP7_75t_L g2034 ( 
.A1(n_2005),
.A2(n_1967),
.A3(n_1880),
.B(n_1950),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2010),
.B(n_1977),
.Y(n_2035)
);

OAI22xp33_ASAP7_75t_L g2036 ( 
.A1(n_2009),
.A2(n_1994),
.B1(n_2005),
.B2(n_1990),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_2025),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_2025),
.Y(n_2038)
);

AOI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_2013),
.A2(n_2010),
.B(n_2020),
.Y(n_2039)
);

INVxp67_ASAP7_75t_L g2040 ( 
.A(n_2024),
.Y(n_2040)
);

AOI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_2014),
.A2(n_1972),
.B(n_1969),
.Y(n_2041)
);

INVx2_ASAP7_75t_SL g2042 ( 
.A(n_2024),
.Y(n_2042)
);

AOI222xp33_ASAP7_75t_L g2043 ( 
.A1(n_2022),
.A2(n_2019),
.B1(n_2016),
.B2(n_2007),
.C1(n_2026),
.C2(n_2029),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_2023),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_L g2045 ( 
.A(n_2027),
.B(n_1992),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2021),
.Y(n_2046)
);

AOI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_2017),
.A2(n_1993),
.B1(n_1970),
.B2(n_1978),
.Y(n_2047)
);

OR4x1_ASAP7_75t_L g2048 ( 
.A(n_2030),
.B(n_2033),
.C(n_2021),
.D(n_2008),
.Y(n_2048)
);

NAND4xp25_ASAP7_75t_L g2049 ( 
.A(n_2011),
.B(n_1992),
.C(n_1993),
.D(n_1972),
.Y(n_2049)
);

OAI21xp33_ASAP7_75t_L g2050 ( 
.A1(n_2018),
.A2(n_1970),
.B(n_1977),
.Y(n_2050)
);

AOI222xp33_ASAP7_75t_L g2051 ( 
.A1(n_2028),
.A2(n_2032),
.B1(n_2031),
.B2(n_2023),
.C1(n_1882),
.C2(n_1969),
.Y(n_2051)
);

INVx2_ASAP7_75t_SL g2052 ( 
.A(n_2034),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2015),
.B(n_1978),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2012),
.Y(n_2054)
);

OAI21xp5_ASAP7_75t_L g2055 ( 
.A1(n_2013),
.A2(n_1972),
.B(n_1969),
.Y(n_2055)
);

OAI21xp33_ASAP7_75t_L g2056 ( 
.A1(n_2013),
.A2(n_1972),
.B(n_1969),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_2025),
.Y(n_2057)
);

OAI221xp5_ASAP7_75t_SL g2058 ( 
.A1(n_2039),
.A2(n_2001),
.B1(n_1991),
.B2(n_1982),
.C(n_1852),
.Y(n_2058)
);

XOR2x2_ASAP7_75t_L g2059 ( 
.A(n_2035),
.B(n_1735),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_2051),
.B(n_2002),
.Y(n_2060)
);

AOI22xp33_ASAP7_75t_L g2061 ( 
.A1(n_2052),
.A2(n_2002),
.B1(n_1999),
.B2(n_2001),
.Y(n_2061)
);

INVxp67_ASAP7_75t_L g2062 ( 
.A(n_2042),
.Y(n_2062)
);

OAI322xp33_ASAP7_75t_L g2063 ( 
.A1(n_2036),
.A2(n_1960),
.A3(n_1958),
.B1(n_1937),
.B2(n_1964),
.C1(n_1962),
.C2(n_1852),
.Y(n_2063)
);

NOR2xp33_ASAP7_75t_L g2064 ( 
.A(n_2040),
.B(n_2045),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2037),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_SL g2066 ( 
.A1(n_2048),
.A2(n_2002),
.B1(n_1999),
.B2(n_1991),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2038),
.Y(n_2067)
);

OAI21xp5_ASAP7_75t_L g2068 ( 
.A1(n_2051),
.A2(n_2002),
.B(n_1999),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2043),
.B(n_1999),
.Y(n_2069)
);

NOR3xp33_ASAP7_75t_L g2070 ( 
.A(n_2056),
.B(n_2054),
.C(n_2055),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_2053),
.B(n_1982),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2062),
.B(n_2043),
.Y(n_2072)
);

NOR2xp67_ASAP7_75t_L g2073 ( 
.A(n_2068),
.B(n_2049),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2061),
.B(n_2057),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_2065),
.Y(n_2075)
);

AOI21xp33_ASAP7_75t_SL g2076 ( 
.A1(n_2070),
.A2(n_2060),
.B(n_2069),
.Y(n_2076)
);

OAI211xp5_ASAP7_75t_L g2077 ( 
.A1(n_2066),
.A2(n_2055),
.B(n_2049),
.C(n_2041),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_2067),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_2071),
.B(n_2044),
.Y(n_2079)
);

AND4x1_ASAP7_75t_L g2080 ( 
.A(n_2064),
.B(n_2047),
.C(n_2046),
.D(n_2050),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_2058),
.B(n_1891),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_2066),
.B(n_1937),
.Y(n_2082)
);

AOI21xp5_ASAP7_75t_L g2083 ( 
.A1(n_2063),
.A2(n_1964),
.B(n_1962),
.Y(n_2083)
);

NAND4xp25_ASAP7_75t_SL g2084 ( 
.A(n_2059),
.B(n_1895),
.C(n_1918),
.D(n_1871),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2079),
.Y(n_2085)
);

INVxp67_ASAP7_75t_L g2086 ( 
.A(n_2072),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_SL g2087 ( 
.A(n_2073),
.B(n_1635),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_R g2088 ( 
.A(n_2074),
.B(n_1639),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_2077),
.A2(n_1747),
.B1(n_1740),
.B2(n_1831),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2075),
.Y(n_2090)
);

OAI211xp5_ASAP7_75t_L g2091 ( 
.A1(n_2076),
.A2(n_1691),
.B(n_1719),
.C(n_1724),
.Y(n_2091)
);

NAND4xp25_ASAP7_75t_L g2092 ( 
.A(n_2087),
.B(n_2076),
.C(n_2078),
.D(n_2082),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2085),
.Y(n_2093)
);

INVx1_ASAP7_75t_SL g2094 ( 
.A(n_2088),
.Y(n_2094)
);

AO22x2_ASAP7_75t_L g2095 ( 
.A1(n_2086),
.A2(n_2080),
.B1(n_2081),
.B2(n_2083),
.Y(n_2095)
);

OAI211xp5_ASAP7_75t_SL g2096 ( 
.A1(n_2091),
.A2(n_2084),
.B(n_1724),
.C(n_1715),
.Y(n_2096)
);

OAI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_2089),
.A2(n_1875),
.B1(n_1918),
.B2(n_1895),
.Y(n_2097)
);

NOR3xp33_ASAP7_75t_L g2098 ( 
.A(n_2090),
.B(n_1691),
.C(n_1740),
.Y(n_2098)
);

NOR3xp33_ASAP7_75t_L g2099 ( 
.A(n_2086),
.B(n_1691),
.C(n_1662),
.Y(n_2099)
);

AND3x4_ASAP7_75t_L g2100 ( 
.A(n_2099),
.B(n_1878),
.C(n_1844),
.Y(n_2100)
);

AO22x2_ASAP7_75t_L g2101 ( 
.A1(n_2093),
.A2(n_1899),
.B1(n_1916),
.B2(n_1875),
.Y(n_2101)
);

NOR2x1_ASAP7_75t_L g2102 ( 
.A(n_2092),
.B(n_1916),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_2094),
.B(n_1898),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2095),
.Y(n_2104)
);

NOR2x1_ASAP7_75t_L g2105 ( 
.A(n_2096),
.B(n_1916),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2103),
.B(n_2098),
.Y(n_2106)
);

AOI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_2104),
.A2(n_2097),
.B1(n_1639),
.B2(n_1844),
.Y(n_2107)
);

NAND3xp33_ASAP7_75t_L g2108 ( 
.A(n_2102),
.B(n_1720),
.C(n_1716),
.Y(n_2108)
);

A2O1A1Ixp33_ASAP7_75t_L g2109 ( 
.A1(n_2105),
.A2(n_1921),
.B(n_1912),
.C(n_1915),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2106),
.Y(n_2110)
);

XNOR2xp5_ASAP7_75t_L g2111 ( 
.A(n_2107),
.B(n_2100),
.Y(n_2111)
);

AO22x1_ASAP7_75t_L g2112 ( 
.A1(n_2110),
.A2(n_2101),
.B1(n_2108),
.B2(n_2109),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2111),
.Y(n_2113)
);

OAI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_2113),
.A2(n_1639),
.B1(n_1912),
.B2(n_1915),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2112),
.Y(n_2115)
);

OAI22x1_ASAP7_75t_L g2116 ( 
.A1(n_2115),
.A2(n_1716),
.B1(n_1710),
.B2(n_1718),
.Y(n_2116)
);

INVxp67_ASAP7_75t_SL g2117 ( 
.A(n_2114),
.Y(n_2117)
);

OA21x2_ASAP7_75t_L g2118 ( 
.A1(n_2117),
.A2(n_2116),
.B(n_1914),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2117),
.Y(n_2119)
);

OAI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_2119),
.A2(n_1921),
.B1(n_1913),
.B2(n_1914),
.Y(n_2120)
);

OAI21xp33_ASAP7_75t_L g2121 ( 
.A1(n_2120),
.A2(n_2118),
.B(n_1698),
.Y(n_2121)
);

OAI22xp33_ASAP7_75t_L g2122 ( 
.A1(n_2121),
.A2(n_2118),
.B1(n_1698),
.B2(n_1639),
.Y(n_2122)
);

AOI221xp5_ASAP7_75t_L g2123 ( 
.A1(n_2122),
.A2(n_2118),
.B1(n_1913),
.B2(n_1855),
.C(n_1862),
.Y(n_2123)
);

AOI211xp5_ASAP7_75t_L g2124 ( 
.A1(n_2123),
.A2(n_1717),
.B(n_1725),
.C(n_1710),
.Y(n_2124)
);


endmodule