module fake_jpeg_1195_n_207 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_207);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_207;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_4),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_14),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_66),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_57),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_23),
.C(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_57),
.Y(n_94)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_85),
.B(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_60),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_89),
.Y(n_98)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_93),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_64),
.B1(n_71),
.B2(n_50),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_89),
.B1(n_73),
.B2(n_65),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_66),
.Y(n_99)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_95),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_53),
.B1(n_71),
.B2(n_64),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_106),
.B1(n_108),
.B2(n_113),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_83),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_69),
.B1(n_66),
.B2(n_61),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_110),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_72),
.B1(n_56),
.B2(n_69),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_58),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_89),
.B1(n_90),
.B2(n_70),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_120),
.B1(n_125),
.B2(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_127),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_112),
.C(n_97),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_124),
.C(n_67),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_70),
.B1(n_51),
.B2(n_62),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_87),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_100),
.A2(n_68),
.B1(n_63),
.B2(n_95),
.Y(n_125)
);

BUFx2_ASAP7_75t_SL g126 ( 
.A(n_111),
.Y(n_126)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_0),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_128),
.B(n_131),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_1),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_134),
.Y(n_145)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_1),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_147),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_96),
.B(n_87),
.Y(n_140)
);

NAND3xp33_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_141),
.C(n_143),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_73),
.B(n_55),
.Y(n_141)
);

XOR2x2_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_67),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_157),
.C(n_12),
.Y(n_167)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_24),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_154),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_55),
.B1(n_3),
.B2(n_5),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_152),
.B1(n_153),
.B2(n_158),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_116),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_123),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_32),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_55),
.B1(n_3),
.B2(n_5),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_114),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_122),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_2),
.B(n_8),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_29),
.B(n_46),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_33),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_26),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_115),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_158)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_167),
.B(n_172),
.Y(n_177)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_13),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_171),
.B(n_175),
.Y(n_183)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_173),
.B(n_174),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_31),
.B(n_45),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_SL g175 ( 
.A1(n_155),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.C1(n_17),
.C2(n_18),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_176),
.A2(n_139),
.B1(n_141),
.B2(n_140),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_184),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_SL g182 ( 
.A(n_161),
.B(n_166),
.C(n_160),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_162),
.C(n_170),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_161),
.A2(n_156),
.B1(n_144),
.B2(n_139),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_167),
.B(n_157),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_39),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_159),
.A3(n_172),
.B1(n_163),
.B2(n_162),
.C1(n_170),
.C2(n_176),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_179),
.B(n_177),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_185),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_188),
.B(n_189),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_192),
.C(n_178),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_40),
.C(n_25),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_178),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_193),
.Y(n_198)
);

NOR2xp67_ASAP7_75t_SL g199 ( 
.A(n_194),
.B(n_190),
.Y(n_199)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_195),
.A2(n_180),
.B1(n_187),
.B2(n_19),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_183),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_198),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_196),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_203),
.A2(n_197),
.B(n_34),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_204),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_36),
.B1(n_41),
.B2(n_43),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_49),
.Y(n_207)
);


endmodule