module real_aes_9270_n_329 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_329);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_329;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_602;
wire n_402;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_1185;
wire n_661;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_1457;
wire n_719;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1679;
wire n_460;
wire n_1595;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1025;
wire n_532;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1678;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_1369;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_0), .A2(n_142), .B1(n_523), .B2(n_663), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_0), .A2(n_142), .B1(n_538), .B2(n_640), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_1), .A2(n_77), .B1(n_688), .B2(n_1202), .Y(n_1201) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1), .Y(n_1209) );
INVxp33_ASAP7_75t_L g776 ( .A(n_2), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g814 ( .A1(n_2), .A2(n_753), .B(n_815), .Y(n_814) );
INVxp67_ASAP7_75t_SL g1272 ( .A(n_3), .Y(n_1272) );
AOI22xp33_ASAP7_75t_L g1288 ( .A1(n_3), .A2(n_8), .B1(n_647), .B2(n_1289), .Y(n_1288) );
AOI22xp33_ASAP7_75t_L g1284 ( .A1(n_4), .A2(n_209), .B1(n_543), .B2(n_672), .Y(n_1284) );
AOI22xp33_ASAP7_75t_L g1295 ( .A1(n_4), .A2(n_209), .B1(n_493), .B2(n_1296), .Y(n_1295) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_5), .A2(n_150), .B1(n_493), .B2(n_915), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g962 ( .A1(n_5), .A2(n_150), .B1(n_614), .B2(n_618), .Y(n_962) );
INVx1_ASAP7_75t_L g1264 ( .A(n_6), .Y(n_1264) );
INVx1_ASAP7_75t_L g1181 ( .A(n_7), .Y(n_1181) );
AOI22xp33_ASAP7_75t_L g1191 ( .A1(n_7), .A2(n_233), .B1(n_647), .B2(n_1192), .Y(n_1191) );
INVx1_ASAP7_75t_L g1271 ( .A(n_8), .Y(n_1271) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_9), .A2(n_265), .B1(n_472), .B2(n_742), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_9), .A2(n_265), .B1(n_760), .B2(n_761), .Y(n_759) );
INVx1_ASAP7_75t_L g1420 ( .A(n_10), .Y(n_1420) );
CKINVDCx5p33_ASAP7_75t_R g1023 ( .A(n_11), .Y(n_1023) );
AOI22xp33_ASAP7_75t_SL g1109 ( .A1(n_12), .A2(n_272), .B1(n_915), .B2(n_1110), .Y(n_1109) );
INVxp67_ASAP7_75t_L g1119 ( .A(n_12), .Y(n_1119) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_13), .A2(n_200), .B1(n_540), .B2(n_541), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_13), .A2(n_200), .B1(n_492), .B2(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g738 ( .A(n_14), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_14), .A2(n_51), .B1(n_744), .B2(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g1263 ( .A(n_15), .Y(n_1263) );
AOI22xp33_ASAP7_75t_L g1291 ( .A1(n_15), .A2(n_61), .B1(n_959), .B2(n_1286), .Y(n_1291) );
INVx1_ASAP7_75t_L g524 ( .A(n_16), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_16), .A2(n_220), .B1(n_432), .B2(n_577), .Y(n_576) );
INVxp33_ASAP7_75t_SL g729 ( .A(n_17), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_17), .A2(n_88), .B1(n_563), .B2(n_765), .Y(n_764) );
AO221x2_ASAP7_75t_L g1418 ( .A1(n_18), .A2(n_245), .B1(n_1395), .B2(n_1417), .C(n_1419), .Y(n_1418) );
INVx1_ASAP7_75t_L g1355 ( .A(n_19), .Y(n_1355) );
OAI22xp5_ASAP7_75t_L g1368 ( .A1(n_19), .A2(n_295), .B1(n_605), .B2(n_610), .Y(n_1368) );
CKINVDCx16_ASAP7_75t_R g1439 ( .A(n_20), .Y(n_1439) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_21), .A2(n_323), .B1(n_523), .B2(n_663), .Y(n_1200) );
INVx1_ASAP7_75t_L g1206 ( .A(n_21), .Y(n_1206) );
INVx1_ASAP7_75t_L g1654 ( .A(n_22), .Y(n_1654) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_23), .A2(n_69), .B1(n_545), .B2(n_889), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_23), .A2(n_69), .B1(n_904), .B2(n_907), .Y(n_903) );
OAI211xp5_ASAP7_75t_L g972 ( .A1(n_24), .A2(n_407), .B(n_847), .C(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g991 ( .A(n_24), .Y(n_991) );
INVx1_ASAP7_75t_L g868 ( .A(n_25), .Y(n_868) );
INVx1_ASAP7_75t_L g1322 ( .A(n_26), .Y(n_1322) );
AOI22xp33_ASAP7_75t_SL g1335 ( .A1(n_26), .A2(n_179), .B1(n_915), .B2(n_916), .Y(n_1335) );
CKINVDCx5p33_ASAP7_75t_R g1074 ( .A(n_27), .Y(n_1074) );
INVx1_ASAP7_75t_L g1095 ( .A(n_28), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g1116 ( .A1(n_28), .A2(n_30), .B1(n_432), .B2(n_577), .Y(n_1116) );
CKINVDCx5p33_ASAP7_75t_R g1002 ( .A(n_29), .Y(n_1002) );
INVx1_ASAP7_75t_L g1096 ( .A(n_30), .Y(n_1096) );
INVx1_ASAP7_75t_L g1648 ( .A(n_31), .Y(n_1648) );
CKINVDCx5p33_ASAP7_75t_R g1075 ( .A(n_32), .Y(n_1075) );
INVx1_ASAP7_75t_L g1033 ( .A(n_33), .Y(n_1033) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_33), .A2(n_165), .B1(n_614), .B2(n_618), .Y(n_1076) );
INVx1_ASAP7_75t_L g725 ( .A(n_34), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_35), .A2(n_317), .B1(n_569), .B2(n_570), .Y(n_568) );
INVxp67_ASAP7_75t_SL g580 ( .A(n_35), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_36), .A2(n_99), .B1(n_440), .B2(n_474), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_36), .A2(n_99), .B1(n_502), .B2(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g335 ( .A(n_37), .Y(n_335) );
XNOR2xp5_ASAP7_75t_L g1013 ( .A(n_38), .B(n_1014), .Y(n_1013) );
AOI221xp5_ASAP7_75t_L g933 ( .A1(n_39), .A2(n_213), .B1(n_540), .B2(n_548), .C(n_934), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_39), .A2(n_213), .B1(n_915), .B2(n_916), .Y(n_950) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_40), .A2(n_59), .B1(n_344), .B2(n_416), .Y(n_703) );
OAI22xp33_ASAP7_75t_L g714 ( .A1(n_40), .A2(n_312), .B1(n_605), .B2(n_610), .Y(n_714) );
INVxp67_ASAP7_75t_L g449 ( .A(n_41), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_41), .A2(n_255), .B1(n_502), .B2(n_503), .Y(n_501) );
INVxp67_ASAP7_75t_SL g602 ( .A(n_42), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_42), .A2(n_172), .B1(n_647), .B2(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g1098 ( .A(n_43), .Y(n_1098) );
OAI22xp5_ASAP7_75t_L g1142 ( .A1(n_44), .A2(n_101), .B1(n_605), .B2(n_930), .Y(n_1142) );
AOI22xp33_ASAP7_75t_SL g1161 ( .A1(n_44), .A2(n_101), .B1(n_535), .B2(n_742), .Y(n_1161) );
INVxp67_ASAP7_75t_SL g404 ( .A(n_45), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_45), .A2(n_328), .B1(n_432), .B2(n_435), .Y(n_431) );
AOI22xp33_ASAP7_75t_SL g533 ( .A1(n_46), .A2(n_168), .B1(n_534), .B2(n_536), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_46), .A2(n_168), .B1(n_561), .B2(n_563), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_47), .A2(n_313), .B1(n_1157), .B2(n_1159), .Y(n_1156) );
AOI22xp33_ASAP7_75t_SL g1168 ( .A1(n_47), .A2(n_214), .B1(n_761), .B2(n_1169), .Y(n_1168) );
INVxp67_ASAP7_75t_SL g736 ( .A(n_48), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_48), .A2(n_261), .B1(n_742), .B2(n_747), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_49), .A2(n_281), .B1(n_672), .B2(n_673), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_49), .A2(n_281), .B1(n_559), .B2(n_684), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g1326 ( .A1(n_50), .A2(n_175), .B1(n_675), .B2(n_959), .Y(n_1326) );
AOI22xp33_ASAP7_75t_L g1331 ( .A1(n_50), .A2(n_175), .B1(n_523), .B2(n_663), .Y(n_1331) );
INVxp33_ASAP7_75t_SL g733 ( .A(n_51), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_52), .A2(n_74), .B1(n_614), .B2(n_618), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_52), .A2(n_74), .B1(n_492), .B2(n_559), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g1445 ( .A1(n_53), .A2(n_296), .B1(n_1395), .B2(n_1417), .Y(n_1445) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_54), .A2(n_56), .B1(n_461), .B2(n_465), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_54), .A2(n_56), .B1(n_486), .B2(n_488), .Y(n_485) );
INVxp67_ASAP7_75t_SL g864 ( .A(n_55), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_55), .A2(n_65), .B1(n_913), .B2(n_916), .Y(n_912) );
INVxp33_ASAP7_75t_SL g1149 ( .A(n_57), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_57), .A2(n_146), .B1(n_760), .B2(n_761), .Y(n_1171) );
INVxp67_ASAP7_75t_SL g1224 ( .A(n_58), .Y(n_1224) );
AOI22xp33_ASAP7_75t_L g1234 ( .A1(n_58), .A2(n_198), .B1(n_548), .B2(n_896), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_59), .A2(n_159), .B1(n_691), .B2(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g952 ( .A(n_60), .Y(n_952) );
INVx1_ASAP7_75t_L g1266 ( .A(n_61), .Y(n_1266) );
INVx1_ASAP7_75t_L g1275 ( .A(n_62), .Y(n_1275) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_62), .A2(n_226), .B1(n_396), .B2(n_500), .Y(n_1298) );
OAI211xp5_ASAP7_75t_L g923 ( .A1(n_63), .A2(n_407), .B(n_924), .C(n_926), .Y(n_923) );
INVx1_ASAP7_75t_L g944 ( .A(n_63), .Y(n_944) );
XNOR2xp5_ASAP7_75t_L g1173 ( .A(n_64), .B(n_1174), .Y(n_1173) );
INVxp67_ASAP7_75t_SL g874 ( .A(n_65), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_66), .A2(n_124), .B1(n_455), .B2(n_457), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_66), .A2(n_124), .B1(n_491), .B2(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g1646 ( .A(n_67), .Y(n_1646) );
INVx1_ASAP7_75t_L g701 ( .A(n_68), .Y(n_701) );
CKINVDCx5p33_ASAP7_75t_R g1372 ( .A(n_70), .Y(n_1372) );
INVxp67_ASAP7_75t_SL g787 ( .A(n_71), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_71), .A2(n_249), .B1(n_502), .B2(n_851), .Y(n_850) );
XOR2xp5_ASAP7_75t_L g1130 ( .A(n_72), .B(n_1131), .Y(n_1130) );
INVx1_ASAP7_75t_L g1137 ( .A(n_73), .Y(n_1137) );
OAI222xp33_ASAP7_75t_L g1146 ( .A1(n_73), .A2(n_156), .B1(n_247), .B2(n_577), .C1(n_813), .C2(n_870), .Y(n_1146) );
AOI221xp5_ASAP7_75t_L g996 ( .A1(n_75), .A2(n_234), .B1(n_455), .B2(n_997), .C(n_999), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_75), .A2(n_234), .B1(n_906), .B2(n_916), .Y(n_1006) );
OAI21xp33_ASAP7_75t_SL g1135 ( .A1(n_76), .A2(n_1020), .B(n_1136), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_76), .A2(n_275), .B1(n_465), .B2(n_648), .Y(n_1162) );
INVx1_ASAP7_75t_L g1210 ( .A(n_77), .Y(n_1210) );
CKINVDCx5p33_ASAP7_75t_R g1177 ( .A(n_78), .Y(n_1177) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_79), .A2(n_222), .B1(n_614), .B2(n_618), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_79), .A2(n_222), .B1(n_493), .B2(n_906), .Y(n_1010) );
BUFx2_ASAP7_75t_L g361 ( .A(n_80), .Y(n_361) );
BUFx2_ASAP7_75t_L g451 ( .A(n_80), .Y(n_451) );
INVx1_ASAP7_75t_L g481 ( .A(n_80), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_81), .A2(n_165), .B1(n_1035), .B2(n_1037), .Y(n_1034) );
OAI211xp5_ASAP7_75t_L g1071 ( .A1(n_81), .A2(n_624), .B(n_1072), .C(n_1073), .Y(n_1071) );
INVx1_ASAP7_75t_L g521 ( .A(n_82), .Y(n_521) );
AOI22xp33_ASAP7_75t_SL g549 ( .A1(n_82), .A2(n_173), .B1(n_534), .B2(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_83), .A2(n_293), .B1(n_643), .B2(n_675), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_83), .A2(n_293), .B1(n_523), .B2(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g1308 ( .A(n_84), .Y(n_1308) );
AOI22xp33_ASAP7_75t_L g1328 ( .A1(n_84), .A2(n_321), .B1(n_543), .B2(n_547), .Y(n_1328) );
XNOR2xp5_ASAP7_75t_L g591 ( .A(n_85), .B(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_86), .A2(n_284), .B1(n_534), .B2(n_643), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_86), .A2(n_284), .B1(n_565), .B2(n_692), .Y(n_902) );
CKINVDCx5p33_ASAP7_75t_R g982 ( .A(n_87), .Y(n_982) );
INVx1_ASAP7_75t_L g724 ( .A(n_88), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_89), .A2(n_319), .B1(n_682), .B2(n_692), .Y(n_1108) );
INVxp33_ASAP7_75t_L g1121 ( .A(n_89), .Y(n_1121) );
OAI22xp33_ASAP7_75t_L g929 ( .A1(n_90), .A2(n_224), .B1(n_930), .B2(n_931), .Y(n_929) );
AOI221xp5_ASAP7_75t_L g939 ( .A1(n_90), .A2(n_224), .B1(n_545), .B2(n_897), .C(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g1067 ( .A(n_91), .Y(n_1067) );
OAI211xp5_ASAP7_75t_SL g1080 ( .A1(n_91), .A2(n_528), .B(n_1081), .C(n_1083), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_92), .A2(n_214), .B1(n_1152), .B2(n_1154), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_92), .A2(n_313), .B1(n_1165), .B2(n_1167), .Y(n_1164) );
INVx1_ASAP7_75t_L g1679 ( .A(n_93), .Y(n_1679) );
OAI22xp5_ASAP7_75t_L g1312 ( .A1(n_94), .A2(n_100), .B1(n_1269), .B2(n_1313), .Y(n_1312) );
OAI22xp5_ASAP7_75t_L g1317 ( .A1(n_94), .A2(n_100), .B1(n_435), .B2(n_627), .Y(n_1317) );
CKINVDCx16_ASAP7_75t_R g1441 ( .A(n_95), .Y(n_1441) );
INVx1_ASAP7_75t_L g715 ( .A(n_96), .Y(n_715) );
INVx1_ASAP7_75t_L g935 ( .A(n_97), .Y(n_935) );
INVx1_ASAP7_75t_L g1672 ( .A(n_98), .Y(n_1672) );
CKINVDCx5p33_ASAP7_75t_R g1000 ( .A(n_102), .Y(n_1000) );
INVx1_ASAP7_75t_L g1657 ( .A(n_103), .Y(n_1657) );
OAI22xp33_ASAP7_75t_SL g1685 ( .A1(n_103), .A2(n_202), .B1(n_344), .B2(n_614), .Y(n_1685) );
AO22x2_ASAP7_75t_L g1085 ( .A1(n_104), .A2(n_1086), .B1(n_1123), .B2(n_1124), .Y(n_1085) );
INVx1_ASAP7_75t_L g1123 ( .A(n_104), .Y(n_1123) );
INVx1_ASAP7_75t_L g928 ( .A(n_105), .Y(n_928) );
AOI22xp5_ASAP7_75t_L g1416 ( .A1(n_106), .A2(n_292), .B1(n_1395), .B2(n_1417), .Y(n_1416) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_107), .A2(n_228), .B1(n_488), .B2(n_565), .Y(n_1240) );
INVxp67_ASAP7_75t_SL g1246 ( .A(n_107), .Y(n_1246) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_108), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_108), .A2(n_270), .B1(n_488), .B2(n_500), .Y(n_499) );
XOR2xp5_ASAP7_75t_L g1339 ( .A(n_109), .B(n_1340), .Y(n_1339) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_110), .A2(n_279), .B1(n_906), .B2(n_916), .Y(n_1102) );
AOI22xp33_ASAP7_75t_SL g1111 ( .A1(n_110), .A2(n_279), .B1(n_543), .B2(n_672), .Y(n_1111) );
INVx1_ASAP7_75t_L g1180 ( .A(n_111), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1193 ( .A1(n_111), .A2(n_236), .B1(n_643), .B2(n_651), .Y(n_1193) );
INVx1_ASAP7_75t_L g1228 ( .A(n_112), .Y(n_1228) );
OAI22xp5_ASAP7_75t_L g1247 ( .A1(n_112), .A2(n_273), .B1(n_432), .B2(n_577), .Y(n_1247) );
INVxp33_ASAP7_75t_L g877 ( .A(n_113), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_113), .A2(n_163), .B1(n_534), .B2(n_900), .Y(n_899) );
AOI22xp5_ASAP7_75t_L g1455 ( .A1(n_114), .A2(n_117), .B1(n_1411), .B2(n_1414), .Y(n_1455) );
INVxp67_ASAP7_75t_SL g1092 ( .A(n_115), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_115), .A2(n_197), .B1(n_538), .B2(n_675), .Y(n_1105) );
INVx1_ASAP7_75t_L g1668 ( .A(n_116), .Y(n_1668) );
OAI22xp33_ASAP7_75t_L g1674 ( .A1(n_116), .A2(n_125), .B1(n_605), .B2(n_930), .Y(n_1674) );
XNOR2xp5_ASAP7_75t_L g355 ( .A(n_117), .B(n_356), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g1456 ( .A1(n_118), .A2(n_309), .B1(n_1389), .B2(n_1457), .Y(n_1456) );
INVx1_ASAP7_75t_L g863 ( .A(n_119), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_120), .A2(n_191), .B1(n_1025), .B2(n_1027), .Y(n_1024) );
INVx1_ASAP7_75t_L g1051 ( .A(n_120), .Y(n_1051) );
INVx1_ASAP7_75t_L g1353 ( .A(n_121), .Y(n_1353) );
OAI22xp5_ASAP7_75t_L g1374 ( .A1(n_121), .A2(n_263), .B1(n_930), .B2(n_931), .Y(n_1374) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_122), .A2(n_718), .B1(n_770), .B2(n_771), .Y(n_717) );
INVxp67_ASAP7_75t_L g770 ( .A(n_122), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g1145 ( .A1(n_123), .A2(n_160), .B1(n_344), .B2(n_416), .Y(n_1145) );
AOI22xp33_ASAP7_75t_SL g1170 ( .A1(n_123), .A2(n_247), .B1(n_486), .B2(n_1167), .Y(n_1170) );
INVx1_ASAP7_75t_L g1671 ( .A(n_125), .Y(n_1671) );
INVxp33_ASAP7_75t_SL g1090 ( .A(n_126), .Y(n_1090) );
AOI22xp33_ASAP7_75t_SL g1104 ( .A1(n_126), .A2(n_287), .B1(n_543), .B2(n_672), .Y(n_1104) );
AO221x2_ASAP7_75t_L g1388 ( .A1(n_127), .A2(n_188), .B1(n_1389), .B2(n_1395), .C(n_1396), .Y(n_1388) );
INVx1_ASAP7_75t_L g1394 ( .A(n_128), .Y(n_1394) );
OAI211xp5_ASAP7_75t_L g619 ( .A1(n_129), .A2(n_620), .B(n_624), .C(n_625), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_129), .A2(n_232), .B1(n_655), .B2(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g1540 ( .A(n_130), .Y(n_1540) );
INVxp33_ASAP7_75t_SL g1220 ( .A(n_131), .Y(n_1220) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_131), .A2(n_169), .B1(n_534), .B2(n_550), .Y(n_1235) );
CKINVDCx5p33_ASAP7_75t_R g1306 ( .A(n_132), .Y(n_1306) );
XOR2x2_ASAP7_75t_L g510 ( .A(n_133), .B(n_511), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_134), .A2(n_208), .B1(n_636), .B2(n_637), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_134), .A2(n_208), .B1(n_492), .B2(n_559), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g1285 ( .A1(n_135), .A2(n_221), .B1(n_422), .B2(n_1286), .Y(n_1285) );
AOI22xp33_ASAP7_75t_L g1293 ( .A1(n_135), .A2(n_221), .B1(n_1037), .B2(n_1294), .Y(n_1293) );
XNOR2xp5_ASAP7_75t_L g772 ( .A(n_136), .B(n_773), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g1444 ( .A1(n_136), .A2(n_320), .B1(n_1411), .B2(n_1414), .Y(n_1444) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_137), .Y(n_866) );
INVx1_ASAP7_75t_L g1357 ( .A(n_138), .Y(n_1357) );
AO22x2_ASAP7_75t_SL g1215 ( .A1(n_139), .A2(n_1216), .B1(n_1217), .B2(n_1253), .Y(n_1215) );
CKINVDCx16_ASAP7_75t_R g1216 ( .A(n_139), .Y(n_1216) );
INVx1_ASAP7_75t_L g1364 ( .A(n_140), .Y(n_1364) );
OAI22xp33_ASAP7_75t_SL g1379 ( .A1(n_140), .A2(n_148), .B1(n_344), .B2(n_614), .Y(n_1379) );
INVx1_ASAP7_75t_L g1392 ( .A(n_141), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1405 ( .A(n_141), .B(n_1402), .Y(n_1405) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_143), .A2(n_206), .B1(n_538), .B2(n_640), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_143), .A2(n_206), .B1(n_523), .B2(n_663), .Y(n_1195) );
OAI22xp5_ASAP7_75t_L g970 ( .A1(n_144), .A2(n_154), .B1(n_605), .B2(n_930), .Y(n_970) );
AOI221xp5_ASAP7_75t_L g986 ( .A1(n_144), .A2(n_276), .B1(n_545), .B2(n_987), .C(n_989), .Y(n_986) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_145), .Y(n_387) );
AOI22xp33_ASAP7_75t_SL g471 ( .A1(n_145), .A2(n_203), .B1(n_455), .B2(n_472), .Y(n_471) );
INVxp33_ASAP7_75t_L g1148 ( .A(n_146), .Y(n_1148) );
INVx2_ASAP7_75t_L g347 ( .A(n_147), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_148), .A2(n_258), .B1(n_493), .B2(n_559), .Y(n_1366) );
AOI22xp33_ASAP7_75t_SL g564 ( .A1(n_149), .A2(n_277), .B1(n_565), .B2(n_567), .Y(n_564) );
INVxp33_ASAP7_75t_SL g582 ( .A(n_149), .Y(n_582) );
BUFx3_ASAP7_75t_L g373 ( .A(n_151), .Y(n_373) );
INVx1_ASAP7_75t_L g391 ( .A(n_151), .Y(n_391) );
INVx1_ASAP7_75t_L g782 ( .A(n_152), .Y(n_782) );
INVx1_ASAP7_75t_L g1397 ( .A(n_153), .Y(n_1397) );
INVx1_ASAP7_75t_L g990 ( .A(n_154), .Y(n_990) );
AOI22xp33_ASAP7_75t_SL g1325 ( .A1(n_155), .A2(n_216), .B1(n_543), .B2(n_672), .Y(n_1325) );
AOI22xp33_ASAP7_75t_SL g1332 ( .A1(n_155), .A2(n_216), .B1(n_493), .B2(n_915), .Y(n_1332) );
INVx1_ASAP7_75t_L g1138 ( .A(n_156), .Y(n_1138) );
INVx1_ASAP7_75t_L g1305 ( .A(n_157), .Y(n_1305) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_157), .A2(n_278), .B1(n_675), .B2(n_959), .Y(n_1329) );
INVxp33_ASAP7_75t_L g872 ( .A(n_158), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_158), .A2(n_219), .B1(n_394), .B2(n_565), .Y(n_917) );
OAI211xp5_ASAP7_75t_SL g696 ( .A1(n_159), .A2(n_624), .B(n_697), .C(n_700), .Y(n_696) );
INVx1_ASAP7_75t_L g1140 ( .A(n_160), .Y(n_1140) );
INVxp33_ASAP7_75t_L g777 ( .A(n_161), .Y(n_777) );
AOI221xp5_ASAP7_75t_L g811 ( .A1(n_161), .A2(n_268), .B1(n_636), .B2(n_648), .C(n_812), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g1233 ( .A1(n_162), .A2(n_211), .B1(n_545), .B2(n_987), .Y(n_1233) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_162), .A2(n_211), .B1(n_761), .B2(n_1238), .Y(n_1237) );
INVx1_ASAP7_75t_L g882 ( .A(n_163), .Y(n_882) );
INVx1_ASAP7_75t_L g1538 ( .A(n_164), .Y(n_1538) );
AOI22xp33_ASAP7_75t_SL g1232 ( .A1(n_166), .A2(n_322), .B1(n_534), .B2(n_536), .Y(n_1232) );
AOI22xp33_ASAP7_75t_SL g1239 ( .A1(n_166), .A2(n_322), .B1(n_486), .B2(n_567), .Y(n_1239) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_167), .A2(n_312), .B1(n_640), .B2(n_643), .Y(n_679) );
INVx1_ASAP7_75t_L g707 ( .A(n_167), .Y(n_707) );
INVx1_ASAP7_75t_L g1226 ( .A(n_169), .Y(n_1226) );
INVx1_ASAP7_75t_L g393 ( .A(n_170), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_170), .A2(n_177), .B1(n_461), .B2(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g600 ( .A(n_171), .Y(n_600) );
INVx1_ASAP7_75t_L g603 ( .A(n_172), .Y(n_603) );
INVxp33_ASAP7_75t_SL g514 ( .A(n_173), .Y(n_514) );
XNOR2xp5_ASAP7_75t_L g967 ( .A(n_174), .B(n_968), .Y(n_967) );
INVx1_ASAP7_75t_L g1403 ( .A(n_174), .Y(n_1403) );
INVx1_ASAP7_75t_L g1658 ( .A(n_176), .Y(n_1658) );
OAI211xp5_ASAP7_75t_SL g1683 ( .A1(n_176), .A2(n_620), .B(n_624), .C(n_1684), .Y(n_1683) );
INVxp33_ASAP7_75t_SL g364 ( .A(n_177), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_178), .A2(n_259), .B1(n_605), .B2(n_610), .Y(n_922) );
INVx1_ASAP7_75t_L g961 ( .A(n_178), .Y(n_961) );
INVx1_ASAP7_75t_L g1320 ( .A(n_179), .Y(n_1320) );
INVx1_ASAP7_75t_L g359 ( .A(n_180), .Y(n_359) );
INVx1_ASAP7_75t_L g702 ( .A(n_181), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_182), .A2(n_185), .B1(n_535), .B2(n_744), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_182), .A2(n_185), .B1(n_488), .B2(n_756), .Y(n_755) );
INVxp67_ASAP7_75t_L g1281 ( .A(n_183), .Y(n_1281) );
AOI22xp33_ASAP7_75t_L g1299 ( .A1(n_183), .A2(n_264), .B1(n_915), .B2(n_916), .Y(n_1299) );
INVx1_ASAP7_75t_L g1185 ( .A(n_184), .Y(n_1185) );
OAI22xp33_ASAP7_75t_L g1207 ( .A1(n_184), .A2(n_298), .B1(n_577), .B2(n_870), .Y(n_1207) );
INVxp67_ASAP7_75t_SL g1349 ( .A(n_186), .Y(n_1349) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_186), .A2(n_302), .B1(n_493), .B2(n_688), .Y(n_1362) );
INVx1_ASAP7_75t_L g1428 ( .A(n_187), .Y(n_1428) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_189), .A2(n_318), .B1(n_543), .B2(n_672), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_189), .A2(n_318), .B1(n_689), .B2(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1062 ( .A(n_190), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_190), .A2(n_192), .B1(n_605), .B2(n_930), .Y(n_1078) );
INVx1_ASAP7_75t_L g1045 ( .A(n_191), .Y(n_1045) );
INVx1_ASAP7_75t_L g1058 ( .A(n_192), .Y(n_1058) );
CKINVDCx14_ASAP7_75t_R g919 ( .A(n_193), .Y(n_919) );
INVx1_ASAP7_75t_L g518 ( .A(n_194), .Y(n_518) );
INVx1_ASAP7_75t_L g927 ( .A(n_195), .Y(n_927) );
AOI22xp5_ASAP7_75t_L g1410 ( .A1(n_196), .A2(n_266), .B1(n_1411), .B2(n_1414), .Y(n_1410) );
INVxp33_ASAP7_75t_SL g1089 ( .A(n_197), .Y(n_1089) );
INVxp33_ASAP7_75t_SL g1221 ( .A(n_198), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_199), .A2(n_271), .B1(n_688), .B2(n_689), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_199), .A2(n_271), .B1(n_614), .B2(n_618), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_201), .A2(n_276), .B1(n_610), .B2(n_931), .Y(n_971) );
INVx1_ASAP7_75t_L g983 ( .A(n_201), .Y(n_983) );
INVx1_ASAP7_75t_L g1660 ( .A(n_202), .Y(n_1660) );
INVxp33_ASAP7_75t_SL g376 ( .A(n_203), .Y(n_376) );
INVx1_ASAP7_75t_L g1223 ( .A(n_204), .Y(n_1223) );
INVx1_ASAP7_75t_L g1345 ( .A(n_205), .Y(n_1345) );
INVx1_ASAP7_75t_L g599 ( .A(n_207), .Y(n_599) );
CKINVDCx16_ASAP7_75t_R g1424 ( .A(n_210), .Y(n_1424) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_212), .A2(n_241), .B1(n_640), .B2(n_643), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_212), .A2(n_241), .B1(n_500), .B2(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g937 ( .A(n_215), .Y(n_937) );
CKINVDCx5p33_ASAP7_75t_R g1018 ( .A(n_217), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_218), .A2(n_251), .B1(n_672), .B2(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g713 ( .A(n_218), .Y(n_713) );
INVxp67_ASAP7_75t_SL g867 ( .A(n_219), .Y(n_867) );
INVx1_ASAP7_75t_L g527 ( .A(n_220), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g809 ( .A(n_223), .Y(n_809) );
INVx1_ASAP7_75t_L g1661 ( .A(n_225), .Y(n_1661) );
OAI22xp5_ASAP7_75t_L g1682 ( .A1(n_225), .A2(n_237), .B1(n_416), .B2(n_618), .Y(n_1682) );
INVxp33_ASAP7_75t_L g1278 ( .A(n_226), .Y(n_1278) );
CKINVDCx5p33_ASAP7_75t_R g979 ( .A(n_227), .Y(n_979) );
INVxp33_ASAP7_75t_L g1252 ( .A(n_228), .Y(n_1252) );
BUFx3_ASAP7_75t_L g375 ( .A(n_229), .Y(n_375) );
INVx1_ASAP7_75t_L g381 ( .A(n_229), .Y(n_381) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_230), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_230), .A2(n_240), .B1(n_545), .B2(n_548), .Y(n_544) );
INVx1_ASAP7_75t_L g953 ( .A(n_231), .Y(n_953) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_232), .A2(n_300), .B1(n_344), .B2(n_416), .Y(n_631) );
INVx1_ASAP7_75t_L g1178 ( .A(n_233), .Y(n_1178) );
INVx1_ASAP7_75t_L g1031 ( .A(n_235), .Y(n_1031) );
OAI22xp5_ASAP7_75t_L g1070 ( .A1(n_235), .A2(n_289), .B1(n_344), .B2(n_416), .Y(n_1070) );
INVx1_ASAP7_75t_L g1183 ( .A(n_236), .Y(n_1183) );
OAI22xp5_ASAP7_75t_L g1675 ( .A1(n_237), .A2(n_244), .B1(n_610), .B2(n_931), .Y(n_1675) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_238), .Y(n_343) );
INVx1_ASAP7_75t_L g483 ( .A(n_238), .Y(n_483) );
AND2x2_ASAP7_75t_L g789 ( .A(n_238), .B(n_419), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_238), .B(n_305), .Y(n_803) );
INVx1_ASAP7_75t_L g784 ( .A(n_239), .Y(n_784) );
OAI221xp5_ASAP7_75t_L g796 ( .A1(n_239), .A2(n_327), .B1(n_797), .B2(n_804), .C(n_806), .Y(n_796) );
INVxp33_ASAP7_75t_SL g516 ( .A(n_240), .Y(n_516) );
INVx1_ASAP7_75t_L g1544 ( .A(n_242), .Y(n_1544) );
CKINVDCx5p33_ASAP7_75t_R g1373 ( .A(n_243), .Y(n_1373) );
INVx1_ASAP7_75t_L g1669 ( .A(n_244), .Y(n_1669) );
INVx1_ASAP7_75t_L g1429 ( .A(n_246), .Y(n_1429) );
XNOR2xp5_ASAP7_75t_L g1641 ( .A(n_246), .B(n_1642), .Y(n_1641) );
AOI22xp5_ASAP7_75t_L g1692 ( .A1(n_246), .A2(n_1693), .B1(n_1698), .B2(n_1701), .Y(n_1692) );
INVx2_ASAP7_75t_L g368 ( .A(n_248), .Y(n_368) );
INVxp67_ASAP7_75t_SL g790 ( .A(n_249), .Y(n_790) );
INVx1_ASAP7_75t_L g1259 ( .A(n_250), .Y(n_1259) );
INVxp67_ASAP7_75t_SL g712 ( .A(n_251), .Y(n_712) );
INVx1_ASAP7_75t_L g1542 ( .A(n_252), .Y(n_1542) );
INVxp33_ASAP7_75t_SL g721 ( .A(n_253), .Y(n_721) );
AOI22xp33_ASAP7_75t_SL g767 ( .A1(n_253), .A2(n_257), .B1(n_768), .B2(n_769), .Y(n_767) );
INVx1_ASAP7_75t_L g1680 ( .A(n_254), .Y(n_1680) );
INVxp67_ASAP7_75t_L g444 ( .A(n_255), .Y(n_444) );
CKINVDCx16_ASAP7_75t_R g1426 ( .A(n_256), .Y(n_1426) );
INVxp33_ASAP7_75t_SL g722 ( .A(n_257), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g1376 ( .A1(n_258), .A2(n_295), .B1(n_416), .B2(n_618), .Y(n_1376) );
INVx1_ASAP7_75t_L g941 ( .A(n_259), .Y(n_941) );
INVx1_ASAP7_75t_L g1434 ( .A(n_260), .Y(n_1434) );
INVxp33_ASAP7_75t_SL g734 ( .A(n_261), .Y(n_734) );
INVx1_ASAP7_75t_L g383 ( .A(n_262), .Y(n_383) );
INVx1_ASAP7_75t_L g1351 ( .A(n_263), .Y(n_1351) );
INVx1_ASAP7_75t_L g1279 ( .A(n_264), .Y(n_1279) );
INVx1_ASAP7_75t_L g1365 ( .A(n_267), .Y(n_1365) );
OAI211xp5_ASAP7_75t_SL g1377 ( .A1(n_267), .A2(n_620), .B(n_624), .C(n_1378), .Y(n_1377) );
INVxp67_ASAP7_75t_SL g780 ( .A(n_268), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g1267 ( .A1(n_269), .A2(n_303), .B1(n_1268), .B2(n_1269), .Y(n_1267) );
OAI22xp5_ASAP7_75t_L g1276 ( .A1(n_269), .A2(n_303), .B1(n_432), .B2(n_435), .Y(n_1276) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_270), .Y(n_421) );
INVxp33_ASAP7_75t_L g1118 ( .A(n_272), .Y(n_1118) );
INVx1_ASAP7_75t_L g1229 ( .A(n_273), .Y(n_1229) );
INVx1_ASAP7_75t_L g1319 ( .A(n_274), .Y(n_1319) );
AOI22xp33_ASAP7_75t_L g1334 ( .A1(n_274), .A2(n_308), .B1(n_396), .B2(n_663), .Y(n_1334) );
INVxp67_ASAP7_75t_SL g1141 ( .A(n_275), .Y(n_1141) );
INVxp67_ASAP7_75t_SL g575 ( .A(n_277), .Y(n_575) );
INVx1_ASAP7_75t_L g1311 ( .A(n_278), .Y(n_1311) );
INVx1_ASAP7_75t_L g859 ( .A(n_280), .Y(n_859) );
INVx1_ASAP7_75t_L g726 ( .A(n_282), .Y(n_726) );
OAI22xp33_ASAP7_75t_L g604 ( .A1(n_283), .A2(n_300), .B1(n_605), .B2(n_610), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_283), .A2(n_311), .B1(n_651), .B2(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g1651 ( .A(n_285), .Y(n_1651) );
INVxp67_ASAP7_75t_SL g878 ( .A(n_286), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_286), .A2(n_307), .B1(n_896), .B2(n_897), .Y(n_895) );
INVxp33_ASAP7_75t_SL g1099 ( .A(n_287), .Y(n_1099) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_288), .Y(n_337) );
AND3x2_ASAP7_75t_L g1393 ( .A(n_288), .B(n_335), .C(n_1394), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1400 ( .A(n_288), .B(n_335), .Y(n_1400) );
OAI22xp5_ASAP7_75t_L g1079 ( .A1(n_289), .A2(n_316), .B1(n_610), .B2(n_931), .Y(n_1079) );
INVx2_ASAP7_75t_L g348 ( .A(n_290), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g1694 ( .A1(n_291), .A2(n_1695), .B1(n_1696), .B2(n_1697), .Y(n_1694) );
CKINVDCx5p33_ASAP7_75t_R g1695 ( .A(n_291), .Y(n_1695) );
AOI21xp33_ASAP7_75t_L g807 ( .A1(n_294), .A2(n_466), .B(n_808), .Y(n_807) );
INVxp67_ASAP7_75t_SL g836 ( .A(n_294), .Y(n_836) );
INVx1_ASAP7_75t_L g822 ( .A(n_297), .Y(n_822) );
INVx1_ASAP7_75t_L g1184 ( .A(n_298), .Y(n_1184) );
INVx1_ASAP7_75t_L g730 ( .A(n_299), .Y(n_730) );
CKINVDCx5p33_ASAP7_75t_R g974 ( .A(n_301), .Y(n_974) );
INVxp67_ASAP7_75t_SL g1347 ( .A(n_302), .Y(n_1347) );
INVx1_ASAP7_75t_L g1344 ( .A(n_304), .Y(n_1344) );
INVx1_ASAP7_75t_L g350 ( .A(n_305), .Y(n_350) );
INVx2_ASAP7_75t_L g419 ( .A(n_305), .Y(n_419) );
XNOR2xp5_ASAP7_75t_L g1301 ( .A(n_306), .B(n_1302), .Y(n_1301) );
INVxp67_ASAP7_75t_SL g880 ( .A(n_307), .Y(n_880) );
INVx1_ASAP7_75t_L g1316 ( .A(n_308), .Y(n_1316) );
INVx1_ASAP7_75t_L g820 ( .A(n_310), .Y(n_820) );
INVx1_ASAP7_75t_L g596 ( .A(n_311), .Y(n_596) );
CKINVDCx5p33_ASAP7_75t_R g975 ( .A(n_314), .Y(n_975) );
INVx1_ASAP7_75t_L g1435 ( .A(n_315), .Y(n_1435) );
INVx1_ASAP7_75t_L g1065 ( .A(n_316), .Y(n_1065) );
INVxp33_ASAP7_75t_SL g579 ( .A(n_317), .Y(n_579) );
INVxp67_ASAP7_75t_SL g1115 ( .A(n_319), .Y(n_1115) );
INVx1_ASAP7_75t_L g1309 ( .A(n_321), .Y(n_1309) );
INVx1_ASAP7_75t_L g1212 ( .A(n_323), .Y(n_1212) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_324), .A2(n_326), .B1(n_1242), .B2(n_1243), .Y(n_1241) );
INVxp33_ASAP7_75t_L g1249 ( .A(n_324), .Y(n_1249) );
INVx1_ASAP7_75t_L g779 ( .A(n_325), .Y(n_779) );
INVxp67_ASAP7_75t_SL g1250 ( .A(n_326), .Y(n_1250) );
INVx1_ASAP7_75t_L g783 ( .A(n_327), .Y(n_783) );
INVxp67_ASAP7_75t_SL g399 ( .A(n_328), .Y(n_399) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_351), .B(n_1381), .Y(n_329) );
BUFx12f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_333), .B(n_338), .Y(n_332) );
AND2x4_ASAP7_75t_L g1691 ( .A(n_333), .B(n_339), .Y(n_1691) );
NOR2xp33_ASAP7_75t_SL g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx1_ASAP7_75t_SL g1700 ( .A(n_334), .Y(n_1700) );
NAND2xp5_ASAP7_75t_L g1704 ( .A(n_334), .B(n_336), .Y(n_1704) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g1699 ( .A(n_336), .B(n_1700), .Y(n_1699) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_344), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x6_ASAP7_75t_L g450 ( .A(n_341), .B(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g1122 ( .A(n_341), .B(n_451), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g469 ( .A(n_342), .B(n_350), .Y(n_469) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g1043 ( .A(n_343), .B(n_418), .Y(n_1043) );
INVx8_ASAP7_75t_L g414 ( .A(n_344), .Y(n_414) );
OR2x6_ASAP7_75t_L g344 ( .A(n_345), .B(n_349), .Y(n_344) );
OR2x6_ASAP7_75t_L g416 ( .A(n_345), .B(n_417), .Y(n_416) );
OAI21xp33_ASAP7_75t_L g808 ( .A1(n_345), .A2(n_469), .B(n_809), .Y(n_808) );
HB1xp67_ASAP7_75t_L g936 ( .A(n_345), .Y(n_936) );
INVx2_ASAP7_75t_SL g943 ( .A(n_345), .Y(n_943) );
BUFx6f_ASAP7_75t_L g1001 ( .A(n_345), .Y(n_1001) );
INVx2_ASAP7_75t_SL g1054 ( .A(n_345), .Y(n_1054) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g425 ( .A(n_347), .Y(n_425) );
INVx1_ASAP7_75t_L g437 ( .A(n_347), .Y(n_437) );
INVx2_ASAP7_75t_L g441 ( .A(n_347), .Y(n_441) );
AND2x4_ASAP7_75t_L g448 ( .A(n_347), .B(n_426), .Y(n_448) );
AND2x2_ASAP7_75t_L g464 ( .A(n_347), .B(n_348), .Y(n_464) );
INVx2_ASAP7_75t_L g426 ( .A(n_348), .Y(n_426) );
INVx1_ASAP7_75t_L g434 ( .A(n_348), .Y(n_434) );
INVx1_ASAP7_75t_L g443 ( .A(n_348), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_348), .B(n_441), .Y(n_617) );
INVx1_ASAP7_75t_L g623 ( .A(n_348), .Y(n_623) );
AND2x4_ASAP7_75t_L g433 ( .A(n_349), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g435 ( .A(n_350), .B(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g577 ( .A(n_350), .B(n_436), .Y(n_577) );
XNOR2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_585), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_509), .B1(n_510), .B2(n_584), .Y(n_352) );
INVx1_ASAP7_75t_L g584 ( .A(n_353), .Y(n_584) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AO211x2_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_362), .B(n_411), .C(n_452), .Y(n_356) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_357), .Y(n_529) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_357), .A2(n_632), .B1(n_719), .B2(n_731), .C(n_739), .Y(n_718) );
INVx1_ASAP7_75t_L g885 ( .A(n_357), .Y(n_885) );
OAI31xp33_ASAP7_75t_SL g1077 ( .A1(n_357), .A2(n_1078), .A3(n_1079), .B(n_1080), .Y(n_1077) );
OAI21xp5_ASAP7_75t_L g1132 ( .A1(n_357), .A2(n_1133), .B(n_1142), .Y(n_1132) );
AND2x4_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
AND2x4_ASAP7_75t_L g611 ( .A(n_358), .B(n_360), .Y(n_611) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g497 ( .A(n_359), .B(n_368), .Y(n_497) );
AND2x4_ASAP7_75t_L g507 ( .A(n_359), .B(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g468 ( .A(n_361), .Y(n_468) );
OR2x6_ASAP7_75t_L g1042 ( .A(n_361), .B(n_1043), .Y(n_1042) );
NAND4xp25_ASAP7_75t_SL g362 ( .A(n_363), .B(n_382), .C(n_392), .D(n_407), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B1(n_376), .B2(n_377), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_365), .A2(n_377), .B1(n_733), .B2(n_734), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_365), .A2(n_377), .B1(n_877), .B2(n_878), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_365), .A2(n_377), .B1(n_1089), .B2(n_1090), .Y(n_1088) );
AOI22xp5_ASAP7_75t_L g1179 ( .A1(n_365), .A2(n_377), .B1(n_1180), .B2(n_1181), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_365), .A2(n_377), .B1(n_1220), .B2(n_1221), .Y(n_1219) );
AOI22xp5_ASAP7_75t_SL g1262 ( .A1(n_365), .A2(n_384), .B1(n_1263), .B2(n_1264), .Y(n_1262) );
AND2x4_ASAP7_75t_L g365 ( .A(n_366), .B(n_369), .Y(n_365) );
AND2x6_ASAP7_75t_L g388 ( .A(n_366), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g515 ( .A(n_366), .B(n_369), .Y(n_515) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g709 ( .A(n_367), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g379 ( .A(n_368), .Y(n_379) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_368), .Y(n_386) );
INVx2_ASAP7_75t_L g508 ( .A(n_368), .Y(n_508) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_370), .Y(n_487) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_370), .Y(n_562) );
INVx2_ASAP7_75t_L g566 ( .A(n_370), .Y(n_566) );
INVx1_ASAP7_75t_L g691 ( .A(n_370), .Y(n_691) );
INVx2_ASAP7_75t_SL g758 ( .A(n_370), .Y(n_758) );
INVx2_ASAP7_75t_L g766 ( .A(n_370), .Y(n_766) );
INVx1_ASAP7_75t_L g1294 ( .A(n_370), .Y(n_1294) );
INVx6_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g384 ( .A(n_371), .B(n_385), .Y(n_384) );
BUFx2_ASAP7_75t_L g500 ( .A(n_371), .Y(n_500) );
INVx2_ASAP7_75t_L g664 ( .A(n_371), .Y(n_664) );
AND2x4_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx1_ASAP7_75t_L g406 ( .A(n_372), .Y(n_406) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g380 ( .A(n_373), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g398 ( .A(n_373), .B(n_375), .Y(n_398) );
INVx1_ASAP7_75t_L g403 ( .A(n_374), .Y(n_403) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g390 ( .A(n_375), .B(n_391), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_377), .A2(n_514), .B1(n_515), .B2(n_516), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_377), .A2(n_388), .B1(n_602), .B2(n_603), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_377), .A2(n_388), .B1(n_712), .B2(n_713), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_377), .A2(n_515), .B1(n_776), .B2(n_777), .Y(n_775) );
CKINVDCx6p67_ASAP7_75t_R g930 ( .A(n_377), .Y(n_930) );
AOI22xp5_ASAP7_75t_L g1270 ( .A1(n_377), .A2(n_388), .B1(n_1271), .B2(n_1272), .Y(n_1270) );
AOI22xp5_ASAP7_75t_L g1307 ( .A1(n_377), .A2(n_388), .B1(n_1308), .B2(n_1309), .Y(n_1307) );
AND2x6_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx1_ASAP7_75t_L g409 ( .A(n_378), .Y(n_409) );
INVx1_ASAP7_75t_L g606 ( .A(n_378), .Y(n_606) );
AND2x2_ASAP7_75t_L g925 ( .A(n_378), .B(n_523), .Y(n_925) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x6_ASAP7_75t_L g405 ( .A(n_379), .B(n_406), .Y(n_405) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_380), .Y(n_491) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_380), .Y(n_559) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_380), .Y(n_688) );
BUFx2_ASAP7_75t_L g760 ( .A(n_380), .Y(n_760) );
BUFx6f_ASAP7_75t_L g906 ( .A(n_380), .Y(n_906) );
BUFx3_ASAP7_75t_L g915 ( .A(n_380), .Y(n_915) );
INVx2_ASAP7_75t_SL g1198 ( .A(n_380), .Y(n_1198) );
HB1xp67_ASAP7_75t_L g1238 ( .A(n_380), .Y(n_1238) );
INVx1_ASAP7_75t_L g609 ( .A(n_381), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B1(n_387), .B2(n_388), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_383), .A2(n_413), .B1(n_414), .B2(n_415), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_384), .A2(n_388), .B1(n_518), .B2(n_519), .Y(n_517) );
INVx4_ASAP7_75t_L g610 ( .A(n_384), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_384), .A2(n_388), .B1(n_730), .B2(n_736), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_384), .A2(n_388), .B1(n_779), .B2(n_780), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_384), .A2(n_388), .B1(n_863), .B2(n_880), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_384), .A2(n_388), .B1(n_1098), .B2(n_1099), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_384), .A2(n_388), .B1(n_1140), .B2(n_1141), .Y(n_1139) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_384), .A2(n_388), .B1(n_1177), .B2(n_1178), .Y(n_1176) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_384), .A2(n_388), .B1(n_1223), .B2(n_1224), .Y(n_1222) );
AOI22xp5_ASAP7_75t_SL g1304 ( .A1(n_384), .A2(n_515), .B1(n_1305), .B2(n_1306), .Y(n_1304) );
AND2x2_ASAP7_75t_SL g400 ( .A(n_385), .B(n_401), .Y(n_400) );
AND2x4_ASAP7_75t_L g526 ( .A(n_385), .B(n_401), .Y(n_526) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx4_ASAP7_75t_L g931 ( .A(n_388), .Y(n_931) );
INVx1_ASAP7_75t_L g504 ( .A(n_389), .Y(n_504) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_389), .Y(n_689) );
INVx1_ASAP7_75t_L g852 ( .A(n_389), .Y(n_852) );
BUFx6f_ASAP7_75t_L g916 ( .A(n_389), .Y(n_916) );
INVx2_ASAP7_75t_L g1028 ( .A(n_389), .Y(n_1028) );
INVx1_ASAP7_75t_L g1203 ( .A(n_389), .Y(n_1203) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_390), .Y(n_493) );
INVx1_ASAP7_75t_L g685 ( .A(n_390), .Y(n_685) );
INVx1_ASAP7_75t_L g762 ( .A(n_390), .Y(n_762) );
INVx2_ASAP7_75t_L g841 ( .A(n_390), .Y(n_841) );
INVx1_ASAP7_75t_L g608 ( .A(n_391), .Y(n_608) );
AOI222xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B1(n_399), .B2(n_400), .C1(n_404), .C2(n_405), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx3_ASAP7_75t_L g563 ( .A(n_397), .Y(n_563) );
BUFx4f_ASAP7_75t_L g567 ( .A(n_397), .Y(n_567) );
INVx1_ASAP7_75t_L g598 ( .A(n_397), .Y(n_598) );
INVx2_ASAP7_75t_SL g656 ( .A(n_397), .Y(n_656) );
INVx1_ASAP7_75t_L g1094 ( .A(n_397), .Y(n_1094) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_398), .Y(n_410) );
AOI222xp33_ASAP7_75t_L g595 ( .A1(n_400), .A2(n_405), .B1(n_596), .B2(n_597), .C1(n_599), .C2(n_600), .Y(n_595) );
AOI222xp33_ASAP7_75t_L g737 ( .A1(n_400), .A2(n_405), .B1(n_692), .B2(n_725), .C1(n_726), .C2(n_738), .Y(n_737) );
AOI222xp33_ASAP7_75t_L g781 ( .A1(n_400), .A2(n_405), .B1(n_563), .B2(n_782), .C1(n_783), .C2(n_784), .Y(n_781) );
AOI222xp33_ASAP7_75t_L g1091 ( .A1(n_400), .A2(n_405), .B1(n_1092), .B2(n_1093), .C1(n_1095), .C2(n_1096), .Y(n_1091) );
AOI222xp33_ASAP7_75t_L g1182 ( .A1(n_400), .A2(n_405), .B1(n_563), .B2(n_1183), .C1(n_1184), .C2(n_1185), .Y(n_1182) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g710 ( .A(n_402), .Y(n_710) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI222xp33_ASAP7_75t_L g520 ( .A1(n_405), .A2(n_521), .B1(n_522), .B2(n_524), .C1(n_525), .C2(n_527), .Y(n_520) );
AOI222xp33_ASAP7_75t_L g706 ( .A1(n_405), .A2(n_701), .B1(n_702), .B2(n_707), .C1(n_708), .C2(n_709), .Y(n_706) );
AOI222xp33_ASAP7_75t_L g881 ( .A1(n_405), .A2(n_525), .B1(n_866), .B2(n_868), .C1(n_882), .C2(n_883), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_405), .A2(n_526), .B1(n_927), .B2(n_928), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_405), .A2(n_526), .B1(n_974), .B2(n_975), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_405), .A2(n_526), .B1(n_1074), .B2(n_1075), .Y(n_1083) );
AOI22xp5_ASAP7_75t_L g1136 ( .A1(n_405), .A2(n_709), .B1(n_1137), .B2(n_1138), .Y(n_1136) );
AOI222xp33_ASAP7_75t_L g1225 ( .A1(n_405), .A2(n_525), .B1(n_1226), .B2(n_1227), .C1(n_1228), .C2(n_1229), .Y(n_1225) );
INVx3_ASAP7_75t_L g1269 ( .A(n_405), .Y(n_1269) );
AOI222xp33_ASAP7_75t_L g1370 ( .A1(n_405), .A2(n_709), .B1(n_1357), .B2(n_1371), .C1(n_1372), .C2(n_1373), .Y(n_1370) );
AOI222xp33_ASAP7_75t_L g1677 ( .A1(n_405), .A2(n_709), .B1(n_1672), .B2(n_1678), .C1(n_1679), .C2(n_1680), .Y(n_1677) );
NAND3xp33_ASAP7_75t_SL g594 ( .A(n_407), .B(n_595), .C(n_601), .Y(n_594) );
NAND3xp33_ASAP7_75t_SL g705 ( .A(n_407), .B(n_706), .C(n_711), .Y(n_705) );
NAND4xp25_ASAP7_75t_SL g731 ( .A(n_407), .B(n_732), .C(n_735), .D(n_737), .Y(n_731) );
NAND4xp25_ASAP7_75t_L g1087 ( .A(n_407), .B(n_1088), .C(n_1091), .D(n_1097), .Y(n_1087) );
NAND2xp5_ASAP7_75t_SL g1369 ( .A(n_407), .B(n_1370), .Y(n_1369) );
NAND2xp5_ASAP7_75t_SL g1676 ( .A(n_407), .B(n_1677), .Y(n_1676) );
CKINVDCx8_ASAP7_75t_R g407 ( .A(n_408), .Y(n_407) );
INVx5_ASAP7_75t_L g528 ( .A(n_408), .Y(n_528) );
NOR2xp33_ASAP7_75t_SL g1134 ( .A(n_408), .B(n_1135), .Y(n_1134) );
AND2x4_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_410), .Y(n_489) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_410), .Y(n_523) );
INVx2_ASAP7_75t_L g693 ( .A(n_410), .Y(n_693) );
INVx1_ASAP7_75t_L g1038 ( .A(n_410), .Y(n_1038) );
AOI31xp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_420), .A3(n_438), .B(n_450), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g581 ( .A1(n_414), .A2(n_518), .B1(n_582), .B2(n_583), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_414), .A2(n_583), .B1(n_729), .B2(n_730), .Y(n_728) );
AOI22xp33_ASAP7_75t_SL g871 ( .A1(n_414), .A2(n_872), .B1(n_873), .B2(n_874), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_414), .A2(n_583), .B1(n_952), .B2(n_961), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_414), .A2(n_583), .B1(n_982), .B2(n_983), .Y(n_981) );
AOI22xp33_ASAP7_75t_SL g1120 ( .A1(n_414), .A2(n_415), .B1(n_1098), .B2(n_1121), .Y(n_1120) );
AOI22xp33_ASAP7_75t_SL g1211 ( .A1(n_414), .A2(n_583), .B1(n_1177), .B2(n_1212), .Y(n_1211) );
AOI22xp33_ASAP7_75t_L g1251 ( .A1(n_414), .A2(n_415), .B1(n_1223), .B2(n_1252), .Y(n_1251) );
AOI22xp33_ASAP7_75t_SL g1277 ( .A1(n_414), .A2(n_439), .B1(n_1278), .B2(n_1279), .Y(n_1277) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_414), .A2(n_439), .B1(n_1319), .B2(n_1320), .Y(n_1318) );
AOI22xp33_ASAP7_75t_SL g1280 ( .A1(n_415), .A2(n_445), .B1(n_1264), .B2(n_1281), .Y(n_1280) );
AOI22xp33_ASAP7_75t_L g1321 ( .A1(n_415), .A2(n_445), .B1(n_1306), .B2(n_1322), .Y(n_1321) );
INVx5_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx4_ASAP7_75t_L g583 ( .A(n_416), .Y(n_583) );
AND2x4_ASAP7_75t_L g439 ( .A(n_417), .B(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g445 ( .A(n_417), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g615 ( .A(n_417), .Y(n_615) );
AND2x4_ASAP7_75t_L g873 ( .A(n_417), .B(n_446), .Y(n_873) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g430 ( .A(n_419), .Y(n_430) );
AOI211xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B(n_427), .C(n_431), .Y(n_420) );
AOI211xp5_ASAP7_75t_SL g574 ( .A1(n_422), .A2(n_427), .B(n_575), .C(n_576), .Y(n_574) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g427 ( .A(n_424), .B(n_428), .Y(n_427) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_424), .Y(n_466) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_424), .Y(n_538) );
BUFx2_ASAP7_75t_L g552 ( .A(n_424), .Y(n_552) );
BUFx3_ASAP7_75t_L g644 ( .A(n_424), .Y(n_644) );
BUFx3_ASAP7_75t_L g959 ( .A(n_424), .Y(n_959) );
AND2x4_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
CKINVDCx11_ASAP7_75t_R g624 ( .A(n_427), .Y(n_624) );
AOI211xp5_ASAP7_75t_L g1114 ( .A1(n_427), .A2(n_744), .B(n_1115), .C(n_1116), .Y(n_1114) );
NOR3xp33_ASAP7_75t_L g1144 ( .A(n_427), .B(n_1145), .C(n_1146), .Y(n_1144) );
AOI211xp5_ASAP7_75t_L g1205 ( .A1(n_427), .A2(n_744), .B(n_1206), .C(n_1207), .Y(n_1205) );
AOI211xp5_ASAP7_75t_L g1245 ( .A1(n_427), .A2(n_643), .B(n_1246), .C(n_1247), .Y(n_1245) );
AOI211xp5_ASAP7_75t_L g1274 ( .A1(n_427), .A2(n_958), .B(n_1275), .C(n_1276), .Y(n_1274) );
AOI211xp5_ASAP7_75t_L g1315 ( .A1(n_427), .A2(n_476), .B(n_1316), .C(n_1317), .Y(n_1315) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g630 ( .A(n_429), .Y(n_630) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2x1p5_ASAP7_75t_L g482 ( .A(n_430), .B(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g627 ( .A(n_433), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_433), .A2(n_628), .B1(n_701), .B2(n_702), .Y(n_700) );
AOI222xp33_ASAP7_75t_L g723 ( .A1(n_433), .A2(n_466), .B1(n_724), .B2(n_725), .C1(n_726), .C2(n_727), .Y(n_723) );
INVx2_ASAP7_75t_L g870 ( .A(n_433), .Y(n_870) );
AOI222xp33_ASAP7_75t_L g957 ( .A1(n_433), .A2(n_628), .B1(n_927), .B2(n_928), .C1(n_953), .C2(n_958), .Y(n_957) );
AOI222xp33_ASAP7_75t_SL g978 ( .A1(n_433), .A2(n_727), .B1(n_974), .B2(n_975), .C1(n_979), .C2(n_980), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_433), .A2(n_628), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
AOI22xp5_ASAP7_75t_L g1378 ( .A1(n_433), .A2(n_628), .B1(n_1372), .B2(n_1373), .Y(n_1378) );
AOI22xp33_ASAP7_75t_L g1684 ( .A1(n_433), .A2(n_628), .B1(n_1679), .B2(n_1680), .Y(n_1684) );
INVx1_ASAP7_75t_L g799 ( .A(n_434), .Y(n_799) );
INVx1_ASAP7_75t_L g629 ( .A(n_436), .Y(n_629) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g622 ( .A(n_437), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_437), .B(n_623), .Y(n_995) );
AOI22xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_444), .B1(n_445), .B2(n_449), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_439), .A2(n_445), .B1(n_579), .B2(n_580), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_439), .A2(n_445), .B1(n_721), .B2(n_722), .Y(n_720) );
AOI22xp33_ASAP7_75t_SL g862 ( .A1(n_439), .A2(n_583), .B1(n_863), .B2(n_864), .Y(n_862) );
AOI22xp33_ASAP7_75t_SL g1117 ( .A1(n_439), .A2(n_873), .B1(n_1118), .B2(n_1119), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_439), .A2(n_873), .B1(n_1148), .B2(n_1149), .Y(n_1147) );
AOI22xp33_ASAP7_75t_SL g1208 ( .A1(n_439), .A2(n_873), .B1(n_1209), .B2(n_1210), .Y(n_1208) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_439), .A2(n_445), .B1(n_1249), .B2(n_1250), .Y(n_1248) );
INVx1_ASAP7_75t_L g456 ( .A(n_440), .Y(n_456) );
BUFx2_ASAP7_75t_L g540 ( .A(n_440), .Y(n_540) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_440), .Y(n_547) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_440), .Y(n_647) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_440), .Y(n_672) );
AND2x2_ASAP7_75t_L g788 ( .A(n_440), .B(n_789), .Y(n_788) );
BUFx2_ASAP7_75t_L g896 ( .A(n_440), .Y(n_896) );
INVx1_ASAP7_75t_L g1158 ( .A(n_440), .Y(n_1158) );
AND2x4_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g805 ( .A(n_441), .Y(n_805) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx5_ASAP7_75t_SL g618 ( .A(n_445), .Y(n_618) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g1290 ( .A(n_447), .Y(n_1290) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g459 ( .A(n_448), .Y(n_459) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_448), .Y(n_543) );
INVx1_ASAP7_75t_L g750 ( .A(n_448), .Y(n_750) );
AOI31xp33_ASAP7_75t_L g573 ( .A1(n_450), .A2(n_574), .A3(n_578), .B(n_581), .Y(n_573) );
CKINVDCx16_ASAP7_75t_R g632 ( .A(n_450), .Y(n_632) );
AOI31xp33_ASAP7_75t_L g1204 ( .A1(n_450), .A2(n_1205), .A3(n_1208), .B(n_1211), .Y(n_1204) );
AOI31xp33_ASAP7_75t_L g1244 ( .A1(n_450), .A2(n_1245), .A3(n_1248), .B(n_1251), .Y(n_1244) );
AND2x4_ASAP7_75t_L g506 ( .A(n_451), .B(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g666 ( .A(n_451), .B(n_507), .Y(n_666) );
NAND4xp25_ASAP7_75t_L g452 ( .A(n_453), .B(n_470), .C(n_484), .D(n_498), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_460), .C(n_467), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g636 ( .A(n_456), .Y(n_636) );
INVx1_ASAP7_75t_L g742 ( .A(n_456), .Y(n_742) );
BUFx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g890 ( .A(n_458), .Y(n_890) );
INVx2_ASAP7_75t_L g1352 ( .A(n_458), .Y(n_1352) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx3_ASAP7_75t_L g474 ( .A(n_459), .Y(n_474) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_459), .Y(n_649) );
BUFx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g1153 ( .A(n_462), .Y(n_1153) );
INVx2_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g535 ( .A(n_463), .Y(n_535) );
INVx2_ASAP7_75t_SL g753 ( .A(n_463), .Y(n_753) );
INVx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_464), .Y(n_642) );
BUFx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_SL g477 ( .A(n_466), .Y(n_477) );
NAND3xp33_ASAP7_75t_L g634 ( .A(n_467), .B(n_635), .C(n_639), .Y(n_634) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_467), .B(n_671), .C(n_674), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g740 ( .A(n_467), .B(n_741), .C(n_743), .Y(n_740) );
INVx2_ASAP7_75t_L g893 ( .A(n_467), .Y(n_893) );
BUFx3_ASAP7_75t_L g938 ( .A(n_467), .Y(n_938) );
AOI33xp33_ASAP7_75t_L g1107 ( .A1(n_467), .A2(n_666), .A3(n_1108), .B1(n_1109), .B2(n_1111), .B3(n_1112), .Y(n_1107) );
NAND3xp33_ASAP7_75t_L g1187 ( .A(n_467), .B(n_1188), .C(n_1189), .Y(n_1187) );
NAND3xp33_ASAP7_75t_L g1283 ( .A(n_467), .B(n_1284), .C(n_1285), .Y(n_1283) );
NAND3xp33_ASAP7_75t_L g1324 ( .A(n_467), .B(n_1325), .C(n_1326), .Y(n_1324) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
OR2x6_ASAP7_75t_L g495 ( .A(n_468), .B(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_L g532 ( .A(n_468), .B(n_469), .Y(n_532) );
OR2x2_ASAP7_75t_L g659 ( .A(n_468), .B(n_660), .Y(n_659) );
BUFx2_ASAP7_75t_L g829 ( .A(n_468), .Y(n_829) );
OR2x2_ASAP7_75t_L g946 ( .A(n_468), .B(n_496), .Y(n_946) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_468), .B(n_816), .Y(n_1106) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_475), .C(n_478), .Y(n_470) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g638 ( .A(n_474), .Y(n_638) );
INVx1_ASAP7_75t_L g998 ( .A(n_474), .Y(n_998) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g652 ( .A(n_477), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g645 ( .A(n_478), .B(n_646), .C(n_650), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g745 ( .A(n_478), .B(n_746), .C(n_751), .Y(n_745) );
NAND3xp33_ASAP7_75t_L g894 ( .A(n_478), .B(n_895), .C(n_899), .Y(n_894) );
CKINVDCx8_ASAP7_75t_R g1068 ( .A(n_478), .Y(n_1068) );
INVx5_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx6_ASAP7_75t_L g553 ( .A(n_479), .Y(n_553) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g816 ( .A(n_482), .Y(n_816) );
NAND3xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_490), .C(n_494), .Y(n_484) );
INVx4_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g1169 ( .A(n_487), .Y(n_1169) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx4f_ASAP7_75t_L g502 ( .A(n_491), .Y(n_502) );
INVx1_ASAP7_75t_L g1647 ( .A(n_491), .Y(n_1647) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g571 ( .A(n_493), .Y(n_571) );
BUFx3_ASAP7_75t_L g769 ( .A(n_493), .Y(n_769) );
INVx1_ASAP7_75t_L g1649 ( .A(n_493), .Y(n_1649) );
INVx1_ASAP7_75t_L g842 ( .A(n_494), .Y(n_842) );
AOI33xp33_ASAP7_75t_L g1163 ( .A1(n_494), .A2(n_505), .A3(n_1164), .B1(n_1168), .B2(n_1170), .B3(n_1171), .Y(n_1163) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_495), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g908 ( .A(n_495), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g1016 ( .A1(n_495), .A2(n_911), .B1(n_1017), .B2(n_1029), .Y(n_1016) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g660 ( .A(n_497), .Y(n_660) );
NAND3xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .C(n_505), .Y(n_498) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g853 ( .A(n_505), .Y(n_853) );
BUFx4f_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx4f_ASAP7_75t_L g572 ( .A(n_506), .Y(n_572) );
INVx4_ASAP7_75t_L g911 ( .A(n_506), .Y(n_911) );
INVx2_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
AOI211xp5_ASAP7_75t_SL g511 ( .A1(n_512), .A2(n_529), .B(n_530), .C(n_573), .Y(n_511) );
NAND4xp25_ASAP7_75t_SL g512 ( .A(n_513), .B(n_517), .C(n_520), .D(n_528), .Y(n_512) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
HB1xp67_ASAP7_75t_L g1227 ( .A(n_523), .Y(n_1227) );
BUFx4f_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND4xp25_ASAP7_75t_L g774 ( .A(n_528), .B(n_775), .C(n_778), .D(n_781), .Y(n_774) );
NAND4xp25_ASAP7_75t_L g875 ( .A(n_528), .B(n_876), .C(n_879), .D(n_881), .Y(n_875) );
NAND4xp25_ASAP7_75t_L g1175 ( .A(n_528), .B(n_1176), .C(n_1179), .D(n_1182), .Y(n_1175) );
NAND4xp25_ASAP7_75t_SL g1218 ( .A(n_528), .B(n_1219), .C(n_1222), .D(n_1225), .Y(n_1218) );
NAND4xp25_ASAP7_75t_L g1261 ( .A(n_528), .B(n_1262), .C(n_1265), .D(n_1270), .Y(n_1261) );
NAND4xp25_ASAP7_75t_L g1303 ( .A(n_528), .B(n_1304), .C(n_1307), .D(n_1310), .Y(n_1303) );
AOI221x1_ASAP7_75t_L g773 ( .A1(n_529), .A2(n_774), .B1(n_785), .B2(n_827), .C(n_830), .Y(n_773) );
AOI211x1_ASAP7_75t_SL g1217 ( .A1(n_529), .A2(n_1218), .B(n_1230), .C(n_1244), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_554), .Y(n_530) );
AOI33xp33_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .A3(n_539), .B1(n_544), .B2(n_549), .B3(n_553), .Y(n_531) );
AOI33xp33_ASAP7_75t_L g1150 ( .A1(n_532), .A2(n_553), .A3(n_1151), .B1(n_1156), .B2(n_1161), .B3(n_1162), .Y(n_1150) );
BUFx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g900 ( .A(n_537), .Y(n_900) );
INVx2_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
BUFx6f_ASAP7_75t_L g744 ( .A(n_538), .Y(n_744) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
BUFx3_ASAP7_75t_L g548 ( .A(n_543), .Y(n_548) );
INVx2_ASAP7_75t_SL g898 ( .A(n_543), .Y(n_898) );
INVx2_ASAP7_75t_SL g988 ( .A(n_543), .Y(n_988) );
INVx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g980 ( .A(n_551), .Y(n_980) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_553), .B(n_677), .C(n_679), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g932 ( .A1(n_553), .A2(n_933), .B1(n_938), .B2(n_939), .C(n_945), .Y(n_932) );
AOI221xp5_ASAP7_75t_L g985 ( .A1(n_553), .A2(n_938), .B1(n_986), .B2(n_996), .C(n_1003), .Y(n_985) );
AOI33xp33_ASAP7_75t_L g1231 ( .A1(n_553), .A2(n_892), .A3(n_1232), .B1(n_1233), .B2(n_1234), .B3(n_1235), .Y(n_1231) );
AOI33xp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_556), .A3(n_560), .B1(n_564), .B2(n_568), .B3(n_572), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g754 ( .A(n_555), .B(n_755), .C(n_759), .Y(n_754) );
AOI33xp33_ASAP7_75t_L g1236 ( .A1(n_555), .A2(n_572), .A3(n_1237), .B1(n_1239), .B2(n_1240), .B3(n_1241), .Y(n_1236) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_SL g569 ( .A(n_558), .Y(n_569) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
BUFx3_ASAP7_75t_L g768 ( .A(n_559), .Y(n_768) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
BUFx2_ASAP7_75t_L g883 ( .A(n_567), .Y(n_883) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND3xp33_ASAP7_75t_L g763 ( .A(n_572), .B(n_764), .C(n_767), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B1(n_1336), .B2(n_1380), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
XNOR2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_963), .Y(n_587) );
XOR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_856), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_716), .B1(n_854), .B2(n_855), .Y(n_589) );
INVx2_ASAP7_75t_L g854 ( .A(n_590), .Y(n_854) );
XOR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_667), .Y(n_590) );
NAND3x1_ASAP7_75t_L g592 ( .A(n_593), .B(n_612), .C(n_633), .Y(n_592) );
OAI21xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_604), .B(n_611), .Y(n_593) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g708 ( .A(n_598), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_599), .A2(n_600), .B1(n_626), .B2(n_628), .Y(n_625) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g833 ( .A(n_607), .Y(n_833) );
INVx2_ASAP7_75t_L g846 ( .A(n_607), .Y(n_846) );
BUFx2_ASAP7_75t_L g1019 ( .A(n_607), .Y(n_1019) );
INVx1_ASAP7_75t_L g1653 ( .A(n_607), .Y(n_1653) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
AND2x2_ASAP7_75t_L g835 ( .A(n_608), .B(n_609), .Y(n_835) );
OAI21xp5_ASAP7_75t_SL g704 ( .A1(n_611), .A2(n_705), .B(n_714), .Y(n_704) );
OAI31xp33_ASAP7_75t_L g921 ( .A1(n_611), .A2(n_922), .A3(n_923), .B(n_929), .Y(n_921) );
OAI31xp33_ASAP7_75t_SL g969 ( .A1(n_611), .A2(n_970), .A3(n_971), .B(n_972), .Y(n_969) );
AOI211x1_ASAP7_75t_L g1086 ( .A1(n_611), .A2(n_1087), .B(n_1100), .C(n_1113), .Y(n_1086) );
AOI211xp5_ASAP7_75t_L g1174 ( .A1(n_611), .A2(n_1175), .B(n_1186), .C(n_1204), .Y(n_1174) );
AOI211xp5_ASAP7_75t_L g1260 ( .A1(n_611), .A2(n_1261), .B(n_1273), .C(n_1282), .Y(n_1260) );
AOI211xp5_ASAP7_75t_L g1302 ( .A1(n_611), .A2(n_1303), .B(n_1314), .C(n_1323), .Y(n_1302) );
OAI31xp33_ASAP7_75t_SL g1367 ( .A1(n_611), .A2(n_1368), .A3(n_1369), .B(n_1374), .Y(n_1367) );
OAI31xp33_ASAP7_75t_L g1673 ( .A1(n_611), .A2(n_1674), .A3(n_1675), .B(n_1676), .Y(n_1673) );
OAI31xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_619), .A3(n_631), .B(n_632), .Y(n_612) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
BUFx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g1048 ( .A(n_617), .Y(n_1048) );
INVx1_ASAP7_75t_L g1061 ( .A(n_617), .Y(n_1061) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g1066 ( .A(n_621), .Y(n_1066) );
BUFx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g699 ( .A(n_622), .Y(n_699) );
INVx3_ASAP7_75t_L g813 ( .A(n_622), .Y(n_813) );
INVx2_ASAP7_75t_L g1356 ( .A(n_622), .Y(n_1356) );
NAND4xp25_ASAP7_75t_L g719 ( .A(n_624), .B(n_720), .C(n_723), .D(n_728), .Y(n_719) );
NAND4xp25_ASAP7_75t_L g861 ( .A(n_624), .B(n_862), .C(n_865), .D(n_871), .Y(n_861) );
NAND3xp33_ASAP7_75t_L g956 ( .A(n_624), .B(n_957), .C(n_960), .Y(n_956) );
NAND3xp33_ASAP7_75t_SL g977 ( .A(n_624), .B(n_978), .C(n_981), .Y(n_977) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AOI222xp33_ASAP7_75t_L g865 ( .A1(n_628), .A2(n_744), .B1(n_866), .B2(n_867), .C1(n_868), .C2(n_869), .Y(n_865) );
AND2x4_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
AND2x4_ASAP7_75t_L g727 ( .A(n_629), .B(n_630), .Y(n_727) );
OAI31xp33_ASAP7_75t_SL g694 ( .A1(n_632), .A2(n_695), .A3(n_696), .B(n_703), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g860 ( .A1(n_632), .A2(n_861), .B1(n_875), .B2(n_884), .C(n_886), .Y(n_860) );
OAI21xp5_ASAP7_75t_L g955 ( .A1(n_632), .A2(n_956), .B(n_962), .Y(n_955) );
OAI21xp5_ASAP7_75t_L g976 ( .A1(n_632), .A2(n_977), .B(n_984), .Y(n_976) );
OAI31xp33_ASAP7_75t_SL g1069 ( .A1(n_632), .A2(n_1070), .A3(n_1071), .B(n_1076), .Y(n_1069) );
OAI31xp33_ASAP7_75t_SL g1375 ( .A1(n_632), .A2(n_1376), .A3(n_1377), .B(n_1379), .Y(n_1375) );
OAI31xp33_ASAP7_75t_SL g1681 ( .A1(n_632), .A2(n_1682), .A3(n_1683), .B(n_1685), .Y(n_1681) );
AND4x1_ASAP7_75t_L g633 ( .A(n_634), .B(n_645), .C(n_653), .D(n_661), .Y(n_633) );
INVx1_ASAP7_75t_L g1064 ( .A(n_637), .Y(n_1064) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g675 ( .A(n_641), .Y(n_675) );
INVx2_ASAP7_75t_L g1286 ( .A(n_641), .Y(n_1286) );
INVx3_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
BUFx2_ASAP7_75t_L g651 ( .A(n_642), .Y(n_651) );
AND2x4_ASAP7_75t_L g823 ( .A(n_642), .B(n_789), .Y(n_823) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x4_ASAP7_75t_L g821 ( .A(n_644), .B(n_792), .Y(n_821) );
INVx1_ASAP7_75t_L g1155 ( .A(n_644), .Y(n_1155) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g673 ( .A(n_649), .Y(n_673) );
INVx2_ASAP7_75t_L g678 ( .A(n_649), .Y(n_678) );
INVx2_ASAP7_75t_SL g1192 ( .A(n_649), .Y(n_1192) );
NAND3xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_657), .C(n_658), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g1167 ( .A(n_656), .Y(n_1167) );
INVx1_ASAP7_75t_L g1371 ( .A(n_656), .Y(n_1371) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_658), .B(n_681), .C(n_683), .Y(n_680) );
AOI33xp33_ASAP7_75t_L g1101 ( .A1(n_658), .A2(n_1102), .A3(n_1103), .B1(n_1104), .B2(n_1105), .B3(n_1106), .Y(n_1101) );
NAND3xp33_ASAP7_75t_L g1194 ( .A(n_658), .B(n_1195), .C(n_1196), .Y(n_1194) );
NAND3xp33_ASAP7_75t_L g1292 ( .A(n_658), .B(n_1293), .C(n_1295), .Y(n_1292) );
NAND3xp33_ASAP7_75t_L g1330 ( .A(n_658), .B(n_1331), .C(n_1332), .Y(n_1330) );
INVx3_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OAI22xp5_ASAP7_75t_SL g1359 ( .A1(n_659), .A2(n_911), .B1(n_1360), .B2(n_1363), .Y(n_1359) );
NAND3xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_665), .C(n_666), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_SL g682 ( .A(n_664), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g686 ( .A(n_666), .B(n_687), .C(n_690), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g1199 ( .A(n_666), .B(n_1200), .C(n_1201), .Y(n_1199) );
NAND3xp33_ASAP7_75t_L g1297 ( .A(n_666), .B(n_1298), .C(n_1299), .Y(n_1297) );
NAND3xp33_ASAP7_75t_L g1333 ( .A(n_666), .B(n_1334), .C(n_1335), .Y(n_1333) );
INVx1_ASAP7_75t_L g1662 ( .A(n_666), .Y(n_1662) );
XOR2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_715), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_694), .C(n_704), .Y(n_668) );
AND4x1_ASAP7_75t_L g669 ( .A(n_670), .B(n_676), .C(n_680), .D(n_686), .Y(n_669) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g1036 ( .A(n_688), .Y(n_1036) );
INVx2_ASAP7_75t_L g1166 ( .A(n_688), .Y(n_1166) );
BUFx3_ASAP7_75t_L g1242 ( .A(n_688), .Y(n_1242) );
INVx1_ASAP7_75t_L g1032 ( .A(n_689), .Y(n_1032) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx3_ASAP7_75t_L g1678 ( .A(n_693), .Y(n_1678) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OR2x6_ASAP7_75t_L g818 ( .A(n_699), .B(n_801), .Y(n_818) );
INVx2_ASAP7_75t_L g1268 ( .A(n_709), .Y(n_1268) );
INVx1_ASAP7_75t_L g1313 ( .A(n_709), .Y(n_1313) );
INVx1_ASAP7_75t_L g855 ( .A(n_716), .Y(n_855) );
XNOR2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_772), .Y(n_716) );
INVx1_ASAP7_75t_L g771 ( .A(n_718), .Y(n_771) );
NAND4xp25_ASAP7_75t_SL g739 ( .A(n_740), .B(n_745), .C(n_754), .D(n_763), .Y(n_739) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g1160 ( .A(n_749), .Y(n_1160) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g794 ( .A(n_750), .Y(n_794) );
BUFx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_753), .B(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g907 ( .A(n_762), .Y(n_907) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AOI222xp33_ASAP7_75t_L g819 ( .A1(n_779), .A2(n_820), .B1(n_821), .B2(n_822), .C1(n_823), .C2(n_824), .Y(n_819) );
OAI21xp5_ASAP7_75t_SL g812 ( .A1(n_782), .A2(n_813), .B(n_814), .Y(n_812) );
NAND3xp33_ASAP7_75t_L g785 ( .A(n_786), .B(n_795), .C(n_819), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_788), .B1(n_790), .B2(n_791), .Y(n_786) );
INVx2_ASAP7_75t_L g793 ( .A(n_789), .Y(n_793) );
AND2x4_ASAP7_75t_L g791 ( .A(n_792), .B(n_794), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NOR3xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_811), .C(n_817), .Y(n_795) );
NAND2x1p5_ASAP7_75t_L g797 ( .A(n_798), .B(n_800), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
OR2x6_ASAP7_75t_L g804 ( .A(n_801), .B(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g826 ( .A(n_801), .Y(n_826) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_810), .Y(n_806) );
OAI221xp5_ASAP7_75t_SL g831 ( .A1(n_809), .A2(n_832), .B1(n_834), .B2(n_836), .C(n_837), .Y(n_831) );
OAI22xp33_ASAP7_75t_L g934 ( .A1(n_813), .A2(n_935), .B1(n_936), .B2(n_937), .Y(n_934) );
OAI22xp33_ASAP7_75t_SL g940 ( .A1(n_813), .A2(n_941), .B1(n_942), .B2(n_944), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_813), .A2(n_1000), .B1(n_1001), .B2(n_1002), .Y(n_999) );
INVx1_ASAP7_75t_L g1056 ( .A(n_813), .Y(n_1056) );
OAI22xp33_ASAP7_75t_L g1670 ( .A1(n_813), .A2(n_1053), .B1(n_1671), .B2(n_1672), .Y(n_1670) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
OAI221xp5_ASAP7_75t_SL g843 ( .A1(n_820), .A2(n_822), .B1(n_844), .B2(n_847), .C(n_850), .Y(n_843) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
CKINVDCx8_ASAP7_75t_R g828 ( .A(n_829), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_842), .B1(n_843), .B2(n_853), .Y(n_830) );
BUFx2_ASAP7_75t_L g1030 ( .A(n_832), .Y(n_1030) );
INVx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
BUFx3_ASAP7_75t_L g949 ( .A(n_834), .Y(n_949) );
INVx1_ASAP7_75t_L g1082 ( .A(n_834), .Y(n_1082) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
BUFx2_ASAP7_75t_L g849 ( .A(n_835), .Y(n_849) );
BUFx4f_ASAP7_75t_L g1009 ( .A(n_835), .Y(n_1009) );
INVx1_ASAP7_75t_L g1022 ( .A(n_835), .Y(n_1022) );
INVx2_ASAP7_75t_SL g838 ( .A(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
BUFx2_ASAP7_75t_L g1110 ( .A(n_840), .Y(n_1110) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g1243 ( .A(n_841), .Y(n_1243) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx2_ASAP7_75t_L g948 ( .A(n_846), .Y(n_948) );
INVx2_ASAP7_75t_L g1005 ( .A(n_846), .Y(n_1005) );
INVx2_ASAP7_75t_L g1361 ( .A(n_846), .Y(n_1361) );
HB1xp67_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
OAI221xp5_ASAP7_75t_L g1363 ( .A1(n_848), .A2(n_1005), .B1(n_1364), .B2(n_1365), .C(n_1366), .Y(n_1363) );
INVx2_ASAP7_75t_SL g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
XNOR2x2_ASAP7_75t_L g857 ( .A(n_858), .B(n_918), .Y(n_857) );
XNOR2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g1419 ( .A1(n_859), .A2(n_1399), .B1(n_1404), .B2(n_1420), .Y(n_1419) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
NAND4xp25_ASAP7_75t_L g886 ( .A(n_887), .B(n_894), .C(n_901), .D(n_909), .Y(n_886) );
NAND3xp33_ASAP7_75t_L g887 ( .A(n_888), .B(n_891), .C(n_892), .Y(n_887) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx2_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
INVxp67_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
NAND3xp33_ASAP7_75t_L g901 ( .A(n_902), .B(n_903), .C(n_908), .Y(n_901) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g1659 ( .A1(n_905), .A2(n_1028), .B1(n_1660), .B2(n_1661), .Y(n_1659) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx2_ASAP7_75t_SL g1026 ( .A(n_906), .Y(n_1026) );
NAND3xp33_ASAP7_75t_L g909 ( .A(n_910), .B(n_912), .C(n_917), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
OAI22xp5_ASAP7_75t_SL g945 ( .A1(n_911), .A2(n_946), .B1(n_947), .B2(n_951), .Y(n_945) );
OAI22xp5_ASAP7_75t_SL g1003 ( .A1(n_911), .A2(n_946), .B1(n_1004), .B2(n_1007), .Y(n_1003) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx2_ASAP7_75t_SL g914 ( .A(n_915), .Y(n_914) );
XNOR2xp5_ASAP7_75t_L g918 ( .A(n_919), .B(n_920), .Y(n_918) );
NAND3x1_ASAP7_75t_SL g920 ( .A(n_921), .B(n_932), .C(n_955), .Y(n_920) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
AOI21xp5_ASAP7_75t_L g1265 ( .A1(n_925), .A2(n_1266), .B(n_1267), .Y(n_1265) );
AOI21xp5_ASAP7_75t_L g1310 ( .A1(n_925), .A2(n_1311), .B(n_1312), .Y(n_1310) );
OAI221xp5_ASAP7_75t_L g947 ( .A1(n_935), .A2(n_937), .B1(n_948), .B2(n_949), .C(n_950), .Y(n_947) );
OAI22xp33_ASAP7_75t_L g1354 ( .A1(n_936), .A2(n_1355), .B1(n_1356), .B2(n_1357), .Y(n_1354) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_942), .A2(n_990), .B1(n_991), .B2(n_992), .Y(n_989) );
INVx3_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
OAI33xp33_ASAP7_75t_L g1644 ( .A1(n_946), .A2(n_1645), .A3(n_1650), .B1(n_1656), .B2(n_1659), .B3(n_1662), .Y(n_1644) );
OAI221xp5_ASAP7_75t_L g951 ( .A1(n_948), .A2(n_949), .B1(n_952), .B2(n_953), .C(n_954), .Y(n_951) );
OAI221xp5_ASAP7_75t_L g1004 ( .A1(n_949), .A2(n_1000), .B1(n_1002), .B2(n_1005), .C(n_1006), .Y(n_1004) );
BUFx2_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
XNOR2xp5_ASAP7_75t_L g963 ( .A(n_964), .B(n_1126), .Y(n_963) );
XOR2x2_ASAP7_75t_SL g964 ( .A(n_965), .B(n_1011), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
NAND3x1_ASAP7_75t_L g968 ( .A(n_969), .B(n_976), .C(n_985), .Y(n_968) );
OAI221xp5_ASAP7_75t_L g1007 ( .A1(n_979), .A2(n_982), .B1(n_1005), .B2(n_1008), .C(n_1010), .Y(n_1007) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVx2_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
BUFx3_ASAP7_75t_L g1072 ( .A(n_994), .Y(n_1072) );
OAI22xp33_ASAP7_75t_L g1343 ( .A1(n_994), .A2(n_1001), .B1(n_1344), .B2(n_1345), .Y(n_1343) );
OAI22xp33_ASAP7_75t_L g1664 ( .A1(n_994), .A2(n_1053), .B1(n_1651), .B2(n_1654), .Y(n_1664) );
BUFx6f_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g1050 ( .A(n_998), .Y(n_1050) );
OAI22xp33_ASAP7_75t_SL g1346 ( .A1(n_998), .A2(n_1347), .B1(n_1348), .B2(n_1349), .Y(n_1346) );
INVx1_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
INVx2_ASAP7_75t_L g1655 ( .A(n_1009), .Y(n_1655) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
AOI22xp5_ASAP7_75t_L g1012 ( .A1(n_1013), .A2(n_1084), .B1(n_1085), .B2(n_1125), .Y(n_1012) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1013), .Y(n_1125) );
NAND3xp33_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1069), .C(n_1077), .Y(n_1014) );
NOR2xp33_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1039), .Y(n_1015) );
OAI221xp5_ASAP7_75t_L g1017 ( .A1(n_1018), .A2(n_1019), .B1(n_1020), .B2(n_1023), .C(n_1024), .Y(n_1017) );
OAI22xp33_ASAP7_75t_L g1052 ( .A1(n_1018), .A2(n_1023), .B1(n_1053), .B2(n_1055), .Y(n_1052) );
OAI221xp5_ASAP7_75t_L g1360 ( .A1(n_1020), .A2(n_1344), .B1(n_1345), .B2(n_1361), .C(n_1362), .Y(n_1360) );
INVx2_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
OAI221xp5_ASAP7_75t_L g1029 ( .A1(n_1030), .A2(n_1031), .B1(n_1032), .B2(n_1033), .C(n_1034), .Y(n_1029) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
OAI33xp33_ASAP7_75t_L g1039 ( .A1(n_1040), .A2(n_1044), .A3(n_1052), .B1(n_1057), .B2(n_1063), .B3(n_1068), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
OAI33xp33_ASAP7_75t_L g1342 ( .A1(n_1042), .A2(n_1343), .A3(n_1346), .B1(n_1350), .B2(n_1354), .B3(n_1358), .Y(n_1342) );
OAI33xp33_ASAP7_75t_L g1663 ( .A1(n_1042), .A2(n_1358), .A3(n_1664), .B1(n_1665), .B2(n_1666), .B3(n_1670), .Y(n_1663) );
OAI22xp5_ASAP7_75t_L g1044 ( .A1(n_1045), .A2(n_1046), .B1(n_1049), .B2(n_1051), .Y(n_1044) );
INVx2_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
BUFx3_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
OAI22xp33_ASAP7_75t_L g1057 ( .A1(n_1053), .A2(n_1058), .B1(n_1059), .B2(n_1062), .Y(n_1057) );
INVx2_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
HB1xp67_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
INVx2_ASAP7_75t_L g1348 ( .A(n_1061), .Y(n_1348) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1061), .Y(n_1667) );
OAI22xp33_ASAP7_75t_L g1063 ( .A1(n_1064), .A2(n_1065), .B1(n_1066), .B2(n_1067), .Y(n_1063) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
INVx2_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1086), .Y(n_1124) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1107), .Y(n_1100) );
NAND3xp33_ASAP7_75t_L g1190 ( .A(n_1106), .B(n_1191), .C(n_1193), .Y(n_1190) );
NAND3xp33_ASAP7_75t_L g1287 ( .A(n_1106), .B(n_1288), .C(n_1291), .Y(n_1287) );
NAND3xp33_ASAP7_75t_L g1327 ( .A(n_1106), .B(n_1328), .C(n_1329), .Y(n_1327) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1106), .Y(n_1358) );
AOI31xp33_ASAP7_75t_L g1113 ( .A1(n_1114), .A2(n_1117), .A3(n_1120), .B(n_1122), .Y(n_1113) );
AO21x1_ASAP7_75t_SL g1143 ( .A1(n_1122), .A2(n_1144), .B(n_1147), .Y(n_1143) );
AOI31xp33_ASAP7_75t_L g1273 ( .A1(n_1122), .A2(n_1274), .A3(n_1277), .B(n_1280), .Y(n_1273) );
AOI31xp33_ASAP7_75t_L g1314 ( .A1(n_1122), .A2(n_1315), .A3(n_1318), .B(n_1321), .Y(n_1314) );
XOR2xp5_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1254), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_1128), .A2(n_1129), .B1(n_1214), .B2(n_1215), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
AO22x2_ASAP7_75t_L g1129 ( .A1(n_1130), .A2(n_1172), .B1(n_1173), .B2(n_1213), .Y(n_1129) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1130), .Y(n_1213) );
NAND4xp25_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1143), .C(n_1150), .D(n_1163), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1139), .Y(n_1133) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
INVx2_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
NAND4xp25_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1190), .C(n_1194), .D(n_1199), .Y(n_1186) );
INVx2_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
INVx2_ASAP7_75t_SL g1296 ( .A(n_1198), .Y(n_1296) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1217), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1236), .Y(n_1230) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
OAI22xp5_ASAP7_75t_L g1256 ( .A1(n_1257), .A2(n_1258), .B1(n_1300), .B2(n_1301), .Y(n_1256) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
XNOR2xp5_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1260), .Y(n_1258) );
NAND4xp25_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1287), .C(n_1292), .D(n_1297), .Y(n_1282) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
NAND4xp25_ASAP7_75t_L g1323 ( .A(n_1324), .B(n_1327), .C(n_1330), .D(n_1333), .Y(n_1323) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1336), .Y(n_1380) );
INVx2_ASAP7_75t_SL g1336 ( .A(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
NAND3xp33_ASAP7_75t_L g1340 ( .A(n_1341), .B(n_1367), .C(n_1375), .Y(n_1340) );
NOR2xp33_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1359), .Y(n_1341) );
OAI22xp5_ASAP7_75t_L g1350 ( .A1(n_1348), .A2(n_1351), .B1(n_1352), .B2(n_1353), .Y(n_1350) );
OAI22xp33_ASAP7_75t_L g1665 ( .A1(n_1348), .A2(n_1352), .B1(n_1646), .B2(n_1648), .Y(n_1665) );
OAI22xp33_ASAP7_75t_L g1666 ( .A1(n_1352), .A2(n_1667), .B1(n_1668), .B2(n_1669), .Y(n_1666) );
OAI221xp5_ASAP7_75t_L g1381 ( .A1(n_1382), .A2(n_1635), .B1(n_1638), .B2(n_1686), .C(n_1692), .Y(n_1381) );
NOR3xp33_ASAP7_75t_L g1382 ( .A(n_1383), .B(n_1546), .C(n_1592), .Y(n_1382) );
AOI21xp5_ASAP7_75t_L g1383 ( .A1(n_1384), .A2(n_1497), .B(n_1536), .Y(n_1383) );
AOI221xp5_ASAP7_75t_L g1384 ( .A1(n_1385), .A2(n_1430), .B1(n_1446), .B2(n_1452), .C(n_1460), .Y(n_1384) );
INVxp67_ASAP7_75t_SL g1385 ( .A(n_1386), .Y(n_1385) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_1387), .B(n_1406), .Y(n_1386) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1387), .Y(n_1518) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1387), .Y(n_1554) );
NAND2xp5_ASAP7_75t_L g1565 ( .A(n_1387), .B(n_1549), .Y(n_1565) );
HB1xp67_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
INVx2_ASAP7_75t_SL g1450 ( .A(n_1388), .Y(n_1450) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_1388), .B(n_1443), .Y(n_1495) );
OR2x2_ASAP7_75t_L g1502 ( .A(n_1388), .B(n_1443), .Y(n_1502) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1389), .Y(n_1440) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1389), .Y(n_1539) );
AND2x4_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1393), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1390), .B(n_1393), .Y(n_1417) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
AND2x4_ASAP7_75t_L g1395 ( .A(n_1391), .B(n_1393), .Y(n_1395) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1401 ( .A(n_1392), .B(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1394), .Y(n_1402) );
INVx1_ASAP7_75t_SL g1425 ( .A(n_1395), .Y(n_1425) );
INVx2_ASAP7_75t_L g1458 ( .A(n_1395), .Y(n_1458) );
OAI22xp33_ASAP7_75t_L g1396 ( .A1(n_1397), .A2(n_1398), .B1(n_1403), .B2(n_1404), .Y(n_1396) );
OAI22xp5_ASAP7_75t_L g1427 ( .A1(n_1398), .A2(n_1404), .B1(n_1428), .B2(n_1429), .Y(n_1427) );
OAI22xp33_ASAP7_75t_L g1433 ( .A1(n_1398), .A2(n_1434), .B1(n_1435), .B2(n_1436), .Y(n_1433) );
BUFx3_ASAP7_75t_L g1543 ( .A(n_1398), .Y(n_1543) );
BUFx6f_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
OR2x2_ASAP7_75t_L g1399 ( .A(n_1400), .B(n_1401), .Y(n_1399) );
OR2x2_ASAP7_75t_L g1404 ( .A(n_1400), .B(n_1405), .Y(n_1404) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1400), .Y(n_1413) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1401), .Y(n_1412) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1404), .Y(n_1437) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1405), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1421), .Y(n_1406) );
NAND2xp5_ASAP7_75t_L g1520 ( .A(n_1407), .B(n_1453), .Y(n_1520) );
NAND2xp5_ASAP7_75t_L g1532 ( .A(n_1407), .B(n_1487), .Y(n_1532) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
NOR2xp33_ASAP7_75t_L g1479 ( .A(n_1408), .B(n_1464), .Y(n_1479) );
OR2x2_ASAP7_75t_L g1568 ( .A(n_1408), .B(n_1421), .Y(n_1568) );
OR2x2_ASAP7_75t_L g1617 ( .A(n_1408), .B(n_1454), .Y(n_1617) );
OR2x2_ASAP7_75t_L g1408 ( .A(n_1409), .B(n_1418), .Y(n_1408) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1409), .Y(n_1467) );
AND2x2_ASAP7_75t_L g1472 ( .A(n_1409), .B(n_1421), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1409), .B(n_1485), .Y(n_1484) );
AND2x2_ASAP7_75t_L g1525 ( .A(n_1409), .B(n_1418), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1410), .B(n_1416), .Y(n_1409) );
AND2x4_ASAP7_75t_L g1411 ( .A(n_1412), .B(n_1413), .Y(n_1411) );
AND2x4_ASAP7_75t_L g1414 ( .A(n_1413), .B(n_1415), .Y(n_1414) );
HB1xp67_ASAP7_75t_L g1703 ( .A(n_1415), .Y(n_1703) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1417), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1452 ( .A(n_1418), .B(n_1453), .Y(n_1452) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_1418), .B(n_1467), .Y(n_1466) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1418), .Y(n_1485) );
NOR2xp33_ASAP7_75t_L g1598 ( .A(n_1418), .B(n_1459), .Y(n_1598) );
CKINVDCx6p67_ASAP7_75t_R g1459 ( .A(n_1421), .Y(n_1459) );
NAND2xp5_ASAP7_75t_L g1478 ( .A(n_1421), .B(n_1479), .Y(n_1478) );
OAI331xp33_ASAP7_75t_L g1498 ( .A1(n_1421), .A2(n_1485), .A3(n_1499), .B1(n_1503), .B2(n_1506), .B3(n_1508), .C1(n_1510), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1535 ( .A(n_1421), .B(n_1484), .Y(n_1535) );
AND2x2_ASAP7_75t_L g1551 ( .A(n_1421), .B(n_1466), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1421), .B(n_1467), .Y(n_1581) );
OR2x2_ASAP7_75t_L g1588 ( .A(n_1421), .B(n_1467), .Y(n_1588) );
OR2x6_ASAP7_75t_SL g1421 ( .A(n_1422), .B(n_1427), .Y(n_1421) );
OAI22xp5_ASAP7_75t_L g1422 ( .A1(n_1423), .A2(n_1424), .B1(n_1425), .B2(n_1426), .Y(n_1422) );
OAI22xp5_ASAP7_75t_L g1438 ( .A1(n_1425), .A2(n_1439), .B1(n_1440), .B2(n_1441), .Y(n_1438) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1430), .Y(n_1521) );
A2O1A1Ixp33_ASAP7_75t_SL g1624 ( .A1(n_1430), .A2(n_1607), .B(n_1625), .C(n_1626), .Y(n_1624) );
AND2x2_ASAP7_75t_L g1430 ( .A(n_1431), .B(n_1442), .Y(n_1430) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1431), .Y(n_1451) );
AND2x2_ASAP7_75t_L g1489 ( .A(n_1431), .B(n_1474), .Y(n_1489) );
OR2x2_ASAP7_75t_L g1512 ( .A(n_1431), .B(n_1443), .Y(n_1512) );
AND2x2_ASAP7_75t_L g1516 ( .A(n_1431), .B(n_1443), .Y(n_1516) );
AND2x2_ASAP7_75t_L g1528 ( .A(n_1431), .B(n_1495), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1548 ( .A(n_1431), .B(n_1450), .Y(n_1548) );
NAND2xp5_ASAP7_75t_L g1583 ( .A(n_1431), .B(n_1536), .Y(n_1583) );
INVx3_ASAP7_75t_L g1612 ( .A(n_1431), .Y(n_1612) );
INVx3_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
AND2x2_ASAP7_75t_L g1475 ( .A(n_1432), .B(n_1443), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1432), .B(n_1454), .Y(n_1509) );
OR2x2_ASAP7_75t_L g1633 ( .A(n_1432), .B(n_1502), .Y(n_1633) );
OR2x2_ASAP7_75t_L g1432 ( .A(n_1433), .B(n_1438), .Y(n_1432) );
HB1xp67_ASAP7_75t_L g1545 ( .A(n_1436), .Y(n_1545) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
OAI211xp5_ASAP7_75t_SL g1460 ( .A1(n_1442), .A2(n_1461), .B(n_1468), .C(n_1490), .Y(n_1460) );
AOI22xp33_ASAP7_75t_SL g1601 ( .A1(n_1442), .A2(n_1567), .B1(n_1602), .B2(n_1606), .Y(n_1601) );
O2A1O1Ixp33_ASAP7_75t_L g1606 ( .A1(n_1442), .A2(n_1464), .B(n_1495), .C(n_1551), .Y(n_1606) );
INVx2_ASAP7_75t_L g1442 ( .A(n_1443), .Y(n_1442) );
OR2x2_ASAP7_75t_L g1449 ( .A(n_1443), .B(n_1450), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1507 ( .A(n_1443), .B(n_1450), .Y(n_1507) );
OAI22xp5_ASAP7_75t_L g1552 ( .A1(n_1443), .A2(n_1488), .B1(n_1553), .B2(n_1555), .Y(n_1552) );
AND2x4_ASAP7_75t_L g1443 ( .A(n_1444), .B(n_1445), .Y(n_1443) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
NAND2xp5_ASAP7_75t_L g1447 ( .A(n_1448), .B(n_1451), .Y(n_1447) );
NAND2xp5_ASAP7_75t_L g1623 ( .A(n_1448), .B(n_1550), .Y(n_1623) );
INVx2_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
OR2x2_ASAP7_75t_L g1614 ( .A(n_1449), .B(n_1550), .Y(n_1614) );
INVx2_ASAP7_75t_SL g1474 ( .A(n_1450), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1491 ( .A(n_1451), .B(n_1492), .Y(n_1491) );
NAND2xp5_ASAP7_75t_L g1481 ( .A(n_1453), .B(n_1466), .Y(n_1481) );
NAND2xp5_ASAP7_75t_L g1576 ( .A(n_1453), .B(n_1525), .Y(n_1576) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1454), .B(n_1459), .Y(n_1453) );
INVx4_ASAP7_75t_L g1464 ( .A(n_1454), .Y(n_1464) );
INVx2_ASAP7_75t_L g1471 ( .A(n_1454), .Y(n_1471) );
NOR2xp33_ASAP7_75t_L g1487 ( .A(n_1454), .B(n_1459), .Y(n_1487) );
NAND2xp5_ASAP7_75t_L g1557 ( .A(n_1454), .B(n_1525), .Y(n_1557) );
OR2x2_ASAP7_75t_L g1567 ( .A(n_1454), .B(n_1568), .Y(n_1567) );
AOI322xp5_ASAP7_75t_L g1571 ( .A1(n_1454), .A2(n_1495), .A3(n_1501), .B1(n_1507), .B2(n_1572), .C1(n_1575), .C2(n_1577), .Y(n_1571) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_1454), .B(n_1507), .Y(n_1600) );
AND2x6_ASAP7_75t_L g1454 ( .A(n_1455), .B(n_1456), .Y(n_1454) );
INVx2_ASAP7_75t_L g1457 ( .A(n_1458), .Y(n_1457) );
OAI22xp5_ASAP7_75t_L g1537 ( .A1(n_1458), .A2(n_1538), .B1(n_1539), .B2(n_1540), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_1459), .B(n_1466), .Y(n_1465) );
AND2x2_ASAP7_75t_L g1496 ( .A(n_1459), .B(n_1484), .Y(n_1496) );
AND2x2_ASAP7_75t_L g1523 ( .A(n_1459), .B(n_1524), .Y(n_1523) );
NOR2xp33_ASAP7_75t_L g1556 ( .A(n_1459), .B(n_1557), .Y(n_1556) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1459), .B(n_1485), .Y(n_1603) );
OR2x2_ASAP7_75t_L g1628 ( .A(n_1459), .B(n_1485), .Y(n_1628) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
NAND2xp5_ASAP7_75t_L g1463 ( .A(n_1464), .B(n_1465), .Y(n_1463) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1464), .Y(n_1494) );
AND2x2_ASAP7_75t_L g1500 ( .A(n_1464), .B(n_1501), .Y(n_1500) );
AND2x2_ASAP7_75t_L g1513 ( .A(n_1464), .B(n_1496), .Y(n_1513) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1464), .B(n_1525), .Y(n_1524) );
NOR2xp33_ASAP7_75t_L g1604 ( .A(n_1464), .B(n_1605), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1570 ( .A(n_1465), .B(n_1492), .Y(n_1570) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1466), .Y(n_1505) );
OAI22xp5_ASAP7_75t_SL g1619 ( .A1(n_1467), .A2(n_1620), .B1(n_1621), .B2(n_1623), .Y(n_1619) );
AOI211xp5_ASAP7_75t_L g1468 ( .A1(n_1469), .A2(n_1473), .B(n_1476), .C(n_1480), .Y(n_1468) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
NAND2xp5_ASAP7_75t_L g1470 ( .A(n_1471), .B(n_1472), .Y(n_1470) );
INVx2_ASAP7_75t_L g1550 ( .A(n_1471), .Y(n_1550) );
NAND2xp5_ASAP7_75t_L g1590 ( .A(n_1471), .B(n_1591), .Y(n_1590) );
OAI32xp33_ASAP7_75t_L g1602 ( .A1(n_1471), .A2(n_1495), .A3(n_1551), .B1(n_1603), .B2(n_1604), .Y(n_1602) );
AND2x2_ASAP7_75t_L g1473 ( .A(n_1474), .B(n_1475), .Y(n_1473) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1474), .Y(n_1477) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1474), .Y(n_1492) );
NOR2xp33_ASAP7_75t_L g1579 ( .A(n_1474), .B(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1474), .Y(n_1591) );
OAI22xp5_ASAP7_75t_L g1615 ( .A1(n_1474), .A2(n_1551), .B1(n_1616), .B2(n_1618), .Y(n_1615) );
NAND2xp5_ASAP7_75t_L g1616 ( .A(n_1474), .B(n_1617), .Y(n_1616) );
OAI21xp33_ASAP7_75t_L g1563 ( .A1(n_1475), .A2(n_1564), .B(n_1566), .Y(n_1563) );
NOR2xp33_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1478), .Y(n_1476) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1478), .Y(n_1560) );
AOI21xp33_ASAP7_75t_SL g1480 ( .A1(n_1481), .A2(n_1482), .B(n_1488), .Y(n_1480) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1481), .Y(n_1618) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1482), .Y(n_1584) );
OR2x2_ASAP7_75t_L g1482 ( .A(n_1483), .B(n_1486), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1504 ( .A(n_1483), .B(n_1505), .Y(n_1504) );
NOR2xp33_ASAP7_75t_L g1526 ( .A(n_1483), .B(n_1527), .Y(n_1526) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
NOR3xp33_ASAP7_75t_L g1630 ( .A(n_1485), .B(n_1550), .C(n_1631), .Y(n_1630) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
OAI21xp5_ASAP7_75t_L g1490 ( .A1(n_1491), .A2(n_1493), .B(n_1496), .Y(n_1490) );
AOI221xp5_ASAP7_75t_SL g1578 ( .A1(n_1491), .A2(n_1579), .B1(n_1582), .B2(n_1584), .C(n_1585), .Y(n_1578) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1494), .B(n_1495), .Y(n_1493) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1496), .Y(n_1574) );
NOR5xp2_ASAP7_75t_L g1497 ( .A(n_1498), .B(n_1514), .C(n_1526), .D(n_1529), .E(n_1533), .Y(n_1497) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
A2O1A1Ixp33_ASAP7_75t_L g1634 ( .A1(n_1500), .A2(n_1533), .B(n_1598), .C(n_1612), .Y(n_1634) );
INVx1_ASAP7_75t_L g1501 ( .A(n_1502), .Y(n_1501) );
NOR2xp33_ASAP7_75t_L g1533 ( .A(n_1502), .B(n_1534), .Y(n_1533) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
NOR2x1_ASAP7_75t_R g1562 ( .A(n_1505), .B(n_1550), .Y(n_1562) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
NAND2xp5_ASAP7_75t_L g1530 ( .A(n_1507), .B(n_1531), .Y(n_1530) );
NAND2xp5_ASAP7_75t_L g1595 ( .A(n_1507), .B(n_1535), .Y(n_1595) );
INVxp67_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
NAND2xp5_ASAP7_75t_L g1510 ( .A(n_1511), .B(n_1513), .Y(n_1510) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
OAI22xp5_ASAP7_75t_SL g1514 ( .A1(n_1515), .A2(n_1517), .B1(n_1521), .B2(n_1522), .Y(n_1514) );
AOI21xp33_ASAP7_75t_L g1585 ( .A1(n_1515), .A2(n_1583), .B(n_1586), .Y(n_1585) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
AND2x2_ASAP7_75t_L g1626 ( .A(n_1516), .B(n_1627), .Y(n_1626) );
NAND2xp5_ASAP7_75t_L g1517 ( .A(n_1518), .B(n_1519), .Y(n_1517) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_1518), .B(n_1576), .Y(n_1620) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
OR2x2_ASAP7_75t_L g1553 ( .A(n_1520), .B(n_1554), .Y(n_1553) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
AOI21xp33_ASAP7_75t_L g1558 ( .A1(n_1527), .A2(n_1559), .B(n_1561), .Y(n_1558) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
INVx1_ASAP7_75t_L g1531 ( .A(n_1532), .Y(n_1531) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1536), .Y(n_1608) );
NAND2xp5_ASAP7_75t_L g1611 ( .A(n_1536), .B(n_1612), .Y(n_1611) );
CKINVDCx5p33_ASAP7_75t_R g1631 ( .A(n_1536), .Y(n_1631) );
OR2x6_ASAP7_75t_SL g1536 ( .A(n_1537), .B(n_1541), .Y(n_1536) );
OAI22xp5_ASAP7_75t_L g1541 ( .A1(n_1542), .A2(n_1543), .B1(n_1544), .B2(n_1545), .Y(n_1541) );
BUFx2_ASAP7_75t_SL g1637 ( .A(n_1545), .Y(n_1637) );
NAND4xp25_ASAP7_75t_L g1546 ( .A(n_1547), .B(n_1563), .C(n_1571), .D(n_1578), .Y(n_1546) );
AOI211xp5_ASAP7_75t_SL g1547 ( .A1(n_1548), .A2(n_1549), .B(n_1552), .C(n_1558), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1550), .B(n_1551), .Y(n_1549) );
NAND2xp5_ASAP7_75t_L g1580 ( .A(n_1550), .B(n_1581), .Y(n_1580) );
NOR2x1_ASAP7_75t_L g1627 ( .A(n_1550), .B(n_1628), .Y(n_1627) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1551), .Y(n_1573) );
OAI31xp33_ASAP7_75t_L g1629 ( .A1(n_1551), .A2(n_1577), .A3(n_1630), .B(n_1632), .Y(n_1629) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1556), .Y(n_1555) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1557), .Y(n_1625) );
INVxp67_ASAP7_75t_SL g1559 ( .A(n_1560), .Y(n_1559) );
INVxp33_ASAP7_75t_L g1561 ( .A(n_1562), .Y(n_1561) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
NAND2xp33_ASAP7_75t_L g1566 ( .A(n_1567), .B(n_1569), .Y(n_1566) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1567), .Y(n_1577) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1568), .Y(n_1622) );
INVxp33_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
NAND2xp5_ASAP7_75t_L g1572 ( .A(n_1573), .B(n_1574), .Y(n_1572) );
NOR2xp33_ASAP7_75t_L g1621 ( .A(n_1575), .B(n_1622), .Y(n_1621) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
AOI22xp5_ASAP7_75t_L g1609 ( .A1(n_1582), .A2(n_1610), .B1(n_1613), .B2(n_1619), .Y(n_1609) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
NAND2xp5_ASAP7_75t_L g1586 ( .A(n_1587), .B(n_1589), .Y(n_1586) );
OAI21xp5_ASAP7_75t_SL g1613 ( .A1(n_1587), .A2(n_1614), .B(n_1615), .Y(n_1613) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
NAND5xp2_ASAP7_75t_L g1592 ( .A(n_1593), .B(n_1609), .C(n_1624), .D(n_1629), .E(n_1634), .Y(n_1592) );
OAI31xp33_ASAP7_75t_SL g1593 ( .A1(n_1594), .A2(n_1596), .A3(n_1601), .B(n_1607), .Y(n_1593) );
INVxp67_ASAP7_75t_SL g1594 ( .A(n_1595), .Y(n_1594) );
NOR2xp33_ASAP7_75t_L g1596 ( .A(n_1597), .B(n_1599), .Y(n_1596) );
INVx1_ASAP7_75t_L g1597 ( .A(n_1598), .Y(n_1597) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1600), .Y(n_1599) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1603), .Y(n_1605) );
CKINVDCx14_ASAP7_75t_R g1607 ( .A(n_1608), .Y(n_1607) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
INVx1_ASAP7_75t_L g1632 ( .A(n_1633), .Y(n_1632) );
CKINVDCx5p33_ASAP7_75t_R g1635 ( .A(n_1636), .Y(n_1635) );
INVx1_ASAP7_75t_SL g1636 ( .A(n_1637), .Y(n_1636) );
HB1xp67_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
INVx2_ASAP7_75t_SL g1639 ( .A(n_1640), .Y(n_1639) );
HB1xp67_ASAP7_75t_L g1640 ( .A(n_1641), .Y(n_1640) );
HB1xp67_ASAP7_75t_L g1697 ( .A(n_1642), .Y(n_1697) );
NAND3xp33_ASAP7_75t_L g1642 ( .A(n_1643), .B(n_1673), .C(n_1681), .Y(n_1642) );
NOR2xp33_ASAP7_75t_L g1643 ( .A(n_1644), .B(n_1663), .Y(n_1643) );
OAI22xp5_ASAP7_75t_L g1645 ( .A1(n_1646), .A2(n_1647), .B1(n_1648), .B2(n_1649), .Y(n_1645) );
OAI22xp5_ASAP7_75t_L g1650 ( .A1(n_1651), .A2(n_1652), .B1(n_1654), .B2(n_1655), .Y(n_1650) );
OAI22xp5_ASAP7_75t_L g1656 ( .A1(n_1652), .A2(n_1655), .B1(n_1657), .B2(n_1658), .Y(n_1656) );
INVx2_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
CKINVDCx5p33_ASAP7_75t_R g1686 ( .A(n_1687), .Y(n_1686) );
CKINVDCx5p33_ASAP7_75t_R g1687 ( .A(n_1688), .Y(n_1687) );
INVx2_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1691), .Y(n_1690) );
INVxp33_ASAP7_75t_L g1693 ( .A(n_1694), .Y(n_1693) );
INVx1_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
BUFx2_ASAP7_75t_L g1698 ( .A(n_1699), .Y(n_1698) );
OAI21xp5_ASAP7_75t_L g1702 ( .A1(n_1700), .A2(n_1703), .B(n_1704), .Y(n_1702) );
BUFx2_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
endmodule