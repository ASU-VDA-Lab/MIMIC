module fake_jpeg_11371_n_593 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_593);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_593;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_455;
wire n_137;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_19),
.B(n_2),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_63),
.B(n_72),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_65),
.Y(n_188)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_19),
.B(n_3),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_67),
.B(n_103),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_68),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_69),
.Y(n_156)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_21),
.B(n_3),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_71),
.B(n_79),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_42),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_76),
.B(n_84),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_48),
.Y(n_78)
);

NAND2xp33_ASAP7_75t_SL g193 ( 
.A(n_78),
.B(n_39),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_21),
.B(n_3),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_80),
.Y(n_185)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_81),
.Y(n_171)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_82),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_83),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_42),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_85),
.Y(n_196)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

BUFx16f_ASAP7_75t_L g189 ( 
.A(n_87),
.Y(n_189)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_89),
.Y(n_163)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_91),
.Y(n_164)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_42),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_97),
.B(n_106),
.Y(n_174)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_98),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_99),
.Y(n_195)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_100),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_23),
.B(n_4),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_101),
.B(n_120),
.Y(n_169)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_102),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_23),
.B(n_17),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_104),
.Y(n_201)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_31),
.B(n_4),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_22),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_108),
.B(n_115),
.Y(n_183)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_109),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

CKINVDCx6p67_ASAP7_75t_R g172 ( 
.A(n_114),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_57),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_26),
.Y(n_116)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

BUFx4f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

BUFx8_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_119),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_31),
.B(n_4),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_32),
.B(n_6),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_20),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_53),
.B(n_35),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_122),
.B(n_124),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_44),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_41),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_46),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g167 ( 
.A(n_125),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_94),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_130),
.B(n_132),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_122),
.Y(n_132)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

INVx11_ASAP7_75t_L g215 ( 
.A(n_133),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_82),
.A2(n_98),
.B1(n_114),
.B2(n_60),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_140),
.A2(n_142),
.B1(n_168),
.B2(n_105),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_141),
.B(n_145),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_68),
.A2(n_38),
.B1(n_43),
.B2(n_46),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_78),
.B(n_32),
.Y(n_145)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

INVx5_ASAP7_75t_SL g251 ( 
.A(n_146),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_117),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_151),
.B(n_158),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_64),
.A2(n_125),
.B1(n_123),
.B2(n_77),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_152),
.A2(n_110),
.B1(n_99),
.B2(n_83),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_95),
.Y(n_158)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g227 ( 
.A(n_159),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_74),
.A2(n_43),
.B1(n_38),
.B2(n_46),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_109),
.B(n_36),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_175),
.B(n_197),
.Y(n_259)
);

INVx6_ASAP7_75t_SL g180 ( 
.A(n_85),
.Y(n_180)
);

CKINVDCx9p33_ASAP7_75t_R g239 ( 
.A(n_180),
.Y(n_239)
);

INVx11_ASAP7_75t_L g181 ( 
.A(n_87),
.Y(n_181)
);

BUFx2_ASAP7_75t_SL g262 ( 
.A(n_181),
.Y(n_262)
);

HAxp5_ASAP7_75t_SL g184 ( 
.A(n_65),
.B(n_20),
.CON(n_184),
.SN(n_184)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_184),
.A2(n_193),
.B(n_36),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_90),
.A2(n_39),
.B(n_58),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_187),
.B(n_203),
.Y(n_260)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_87),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_191),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_113),
.B(n_50),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_192),
.B(n_194),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_70),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_80),
.B(n_49),
.Y(n_197)
);

INVx11_ASAP7_75t_L g199 ( 
.A(n_81),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_199),
.Y(n_208)
);

INVx6_ASAP7_75t_SL g203 ( 
.A(n_92),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_96),
.B(n_49),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_207),
.B(n_12),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_183),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_209),
.B(n_237),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_210),
.B(n_260),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_150),
.B(n_47),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_211),
.B(n_220),
.Y(n_301)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_154),
.Y(n_213)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_213),
.Y(n_303)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_135),
.Y(n_214)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_214),
.Y(n_296)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_135),
.Y(n_217)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_217),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_154),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_218),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_219),
.A2(n_223),
.B1(n_230),
.B2(n_231),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_47),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_221),
.Y(n_281)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_222),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_168),
.A2(n_104),
.B1(n_112),
.B2(n_107),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_126),
.B(n_169),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_224),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_184),
.A2(n_27),
.B1(n_59),
.B2(n_58),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_225),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_166),
.B(n_27),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_226),
.Y(n_327)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_143),
.Y(n_228)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_228),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_229),
.A2(n_139),
.B1(n_176),
.B2(n_195),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_142),
.A2(n_69),
.B1(n_38),
.B2(n_43),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_128),
.A2(n_45),
.B1(n_55),
.B2(n_50),
.Y(n_231)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_155),
.Y(n_233)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_233),
.Y(n_295)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_153),
.Y(n_235)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_235),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_140),
.A2(n_53),
.B1(n_55),
.B2(n_45),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_236),
.A2(n_196),
.B1(n_170),
.B2(n_190),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_160),
.B(n_59),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_178),
.B(n_53),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_238),
.B(n_243),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_240),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_136),
.A2(n_53),
.B1(n_56),
.B2(n_52),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_241),
.A2(n_271),
.B1(n_272),
.B2(n_274),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_56),
.Y(n_242)
);

XNOR2x1_ASAP7_75t_L g312 ( 
.A(n_242),
.B(n_247),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_179),
.B(n_52),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_163),
.Y(n_244)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_244),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_133),
.Y(n_245)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_245),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_146),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_246),
.B(n_253),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_41),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g248 ( 
.A(n_204),
.Y(n_248)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

BUFx12f_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_249),
.Y(n_334)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_148),
.Y(n_250)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_156),
.Y(n_252)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_252),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_193),
.B(n_6),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_172),
.B(n_7),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_254),
.B(n_261),
.Y(n_307)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_164),
.Y(n_255)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_255),
.Y(n_305)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_156),
.Y(n_257)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_148),
.Y(n_258)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_258),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_172),
.B(n_7),
.Y(n_261)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_165),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_263),
.B(n_266),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_152),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_265)
);

OA21x2_ASAP7_75t_L g333 ( 
.A1(n_265),
.A2(n_269),
.B(n_127),
.Y(n_333)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_177),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_144),
.Y(n_267)
);

INVx11_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_129),
.B(n_8),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_268),
.B(n_270),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_136),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_198),
.Y(n_270)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_165),
.Y(n_271)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_148),
.Y(n_273)
);

INVx11_ASAP7_75t_L g322 ( 
.A(n_273),
.Y(n_322)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_167),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_172),
.B(n_12),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_275),
.Y(n_328)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_144),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_276),
.A2(n_278),
.B1(n_185),
.B2(n_182),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_200),
.B(n_138),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_274),
.Y(n_292)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_182),
.Y(n_278)
);

O2A1O1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_239),
.A2(n_159),
.B(n_181),
.C(n_191),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_279),
.B(n_284),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_212),
.B(n_187),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_280),
.B(n_285),
.C(n_286),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_196),
.B(n_127),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_242),
.B(n_247),
.C(n_259),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_242),
.B(n_131),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_292),
.B(n_248),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_253),
.A2(n_268),
.B(n_232),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_300),
.B(n_318),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_233),
.B(n_134),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_310),
.B(n_317),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_313),
.A2(n_330),
.B1(n_304),
.B2(n_271),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_247),
.B(n_188),
.C(n_199),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_314),
.B(n_325),
.C(n_208),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_244),
.B(n_134),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_234),
.A2(n_265),
.B(n_239),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_321),
.B(n_167),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_229),
.A2(n_206),
.B1(n_201),
.B2(n_162),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_323),
.A2(n_326),
.B1(n_331),
.B2(n_333),
.Y(n_358)
);

INVx3_ASAP7_75t_SL g367 ( 
.A(n_324),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_255),
.B(n_188),
.C(n_190),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_230),
.A2(n_139),
.B1(n_176),
.B2(n_195),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_223),
.A2(n_186),
.B1(n_149),
.B2(n_206),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_269),
.A2(n_162),
.B1(n_201),
.B2(n_149),
.Y(n_331)
);

AND2x6_ASAP7_75t_L g335 ( 
.A(n_297),
.B(n_264),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_335),
.B(n_345),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_280),
.B(n_270),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_341),
.Y(n_378)
);

INVx13_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_340),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_297),
.B(n_266),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_308),
.Y(n_342)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_342),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_306),
.Y(n_343)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_343),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_297),
.B(n_217),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_344),
.B(n_351),
.Y(n_392)
);

AND2x6_ASAP7_75t_L g345 ( 
.A(n_285),
.B(n_251),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_346),
.B(n_347),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_301),
.B(n_216),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_295),
.Y(n_348)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_348),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_216),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_349),
.Y(n_382)
);

AO22x1_ASAP7_75t_L g350 ( 
.A1(n_311),
.A2(n_236),
.B1(n_251),
.B2(n_221),
.Y(n_350)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_290),
.B(n_214),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_295),
.Y(n_352)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_352),
.Y(n_397)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_309),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_353),
.Y(n_398)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_302),
.Y(n_354)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_354),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_355),
.B(n_377),
.Y(n_407)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_282),
.Y(n_356)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_356),
.Y(n_406)
);

AND2x6_ASAP7_75t_L g357 ( 
.A(n_284),
.B(n_215),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_362),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_288),
.B(n_216),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_359),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_323),
.A2(n_186),
.B1(n_222),
.B2(n_170),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_360),
.A2(n_366),
.B1(n_369),
.B2(n_331),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_312),
.B(n_256),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_361),
.B(n_368),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_307),
.B(n_257),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_302),
.Y(n_363)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_363),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_289),
.B(n_249),
.Y(n_364)
);

AO21x1_ASAP7_75t_L g414 ( 
.A1(n_364),
.A2(n_374),
.B(n_375),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_292),
.B(n_213),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_305),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_370),
.A2(n_245),
.B1(n_293),
.B2(n_250),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_311),
.A2(n_278),
.B1(n_258),
.B2(n_273),
.Y(n_371)
);

OAI22x1_ASAP7_75t_L g408 ( 
.A1(n_371),
.A2(n_215),
.B1(n_322),
.B2(n_291),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_304),
.A2(n_252),
.B1(n_263),
.B2(n_218),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_372),
.A2(n_279),
.B1(n_316),
.B2(n_303),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_320),
.B(n_276),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_376),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_289),
.B(n_248),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_327),
.B(n_249),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_327),
.B(n_299),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_286),
.B(n_267),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_358),
.A2(n_313),
.B1(n_318),
.B2(n_319),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_379),
.A2(n_381),
.B1(n_387),
.B2(n_394),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_358),
.A2(n_333),
.B1(n_298),
.B2(n_314),
.Y(n_381)
);

OAI32xp33_ASAP7_75t_L g383 ( 
.A1(n_341),
.A2(n_333),
.A3(n_310),
.B1(n_317),
.B2(n_312),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_383),
.B(n_377),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_386),
.A2(n_390),
.B1(n_396),
.B2(n_343),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_337),
.A2(n_300),
.B1(n_325),
.B2(n_306),
.Y(n_387)
);

OAI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_342),
.A2(n_299),
.B1(n_294),
.B2(n_316),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_337),
.A2(n_294),
.B1(n_303),
.B2(n_332),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_395),
.A2(n_404),
.B1(n_315),
.B2(n_296),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_372),
.A2(n_283),
.B1(n_305),
.B2(n_282),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_336),
.A2(n_334),
.B(n_309),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_399),
.A2(n_400),
.B(n_370),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_336),
.A2(n_334),
.B(n_256),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_339),
.A2(n_332),
.B1(n_281),
.B2(n_283),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_365),
.A2(n_329),
.B1(n_291),
.B2(n_293),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_405),
.A2(n_412),
.B(n_350),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g436 ( 
.A1(n_408),
.A2(n_367),
.B1(n_182),
.B2(n_185),
.Y(n_436)
);

OA21x2_ASAP7_75t_L g412 ( 
.A1(n_336),
.A2(n_329),
.B(n_315),
.Y(n_412)
);

OAI22xp33_ASAP7_75t_SL g421 ( 
.A1(n_413),
.A2(n_367),
.B1(n_353),
.B2(n_208),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g415 ( 
.A1(n_389),
.A2(n_369),
.B1(n_365),
.B2(n_366),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_415),
.A2(n_405),
.B1(n_400),
.B2(n_399),
.Y(n_461)
);

AO22x1_ASAP7_75t_SL g416 ( 
.A1(n_389),
.A2(n_383),
.B1(n_357),
.B2(n_412),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_416),
.B(n_442),
.Y(n_450)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_388),
.Y(n_417)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_417),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_407),
.B(n_338),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_418),
.B(n_422),
.C(n_428),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_419),
.A2(n_435),
.B(n_436),
.Y(n_448)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_388),
.Y(n_420)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_420),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_421),
.A2(n_427),
.B1(n_412),
.B2(n_379),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_338),
.C(n_361),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_382),
.B(n_351),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_423),
.B(n_424),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_382),
.B(n_362),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_426),
.B(n_438),
.Y(n_460)
);

MAJx2_ASAP7_75t_L g428 ( 
.A(n_391),
.B(n_365),
.C(n_344),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_384),
.B(n_368),
.Y(n_429)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_429),
.Y(n_453)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_402),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_430),
.Y(n_462)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_397),
.Y(n_431)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_431),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_391),
.B(n_355),
.C(n_345),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_432),
.B(n_434),
.C(n_439),
.Y(n_459)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_397),
.Y(n_433)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_433),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_378),
.B(n_373),
.Y(n_434)
);

CKINVDCx10_ASAP7_75t_R g437 ( 
.A(n_385),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_437),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_393),
.B(n_335),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_378),
.B(n_352),
.C(n_348),
.Y(n_439)
);

A2O1A1O1Ixp25_ASAP7_75t_L g440 ( 
.A1(n_380),
.A2(n_350),
.B(n_363),
.C(n_354),
.D(n_343),
.Y(n_440)
);

NOR3xp33_ASAP7_75t_SL g467 ( 
.A(n_440),
.B(n_426),
.C(n_443),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_393),
.B(n_287),
.Y(n_441)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_441),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_384),
.B(n_356),
.Y(n_442)
);

NAND2x1_ASAP7_75t_L g443 ( 
.A(n_392),
.B(n_369),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_443),
.B(n_444),
.Y(n_457)
);

INVx13_ASAP7_75t_L g444 ( 
.A(n_385),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_445),
.B(n_447),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_387),
.B(n_296),
.C(n_367),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_446),
.B(n_406),
.C(n_403),
.Y(n_474)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_403),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_418),
.B(n_411),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_451),
.B(n_455),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_422),
.B(n_411),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_461),
.A2(n_465),
.B1(n_173),
.B2(n_157),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_463),
.A2(n_445),
.B1(n_435),
.B2(n_440),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_429),
.B(n_395),
.Y(n_464)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_464),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_425),
.A2(n_401),
.B1(n_390),
.B2(n_392),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_432),
.B(n_401),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_473),
.C(n_474),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_467),
.A2(n_470),
.B(n_189),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_419),
.A2(n_414),
.B(n_402),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_446),
.A2(n_381),
.B1(n_404),
.B2(n_410),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_471),
.A2(n_447),
.B1(n_420),
.B2(n_431),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_428),
.B(n_414),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_434),
.B(n_410),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_475),
.B(n_439),
.Y(n_478)
);

XOR2x2_ASAP7_75t_L g477 ( 
.A(n_425),
.B(n_406),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_477),
.B(n_416),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_478),
.B(n_473),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_479),
.A2(n_499),
.B1(n_500),
.B2(n_471),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_482),
.A2(n_486),
.B1(n_461),
.B2(n_458),
.Y(n_507)
);

NAND3xp33_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_442),
.C(n_433),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_483),
.B(n_487),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_456),
.B(n_443),
.C(n_416),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_484),
.B(n_485),
.C(n_494),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_456),
.B(n_459),
.C(n_455),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_448),
.A2(n_437),
.B(n_408),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_451),
.B(n_417),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_488),
.B(n_474),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_472),
.B(n_398),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_490),
.B(n_493),
.Y(n_504)
);

AND2x4_ASAP7_75t_SL g491 ( 
.A(n_457),
.B(n_409),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_491),
.B(n_492),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_457),
.B(n_409),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_462),
.B(n_398),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_459),
.B(n_444),
.C(n_340),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_452),
.Y(n_495)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_495),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_466),
.B(n_340),
.C(n_157),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_496),
.B(n_501),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_477),
.Y(n_497)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_497),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_470),
.A2(n_262),
.B(n_227),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_448),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_465),
.A2(n_173),
.B1(n_171),
.B2(n_227),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_450),
.Y(n_501)
);

A2O1A1Ixp33_ASAP7_75t_L g524 ( 
.A1(n_502),
.A2(n_468),
.B(n_449),
.C(n_476),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_453),
.B(n_464),
.Y(n_503)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_503),
.Y(n_508)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_507),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_509),
.B(n_516),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_513),
.A2(n_486),
.B1(n_492),
.B2(n_496),
.Y(n_531)
);

AOI21x1_ASAP7_75t_SL g532 ( 
.A1(n_514),
.A2(n_487),
.B(n_492),
.Y(n_532)
);

FAx1_ASAP7_75t_SL g515 ( 
.A(n_484),
.B(n_450),
.CI(n_467),
.CON(n_515),
.SN(n_515)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_518),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_488),
.B(n_460),
.Y(n_517)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_517),
.Y(n_535)
);

FAx1_ASAP7_75t_SL g518 ( 
.A(n_481),
.B(n_475),
.CI(n_458),
.CON(n_518),
.SN(n_518)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_485),
.B(n_478),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_519),
.B(n_520),
.Y(n_534)
);

FAx1_ASAP7_75t_SL g520 ( 
.A(n_481),
.B(n_463),
.CI(n_469),
.CON(n_520),
.SN(n_520)
);

INVxp33_ASAP7_75t_L g521 ( 
.A(n_498),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_521),
.B(n_491),
.Y(n_527)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_503),
.Y(n_523)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_523),
.Y(n_530)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_524),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_494),
.B(n_502),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_525),
.B(n_480),
.C(n_500),
.Y(n_536)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_527),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_508),
.B(n_489),
.Y(n_529)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_529),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_531),
.A2(n_507),
.B1(n_514),
.B2(n_506),
.Y(n_545)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_532),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_522),
.A2(n_499),
.B(n_491),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_533),
.B(n_538),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_536),
.B(n_542),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_512),
.B(n_480),
.C(n_189),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_510),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_540),
.B(n_525),
.Y(n_543)
);

AOI322xp5_ASAP7_75t_SL g541 ( 
.A1(n_504),
.A2(n_137),
.A3(n_189),
.B1(n_185),
.B2(n_171),
.C1(n_17),
.C2(n_14),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_541),
.B(n_505),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_511),
.A2(n_137),
.B(n_147),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_543),
.B(n_546),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_545),
.A2(n_530),
.B1(n_528),
.B2(n_529),
.Y(n_565)
);

FAx1_ASAP7_75t_SL g546 ( 
.A(n_526),
.B(n_515),
.CI(n_511),
.CON(n_546),
.SN(n_546)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_547),
.B(n_554),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_536),
.B(n_509),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_549),
.B(n_555),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_535),
.B(n_520),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_551),
.B(n_552),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_539),
.B(n_512),
.C(n_519),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_539),
.B(n_516),
.C(n_521),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_531),
.B(n_520),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_538),
.B(n_518),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_556),
.B(n_540),
.C(n_534),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_558),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_543),
.Y(n_560)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_560),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_556),
.A2(n_537),
.B(n_533),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_SL g571 ( 
.A(n_562),
.B(n_564),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g564 ( 
.A(n_552),
.B(n_537),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_565),
.B(n_566),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_557),
.A2(n_530),
.B(n_532),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_549),
.B(n_528),
.C(n_527),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_568),
.B(n_554),
.C(n_548),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_559),
.B(n_546),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_572),
.B(n_574),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_558),
.B(n_568),
.Y(n_574)
);

HAxp5_ASAP7_75t_SL g575 ( 
.A(n_563),
.B(n_515),
.CON(n_575),
.SN(n_575)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_575),
.A2(n_563),
.B(n_555),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_561),
.B(n_546),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_576),
.B(n_577),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_579),
.B(n_581),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_573),
.B(n_567),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_577),
.B(n_560),
.C(n_553),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_582),
.B(n_583),
.Y(n_585)
);

BUFx24_ASAP7_75t_SL g583 ( 
.A(n_571),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_580),
.B(n_573),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_586),
.A2(n_578),
.B(n_569),
.Y(n_587)
);

A2O1A1O1Ixp25_ASAP7_75t_L g589 ( 
.A1(n_587),
.A2(n_588),
.B(n_585),
.C(n_542),
.D(n_548),
.Y(n_589)
);

AOI322xp5_ASAP7_75t_L g588 ( 
.A1(n_584),
.A2(n_550),
.A3(n_575),
.B1(n_570),
.B2(n_544),
.C1(n_524),
.C2(n_518),
.Y(n_588)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_589),
.Y(n_590)
);

AOI322xp5_ASAP7_75t_SL g591 ( 
.A1(n_590),
.A2(n_12),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.C1(n_147),
.C2(n_584),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_591),
.B(n_15),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_592),
.B(n_16),
.Y(n_593)
);


endmodule