module fake_jpeg_21944_n_201 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx8_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_32),
.B1(n_20),
.B2(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_37),
.Y(n_50)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_42),
.A2(n_19),
.B1(n_24),
.B2(n_17),
.Y(n_81)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_51),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_21),
.B1(n_27),
.B2(n_26),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_39),
.B1(n_16),
.B2(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

AOI32xp33_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_36),
.A3(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_56)
);

AOI32xp33_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_92)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_59),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_39),
.B1(n_28),
.B2(n_37),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_58),
.A2(n_61),
.B1(n_80),
.B2(n_81),
.Y(n_99)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_46),
.B1(n_32),
.B2(n_20),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_17),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_67),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_37),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_71),
.B(n_76),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_72),
.A2(n_74),
.B1(n_79),
.B2(n_7),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_33),
.B1(n_23),
.B2(n_35),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_25),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_35),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_5),
.C(n_6),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_23),
.B1(n_24),
.B2(n_17),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_45),
.A2(n_25),
.B1(n_19),
.B2(n_16),
.Y(n_80)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_3),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_23),
.B(n_24),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_85),
.A2(n_91),
.B(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_78),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_62),
.B(n_1),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_81),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_3),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_98),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_7),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_102),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_6),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_104),
.B(n_72),
.Y(n_107)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_105),
.Y(n_111)
);

NAND2x1_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_77),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_106),
.A2(n_110),
.B(n_118),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_112),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_71),
.B(n_77),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_97),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_60),
.B1(n_70),
.B2(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_116),
.B(n_125),
.Y(n_128)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_96),
.B(n_75),
.Y(n_120)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_104),
.A2(n_68),
.B(n_69),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_100),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_86),
.B(n_64),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

OA21x2_ASAP7_75t_SL g125 ( 
.A1(n_91),
.A2(n_8),
.B(n_9),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_82),
.Y(n_126)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_57),
.Y(n_127)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_135),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_98),
.B(n_99),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_114),
.B(n_126),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_141),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_89),
.C(n_90),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_142),
.C(n_106),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_146),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_95),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_111),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_148),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_152),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_158),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_144),
.B(n_106),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_157),
.C(n_161),
.Y(n_168)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_108),
.Y(n_156)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_127),
.B1(n_112),
.B2(n_122),
.C(n_115),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_160),
.Y(n_164)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_118),
.C(n_119),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_153),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_166),
.B(n_167),
.Y(n_175)
);

BUFx12_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_137),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_157),
.C(n_151),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_129),
.B1(n_143),
.B2(n_145),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_155),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_172),
.B(n_140),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_165),
.Y(n_174)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_177),
.C(n_179),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_161),
.C(n_154),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_175),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_138),
.C(n_128),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_181),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_129),
.B1(n_111),
.B2(n_103),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_180),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_162),
.C(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_187),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_163),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_132),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_182),
.A2(n_163),
.B(n_169),
.Y(n_189)
);

OAI21x1_ASAP7_75t_SL g194 ( 
.A1(n_189),
.A2(n_183),
.B(n_185),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_167),
.B(n_117),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_191),
.A2(n_193),
.B(n_89),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_194),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_190),
.A2(n_192),
.B(n_95),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_196),
.C(n_105),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_198),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_116),
.Y(n_201)
);


endmodule