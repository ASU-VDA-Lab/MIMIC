module fake_jpeg_30931_n_256 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_26),
.B(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_57),
.Y(n_73)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_18),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_65),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_1),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_64),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_23),
.B1(n_39),
.B2(n_30),
.Y(n_68)
);

AO21x1_ASAP7_75t_L g133 ( 
.A1(n_68),
.A2(n_87),
.B(n_95),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_70),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_19),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_22),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_20),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_49),
.A2(n_23),
.B1(n_30),
.B2(n_17),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_43),
.A2(n_31),
.B1(n_22),
.B2(n_35),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_34),
.B1(n_25),
.B2(n_20),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_17),
.B1(n_38),
.B2(n_31),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_44),
.B(n_37),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_99),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_45),
.A2(n_17),
.B1(n_37),
.B2(n_33),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_100),
.B1(n_2),
.B2(n_3),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_44),
.B(n_35),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_55),
.A2(n_33),
.B1(n_28),
.B2(n_25),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_46),
.B(n_28),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_34),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_50),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_103),
.B(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_106),
.A2(n_95),
.B1(n_93),
.B2(n_85),
.Y(n_145)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_110),
.B(n_114),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_119),
.Y(n_135)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_17),
.B1(n_61),
.B2(n_63),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_73),
.B(n_17),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_125),
.Y(n_158)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_68),
.A2(n_59),
.B1(n_46),
.B2(n_5),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_117),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_161)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_83),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_121),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_59),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_96),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_130),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_75),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_2),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_14),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_129),
.Y(n_144)
);

AOI32xp33_ASAP7_75t_L g129 ( 
.A1(n_87),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_129)
);

AOI32xp33_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_104),
.A3(n_107),
.B1(n_112),
.B2(n_115),
.Y(n_149)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_6),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_96),
.C(n_78),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_82),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_132),
.A2(n_85),
.B1(n_93),
.B2(n_71),
.Y(n_159)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_140),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_124),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_149),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_157),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_118),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_10),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_151),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_125),
.A2(n_92),
.B1(n_79),
.B2(n_78),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_161),
.B1(n_131),
.B2(n_119),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_92),
.B1(n_79),
.B2(n_75),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_159),
.A2(n_117),
.B(n_133),
.Y(n_165)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_103),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_166),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_165),
.A2(n_171),
.B1(n_180),
.B2(n_160),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_133),
.B(n_123),
.C(n_114),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_158),
.B(n_103),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_176),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_154),
.B(n_127),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_169),
.B(n_135),
.Y(n_185)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_170),
.B(n_179),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_158),
.A2(n_133),
.B(n_105),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_172),
.A2(n_143),
.B(n_145),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_150),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_173),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_109),
.C(n_108),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_137),
.C(n_142),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_116),
.B1(n_126),
.B2(n_134),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_181),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_157),
.B1(n_152),
.B2(n_147),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_152),
.A2(n_147),
.B1(n_161),
.B2(n_140),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_110),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_183),
.Y(n_188)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_11),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_162),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_185),
.B(n_187),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_195),
.C(n_177),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_181),
.A2(n_137),
.B(n_156),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_190),
.B(n_192),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_153),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_198),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_156),
.C(n_153),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_184),
.B(n_155),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_197),
.B(n_168),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_130),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_176),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_200),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_130),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_202),
.B(n_172),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_203),
.A2(n_168),
.B1(n_179),
.B2(n_171),
.Y(n_207)
);

AO221x1_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_201),
.B1(n_186),
.B2(n_163),
.C(n_170),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_204),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_196),
.A2(n_168),
.B1(n_166),
.B2(n_165),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_205),
.A2(n_207),
.B1(n_218),
.B2(n_191),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_209),
.B(n_216),
.Y(n_229)
);

AO221x1_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_183),
.B1(n_182),
.B2(n_173),
.C(n_150),
.Y(n_211)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_189),
.C(n_214),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_167),
.Y(n_213)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_174),
.Y(n_214)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g222 ( 
.A(n_217),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_196),
.A2(n_191),
.B1(n_187),
.B2(n_195),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_226),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_225),
.C(n_208),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_193),
.C(n_185),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_193),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_197),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_209),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_234),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_210),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_233),
.C(n_236),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_216),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_229),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_235),
.A2(n_237),
.B(n_204),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_215),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_228),
.A2(n_208),
.B(n_217),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_235),
.A2(n_219),
.B1(n_205),
.B2(n_227),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_239),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_230),
.A2(n_222),
.B1(n_207),
.B2(n_221),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_220),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_242),
.B(n_243),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_230),
.A2(n_224),
.B1(n_186),
.B2(n_234),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_213),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_247),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_211),
.C(n_160),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_240),
.A2(n_11),
.B(n_12),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_13),
.B(n_238),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_252),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_242),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_250),
.A2(n_249),
.B(n_241),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_253),
.B(n_241),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_254),
.Y(n_256)
);


endmodule