module fake_aes_238_n_23 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_23);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_23;
wire n_20;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
AND2x4_ASAP7_75t_L g9 ( .A(n_0), .B(n_6), .Y(n_9) );
BUFx3_ASAP7_75t_L g10 ( .A(n_3), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
BUFx2_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_1), .B(n_4), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
AOI21x1_ASAP7_75t_L g15 ( .A1(n_11), .A2(n_7), .B(n_8), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_12), .Y(n_16) );
OAI21x1_ASAP7_75t_SL g17 ( .A1(n_11), .A2(n_1), .B(n_3), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_16), .B(n_10), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_15), .B(n_9), .Y(n_19) );
OAI21xp5_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_15), .B(n_9), .Y(n_20) );
AO22x2_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_17), .B1(n_18), .B2(n_13), .Y(n_21) );
OA22x2_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_13), .B1(n_14), .B2(n_5), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
endmodule