module fake_jpeg_28143_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g16 ( 
.A(n_10),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_38),
.Y(n_46)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_47),
.B(n_62),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_26),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_65),
.Y(n_73)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_40),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_74),
.B(n_31),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_30),
.B1(n_19),
.B2(n_26),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_51),
.A2(n_30),
.B1(n_17),
.B2(n_16),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_71),
.B1(n_45),
.B2(n_68),
.Y(n_100)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_30),
.B1(n_17),
.B2(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_75),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_77),
.B(n_78),
.Y(n_108)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_83),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_50),
.B(n_57),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_39),
.C(n_44),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_45),
.B1(n_35),
.B2(n_17),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_81),
.A2(n_87),
.B1(n_63),
.B2(n_37),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_50),
.B(n_22),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_27),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_89),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_54),
.A2(n_45),
.B1(n_43),
.B2(n_41),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_21),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_42),
.Y(n_97)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_73),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_96),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_112),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_73),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_99),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_118),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_102),
.B(n_23),
.Y(n_151)
);

AO21x1_ASAP7_75t_L g144 ( 
.A1(n_104),
.A2(n_114),
.B(n_34),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_34),
.B(n_31),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_31),
.B(n_34),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_44),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_120),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_43),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_22),
.Y(n_146)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_44),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_115),
.B(n_123),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_74),
.A2(n_63),
.B1(n_27),
.B2(n_37),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_20),
.B1(n_82),
.B2(n_85),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_124),
.B1(n_81),
.B2(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_44),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_66),
.A2(n_37),
.B1(n_44),
.B2(n_42),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_130),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_84),
.B(n_80),
.C(n_77),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_129),
.A2(n_136),
.B(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_120),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_131),
.B(n_133),
.Y(n_186)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_145),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_88),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_115),
.B(n_86),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_134),
.B(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_78),
.C(n_70),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_105),
.C(n_103),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_138),
.A2(n_121),
.B1(n_101),
.B2(n_106),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_112),
.A2(n_116),
.B1(n_109),
.B2(n_104),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_105),
.B1(n_103),
.B2(n_85),
.Y(n_171)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_22),
.A3(n_23),
.B1(n_75),
.B2(n_72),
.Y(n_140)
);

AOI32xp33_ASAP7_75t_L g174 ( 
.A1(n_140),
.A2(n_24),
.A3(n_28),
.B1(n_33),
.B2(n_18),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_79),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_141),
.B(n_142),
.Y(n_163)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp33_ASAP7_75t_SL g155 ( 
.A(n_144),
.B(n_102),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_SL g145 ( 
.A(n_107),
.B(n_42),
.C(n_44),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_146),
.B(n_18),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_113),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_151),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_82),
.Y(n_149)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_33),
.Y(n_153)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

AO22x1_ASAP7_75t_L g202 ( 
.A1(n_155),
.A2(n_174),
.B1(n_144),
.B2(n_135),
.Y(n_202)
);

AOI22x1_ASAP7_75t_SL g157 ( 
.A1(n_152),
.A2(n_100),
.B1(n_114),
.B2(n_99),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_157),
.A2(n_171),
.B(n_182),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_146),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_158),
.B(n_166),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_162),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_97),
.Y(n_166)
);

AO22x1_ASAP7_75t_SL g167 ( 
.A1(n_154),
.A2(n_114),
.B1(n_97),
.B2(n_121),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_76),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_188),
.C(n_136),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_177),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_141),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_173),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_129),
.A2(n_23),
.B(n_20),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_151),
.B(n_143),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_178),
.B1(n_180),
.B2(n_127),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_139),
.B(n_18),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_142),
.A2(n_106),
.B1(n_92),
.B2(n_49),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_126),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_181),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_138),
.A2(n_61),
.B1(n_49),
.B2(n_93),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_0),
.B(n_1),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_125),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_18),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_93),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_125),
.B(n_39),
.C(n_61),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_169),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_193),
.Y(n_230)
);

OA22x2_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_143),
.B1(n_126),
.B2(n_140),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_202),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_147),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_130),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_194),
.A2(n_212),
.B(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_201),
.Y(n_240)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_207),
.C(n_188),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_148),
.B1(n_93),
.B2(n_76),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_160),
.B1(n_162),
.B2(n_171),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_159),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_208),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_39),
.C(n_76),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_213),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_217),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_164),
.B(n_33),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_33),
.Y(n_214)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_158),
.B(n_183),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_215),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_25),
.B(n_1),
.Y(n_216)
);

A2O1A1O1Ixp25_ASAP7_75t_L g217 ( 
.A1(n_181),
.A2(n_18),
.B(n_25),
.C(n_28),
.D(n_8),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_187),
.B(n_7),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_218),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_166),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_223),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_222),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_177),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_231),
.C(n_232),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_206),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_235),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_194),
.A2(n_180),
.B1(n_184),
.B2(n_170),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_227),
.B(n_196),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_167),
.C(n_185),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_167),
.C(n_172),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_182),
.C(n_175),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_190),
.C(n_216),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_199),
.Y(n_235)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_241),
.Y(n_264)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_244),
.B(n_258),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_250),
.Y(n_266)
);

NOR3xp33_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_204),
.C(n_217),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_252),
.Y(n_278)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_254),
.Y(n_274)
);

BUFx24_ASAP7_75t_SL g252 ( 
.A(n_228),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_223),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_212),
.C(n_189),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_260),
.C(n_219),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_220),
.A2(n_194),
.B1(n_202),
.B2(n_192),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_261),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_201),
.C(n_192),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_224),
.A2(n_192),
.B1(n_28),
.B2(n_8),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_243),
.A2(n_28),
.B1(n_8),
.B2(n_9),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_5),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_263),
.A2(n_236),
.B(n_238),
.Y(n_265)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_221),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_267),
.B(n_270),
.Y(n_285)
);

BUFx12_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_268),
.B(n_269),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_257),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_232),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_279),
.Y(n_286)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_264),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_273),
.B(n_275),
.Y(n_295)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_246),
.A2(n_237),
.B1(n_239),
.B2(n_234),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_263),
.B1(n_253),
.B2(n_249),
.Y(n_284)
);

AO22x1_ASAP7_75t_L g277 ( 
.A1(n_245),
.A2(n_219),
.B1(n_222),
.B2(n_2),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

INVx11_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_294),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_280),
.A2(n_255),
.B1(n_260),
.B2(n_253),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_283),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_11),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_265),
.A2(n_5),
.B(n_13),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_287),
.A2(n_289),
.B(n_11),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_6),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_272),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_6),
.C(n_13),
.Y(n_292)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_274),
.A2(n_15),
.B(n_13),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_12),
.Y(n_307)
);

OA21x2_ASAP7_75t_SL g297 ( 
.A1(n_295),
.A2(n_288),
.B(n_291),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_297),
.A2(n_305),
.B(n_3),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_290),
.A2(n_281),
.B(n_271),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_298),
.A2(n_300),
.B(n_304),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_280),
.B(n_270),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_306),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_277),
.B1(n_268),
.B2(n_11),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_307),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_267),
.B(n_15),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_282),
.B(n_292),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_285),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_299),
.B(n_285),
.Y(n_309)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_317),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_314),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_0),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_316),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_2),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_3),
.Y(n_320)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

AOI21x1_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_3),
.B(n_4),
.Y(n_323)
);

OA21x2_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_312),
.B(n_310),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_324),
.B(n_325),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_313),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_321),
.C(n_322),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_328),
.A2(n_326),
.B1(n_314),
.B2(n_318),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_3),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_4),
.Y(n_331)
);


endmodule