module fake_jpeg_26786_n_181 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_181);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_57),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_24),
.B1(n_19),
.B2(n_20),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_51),
.B1(n_43),
.B2(n_38),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_50),
.B(n_16),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_24),
.B1(n_30),
.B2(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_18),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_21),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_21),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_32),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_69),
.Y(n_91)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_62),
.Y(n_93)
);

OR2x2_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_31),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_67),
.B(n_74),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_30),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_81),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_22),
.B(n_15),
.C(n_29),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_77),
.B1(n_47),
.B2(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_71),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_25),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_22),
.B(n_15),
.C(n_29),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_34),
.B1(n_24),
.B2(n_43),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_47),
.B1(n_57),
.B2(n_34),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_36),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_38),
.C(n_36),
.Y(n_96)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_23),
.B(n_27),
.C(n_31),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_0),
.B(n_1),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_33),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_85),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_33),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_25),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_78),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_104),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_34),
.B1(n_38),
.B2(n_36),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_99),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_42),
.B1(n_27),
.B2(n_23),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_67),
.B(n_85),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_37),
.C(n_42),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_37),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_105),
.B(n_73),
.Y(n_118)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_109),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_63),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_70),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_102),
.B1(n_68),
.B2(n_79),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_113),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_103),
.A2(n_81),
.B(n_84),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_117),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_115),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_84),
.B(n_80),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_121),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_69),
.B1(n_74),
.B2(n_64),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_123),
.B1(n_91),
.B2(n_92),
.Y(n_128)
);

OA21x2_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_89),
.B(n_105),
.Y(n_120)
);

OAI321xp33_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_97),
.A3(n_94),
.B1(n_102),
.B2(n_42),
.C(n_37),
.Y(n_135)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_94),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_108),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_124),
.A2(n_98),
.B1(n_96),
.B2(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_131),
.B(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_122),
.B1(n_121),
.B2(n_115),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_136),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_106),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_122),
.B1(n_119),
.B2(n_93),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_140),
.A2(n_151),
.B1(n_1),
.B2(n_2),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_116),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_150),
.C(n_139),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_145),
.Y(n_157)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_149),
.B1(n_62),
.B2(n_2),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_120),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_114),
.B1(n_112),
.B2(n_117),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_134),
.C(n_127),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_155),
.C(n_158),
.Y(n_162)
);

AOI322xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_134),
.A3(n_139),
.B1(n_135),
.B2(n_129),
.C1(n_123),
.C2(n_137),
.Y(n_153)
);

OAI31xp33_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_13),
.A3(n_11),
.B(n_10),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_14),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_93),
.C(n_37),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_37),
.C(n_75),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_160),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_144),
.B(n_148),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_164),
.Y(n_170)
);

OAI21x1_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_142),
.B(n_9),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_9),
.Y(n_165)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_3),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_167),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_152),
.B1(n_4),
.B2(n_5),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_162),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_172),
.C(n_7),
.Y(n_175)
);

AOI21x1_ASAP7_75t_L g173 ( 
.A1(n_170),
.A2(n_162),
.B(n_166),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_175),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_176),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_169),
.A2(n_4),
.B(n_6),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_171),
.B(n_168),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_178),
.C(n_172),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_7),
.Y(n_181)
);


endmodule