module fake_jpeg_12493_n_520 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_520);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_520;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_8),
.B(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_60),
.Y(n_171)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_63),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_64),
.B(n_77),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_16),
.C(n_15),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_65),
.B(n_27),
.C(n_39),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_66),
.Y(n_170)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_67),
.Y(n_186)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g168 ( 
.A(n_68),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_25),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_69),
.B(n_70),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_25),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_71),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_75),
.Y(n_127)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_16),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_78),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_14),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_79),
.B(n_98),
.Y(n_176)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_82),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_83),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_84),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_28),
.B(n_0),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_85),
.B(n_106),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_40),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_92),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_87),
.Y(n_204)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_88),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_19),
.Y(n_89)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_90),
.Y(n_199)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g192 ( 
.A(n_91),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_22),
.Y(n_92)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_93),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_97),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_30),
.B(n_13),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_40),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_105),
.Y(n_148)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_103),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_30),
.B(n_13),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_32),
.B(n_0),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_32),
.B(n_1),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_108),
.B(n_113),
.Y(n_161)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_22),
.Y(n_109)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_23),
.Y(n_110)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_20),
.Y(n_112)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_36),
.B(n_1),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_22),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_115),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_40),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_40),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_116),
.B(n_119),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_23),
.Y(n_117)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_41),
.B(n_1),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_118),
.B(n_2),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_41),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_54),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_120),
.B(n_125),
.Y(n_183)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_20),
.Y(n_121)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_44),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_85),
.A2(n_24),
.B1(n_58),
.B2(n_53),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_130),
.A2(n_147),
.B1(n_163),
.B2(n_175),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_84),
.A2(n_53),
.B1(n_58),
.B2(n_24),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_134),
.A2(n_149),
.B1(n_154),
.B2(n_158),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_113),
.A2(n_58),
.B1(n_24),
.B2(n_27),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_67),
.A2(n_50),
.B1(n_45),
.B2(n_38),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_150),
.B(n_138),
.C(n_140),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_73),
.A2(n_21),
.B1(n_50),
.B2(n_45),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_78),
.A2(n_38),
.B1(n_37),
.B2(n_31),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g162 ( 
.A1(n_82),
.A2(n_52),
.B(n_39),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_162),
.B(n_189),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_96),
.A2(n_37),
.B1(n_31),
.B2(n_21),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_60),
.A2(n_52),
.B1(n_35),
.B2(n_4),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_164),
.A2(n_167),
.B1(n_178),
.B2(n_188),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_61),
.A2(n_35),
.B1(n_3),
.B2(n_4),
.Y(n_167)
);

HAxp5_ASAP7_75t_SL g169 ( 
.A(n_68),
.B(n_2),
.CON(n_169),
.SN(n_169)
);

AOI21xp33_ASAP7_75t_L g213 ( 
.A1(n_169),
.A2(n_80),
.B(n_66),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_65),
.A2(n_110),
.B1(n_100),
.B2(n_76),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_62),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_187),
.B(n_193),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_72),
.A2(n_90),
.B1(n_97),
.B2(n_89),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_120),
.B(n_7),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_122),
.B(n_7),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_191),
.B(n_195),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_124),
.B(n_9),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_114),
.B(n_9),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_114),
.B(n_9),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_196),
.B(n_201),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_72),
.A2(n_9),
.B1(n_10),
.B2(n_107),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_197),
.A2(n_208),
.B1(n_131),
.B2(n_181),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_81),
.B(n_10),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_103),
.B(n_10),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_202),
.B(n_203),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_75),
.B(n_88),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_117),
.B(n_109),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_209),
.Y(n_232)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_63),
.Y(n_207)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_93),
.A2(n_91),
.B1(n_71),
.B2(n_94),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_111),
.B(n_123),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_129),
.B(n_80),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_210),
.Y(n_330)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_211),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_174),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_212),
.B(n_228),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_213),
.B(n_220),
.Y(n_291)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_214),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_161),
.B(n_83),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_216),
.B(n_223),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_217),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_218),
.Y(n_327)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_219),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_172),
.B(n_146),
.Y(n_220)
);

INVx6_ASAP7_75t_SL g221 ( 
.A(n_168),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_221),
.Y(n_316)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_222),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_157),
.B(n_87),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_135),
.Y(n_224)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_224),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_177),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_226),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_134),
.A2(n_95),
.B1(n_101),
.B2(n_102),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_227),
.A2(n_251),
.B1(n_263),
.B2(n_256),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_180),
.B(n_104),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_169),
.A2(n_155),
.B1(n_133),
.B2(n_132),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_229),
.A2(n_238),
.B1(n_244),
.B2(n_259),
.Y(n_311)
);

AOI21xp33_ASAP7_75t_L g231 ( 
.A1(n_176),
.A2(n_148),
.B(n_151),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_231),
.Y(n_333)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_177),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_233),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_185),
.A2(n_160),
.B(n_136),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_234),
.A2(n_276),
.B(n_210),
.Y(n_308)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_128),
.Y(n_235)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_127),
.Y(n_236)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_236),
.Y(n_313)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_237),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_163),
.A2(n_141),
.B1(n_179),
.B2(n_173),
.Y(n_238)
);

AND2x2_ASAP7_75t_SL g239 ( 
.A(n_139),
.B(n_194),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_239),
.B(n_240),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g240 ( 
.A(n_156),
.B(n_171),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_126),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_241),
.B(n_261),
.Y(n_289)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_242),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_183),
.A2(n_165),
.B(n_149),
.C(n_158),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_243),
.A2(n_228),
.B(n_240),
.C(n_220),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_133),
.A2(n_155),
.B1(n_132),
.B2(n_171),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_L g247 ( 
.A1(n_154),
.A2(n_197),
.B(n_188),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_247),
.B(n_249),
.Y(n_300)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_152),
.Y(n_248)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_248),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_199),
.B(n_145),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_250),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_208),
.A2(n_164),
.B1(n_167),
.B2(n_153),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_145),
.B(n_127),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_252),
.B(n_277),
.Y(n_314)
);

AO22x1_ASAP7_75t_L g254 ( 
.A1(n_182),
.A2(n_144),
.B1(n_173),
.B2(n_159),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_254),
.A2(n_249),
.B(n_271),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_153),
.B(n_179),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_257),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_144),
.B(n_159),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_143),
.Y(n_258)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_258),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_192),
.A2(n_140),
.B1(n_186),
.B2(n_182),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_184),
.Y(n_260)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_260),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_137),
.B(n_131),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_143),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_264),
.B(n_266),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_204),
.B(n_166),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_269),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_137),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_142),
.Y(n_267)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_267),
.Y(n_299)
);

BUFx12f_ASAP7_75t_L g268 ( 
.A(n_186),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_268),
.B(n_271),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_204),
.B(n_142),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_240),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_181),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_137),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_279),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_166),
.B(n_200),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_275),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_200),
.B(n_143),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_205),
.A2(n_84),
.B1(n_34),
.B2(n_73),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_205),
.B(n_157),
.C(n_161),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_128),
.Y(n_278)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_278),
.Y(n_305)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_128),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_174),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_234),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_215),
.A2(n_252),
.B(n_243),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_283),
.A2(n_308),
.B(n_318),
.Y(n_343)
);

O2A1O1Ixp33_ASAP7_75t_L g285 ( 
.A1(n_239),
.A2(n_247),
.B(n_246),
.C(n_221),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_285),
.A2(n_317),
.B(n_329),
.Y(n_345)
);

OA22x2_ASAP7_75t_L g369 ( 
.A1(n_286),
.A2(n_298),
.B1(n_316),
.B2(n_297),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_227),
.A2(n_251),
.B1(n_273),
.B2(n_232),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_273),
.A2(n_223),
.B1(n_216),
.B2(n_270),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_303),
.A2(n_242),
.B1(n_233),
.B2(n_214),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_304),
.B(n_314),
.C(n_283),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_253),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_312),
.B(n_319),
.Y(n_353)
);

O2A1O1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_239),
.A2(n_210),
.B(n_249),
.C(n_220),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_225),
.B(n_255),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_321),
.B(n_332),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_319),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_274),
.A2(n_269),
.B1(n_265),
.B2(n_245),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_325),
.A2(n_331),
.B1(n_329),
.B2(n_282),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_257),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_217),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_240),
.A2(n_254),
.B(n_275),
.C(n_230),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_262),
.A2(n_237),
.B1(n_224),
.B2(n_250),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_211),
.B(n_260),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_300),
.A2(n_254),
.B1(n_258),
.B2(n_268),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_335),
.A2(n_306),
.B(n_324),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_336),
.B(n_339),
.Y(n_380)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_327),
.Y(n_337)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_337),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_290),
.Y(n_338)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_338),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_281),
.B(n_219),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_340),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_310),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_341),
.B(n_342),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_332),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_332),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_344),
.B(n_347),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_314),
.B(n_222),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_346),
.B(n_356),
.C(n_364),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_333),
.B(n_217),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_299),
.Y(n_348)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_312),
.B(n_268),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_349),
.B(n_351),
.Y(n_390)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_299),
.Y(n_350)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_350),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_289),
.B(n_218),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_360),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_325),
.A2(n_285),
.B1(n_300),
.B2(n_291),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_354),
.A2(n_359),
.B1(n_371),
.B2(n_290),
.Y(n_387)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_290),
.Y(n_355)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_355),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_286),
.A2(n_303),
.B1(n_282),
.B2(n_292),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_357),
.A2(n_361),
.B1(n_362),
.B2(n_366),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_358),
.B(n_368),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_300),
.A2(n_291),
.B1(n_304),
.B2(n_292),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_307),
.B(n_293),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_293),
.A2(n_307),
.B1(n_318),
.B2(n_291),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_308),
.A2(n_304),
.B1(n_330),
.B2(n_311),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_294),
.B(n_331),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_363),
.B(n_365),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_294),
.C(n_295),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_294),
.B(n_305),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_317),
.A2(n_321),
.B1(n_305),
.B2(n_297),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_309),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_369),
.B(n_373),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_296),
.B(n_301),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_370),
.B(n_374),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_320),
.A2(n_315),
.B1(n_334),
.B2(n_322),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_302),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_372),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_313),
.B(n_287),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_302),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_287),
.B(n_288),
.Y(n_375)
);

AND2x2_ASAP7_75t_SL g391 ( 
.A(n_375),
.B(n_326),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_352),
.A2(n_322),
.B1(n_315),
.B2(n_327),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_377),
.B(n_395),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_343),
.A2(n_345),
.B(n_362),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_378),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_375),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_387),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_392),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_339),
.A2(n_288),
.B1(n_284),
.B2(n_306),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_389),
.A2(n_401),
.B1(n_407),
.B2(n_369),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_391),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_345),
.A2(n_284),
.B(n_326),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_354),
.A2(n_359),
.B1(n_360),
.B2(n_353),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_373),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_356),
.B(n_346),
.C(n_353),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_398),
.B(n_367),
.C(n_369),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_357),
.A2(n_366),
.B1(n_363),
.B2(n_361),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_369),
.A2(n_358),
.B1(n_349),
.B2(n_335),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_406),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_371),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_369),
.A2(n_367),
.B1(n_342),
.B2(n_344),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_403),
.Y(n_409)
);

AO32x1_ASAP7_75t_L g410 ( 
.A1(n_381),
.A2(n_343),
.A3(n_367),
.B1(n_365),
.B2(n_364),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_410),
.A2(n_383),
.B(n_400),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_412),
.A2(n_418),
.B1(n_419),
.B2(n_377),
.Y(n_446)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_404),
.Y(n_414)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_414),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_421),
.C(n_422),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_406),
.A2(n_408),
.B1(n_379),
.B2(n_384),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_416),
.A2(n_388),
.B(n_380),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_401),
.A2(n_350),
.B1(n_368),
.B2(n_337),
.Y(n_418)
);

OAI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_407),
.A2(n_393),
.B1(n_396),
.B2(n_402),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_376),
.B(n_372),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_376),
.B(n_374),
.C(n_355),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_405),
.Y(n_423)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_423),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_337),
.Y(n_424)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_424),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_376),
.B(n_398),
.C(n_395),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_425),
.B(n_398),
.C(n_393),
.Y(n_438)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_394),
.Y(n_427)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_427),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_385),
.B(n_386),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_428),
.Y(n_444)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_384),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_396),
.B(n_381),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_431),
.B(n_386),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_435),
.B(n_445),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_440),
.C(n_441),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_439),
.B(n_451),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_425),
.B(n_378),
.C(n_383),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_421),
.B(n_400),
.C(n_387),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_429),
.A2(n_420),
.B1(n_417),
.B2(n_408),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_442),
.B(n_417),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_390),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_443),
.B(n_447),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_415),
.B(n_382),
.C(n_392),
.Y(n_445)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_446),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_410),
.B(n_390),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_448),
.A2(n_449),
.B(n_450),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_426),
.A2(n_380),
.B(n_382),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_426),
.A2(n_391),
.B1(n_405),
.B2(n_399),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_428),
.B(n_391),
.Y(n_451)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_452),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_444),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_454),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_440),
.B(n_420),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_459),
.B(n_441),
.Y(n_473)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_437),
.Y(n_460)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_460),
.Y(n_479)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_432),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_461),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_448),
.A2(n_411),
.B(n_413),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_462),
.A2(n_467),
.B(n_411),
.Y(n_475)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_432),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_463),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_433),
.B(n_424),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_464),
.B(n_466),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_433),
.B(n_418),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_449),
.A2(n_411),
.B(n_413),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_438),
.C(n_436),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_469),
.B(n_470),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_436),
.C(n_443),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_473),
.B(n_478),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_475),
.A2(n_462),
.B(n_457),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_455),
.B(n_445),
.C(n_447),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_480),
.C(n_459),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_435),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_455),
.B(n_450),
.C(n_451),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_471),
.A2(n_453),
.B1(n_429),
.B2(n_454),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_481),
.A2(n_474),
.B1(n_468),
.B2(n_479),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_473),
.B(n_465),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_485),
.Y(n_496)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_472),
.Y(n_484)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_484),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_486),
.B(n_489),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_480),
.B(n_457),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_491),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_471),
.A2(n_434),
.B1(n_466),
.B2(n_475),
.Y(n_488)
);

OA21x2_ASAP7_75t_L g489 ( 
.A1(n_478),
.A2(n_442),
.B(n_434),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_470),
.B(n_456),
.Y(n_491)
);

BUFx24_ASAP7_75t_SL g492 ( 
.A(n_482),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_499),
.Y(n_505)
);

FAx1_ASAP7_75t_SL g495 ( 
.A(n_485),
.B(n_477),
.CI(n_469),
.CON(n_495),
.SN(n_495)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_497),
.Y(n_506)
);

FAx1_ASAP7_75t_SL g497 ( 
.A(n_486),
.B(n_456),
.CI(n_464),
.CON(n_497),
.SN(n_497)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_498),
.A2(n_488),
.B1(n_489),
.B2(n_479),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_476),
.C(n_474),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_476),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_501),
.B(n_500),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_496),
.B(n_491),
.C(n_490),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_502),
.B(n_503),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_500),
.B(n_490),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_504),
.B(n_507),
.C(n_508),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_499),
.B(n_489),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_506),
.A2(n_495),
.B(n_494),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_511),
.A2(n_512),
.B(n_513),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_505),
.B(n_501),
.C(n_493),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_506),
.A2(n_493),
.B(n_497),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_509),
.B(n_503),
.Y(n_515)
);

AO21x1_ASAP7_75t_L g516 ( 
.A1(n_515),
.A2(n_502),
.B(n_481),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_514),
.C(n_510),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_517),
.B(n_430),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_518),
.B(n_414),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_519),
.B(n_409),
.Y(n_520)
);


endmodule