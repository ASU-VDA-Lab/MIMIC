module fake_ibex_1464_n_929 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_929);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_929;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_510;
wire n_193;
wire n_418;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_798;
wire n_732;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_543;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_817;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_288;
wire n_247;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_298;
wire n_231;
wire n_202;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

INVxp33_ASAP7_75t_SL g163 ( 
.A(n_81),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_70),
.Y(n_164)
);

NOR2xp67_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_151),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_6),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_53),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_18),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_49),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_84),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_114),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_16),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_102),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_38),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_66),
.Y(n_178)
);

NOR2xp67_ASAP7_75t_L g179 ( 
.A(n_93),
.B(n_2),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_27),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

BUFx2_ASAP7_75t_SL g184 ( 
.A(n_107),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_15),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_17),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_50),
.B(n_74),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_101),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_69),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_32),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_10),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_51),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_23),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_25),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_139),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_55),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_133),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_33),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_37),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_129),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_137),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_128),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_16),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_92),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_144),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_87),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_97),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_18),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_135),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_32),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_109),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_82),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_123),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_64),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_149),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_54),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_140),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_117),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_150),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_111),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_13),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_71),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_99),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_13),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_112),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_119),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_79),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_75),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_44),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_24),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_121),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_59),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_138),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_100),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_85),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_56),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_131),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_21),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_10),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_7),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_24),
.Y(n_241)
);

INVx4_ASAP7_75t_R g242 ( 
.A(n_22),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_26),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_41),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_147),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_90),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_143),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_96),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_94),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_80),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_47),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_52),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_33),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_7),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_22),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_39),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_45),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_152),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_34),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_125),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_115),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_136),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_155),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_124),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_108),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_68),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_110),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_25),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_88),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_89),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_113),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_130),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_14),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_158),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_46),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_120),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_175),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_277)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_275),
.A2(n_83),
.B(n_159),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_240),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_189),
.B(n_0),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_195),
.Y(n_281)
);

OAI21x1_ASAP7_75t_L g282 ( 
.A1(n_275),
.A2(n_86),
.B(n_157),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_181),
.Y(n_283)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_189),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_175),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_240),
.B(n_1),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_167),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_185),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_181),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_189),
.B(n_3),
.Y(n_292)
);

AND2x4_ASAP7_75t_L g293 ( 
.A(n_211),
.B(n_4),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_162),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_207),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_183),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_171),
.Y(n_297)
);

AND2x2_ASAP7_75t_SL g298 ( 
.A(n_166),
.B(n_40),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_207),
.B(n_4),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_5),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_183),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_169),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_271),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_186),
.B(n_6),
.Y(n_305)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_195),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_193),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_170),
.B(n_8),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_180),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_172),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_173),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_190),
.Y(n_312)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_195),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_194),
.B(n_8),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_195),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_182),
.Y(n_316)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_201),
.A2(n_91),
.B(n_156),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_201),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_193),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_196),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_193),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_227),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_205),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_191),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_205),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_232),
.Y(n_326)
);

AND2x4_ASAP7_75t_L g327 ( 
.A(n_232),
.B(n_9),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_198),
.B(n_11),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_178),
.A2(n_12),
.B1(n_14),
.B2(n_17),
.Y(n_329)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_205),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_246),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_197),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_209),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_256),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_193),
.Y(n_335)
);

OAI21x1_ASAP7_75t_L g336 ( 
.A1(n_256),
.A2(n_95),
.B(n_154),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_261),
.Y(n_337)
);

AND2x4_ASAP7_75t_L g338 ( 
.A(n_261),
.B(n_19),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_208),
.B(n_19),
.Y(n_339)
);

OAI22x1_ASAP7_75t_L g340 ( 
.A1(n_203),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_199),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_206),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_210),
.B(n_20),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_212),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_213),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_214),
.Y(n_346)
);

OA21x2_ASAP7_75t_L g347 ( 
.A1(n_215),
.A2(n_98),
.B(n_153),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_216),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_209),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_217),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_293),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_281),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_327),
.B(n_218),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_284),
.B(n_224),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_327),
.Y(n_355)
);

CKINVDCx6p67_ASAP7_75t_R g356 ( 
.A(n_298),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_327),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_281),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_281),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_338),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_281),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_284),
.B(n_279),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_338),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_338),
.B(n_222),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_315),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_284),
.B(n_230),
.Y(n_366)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_286),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_302),
.Y(n_368)
);

OR2x6_ASAP7_75t_L g369 ( 
.A(n_277),
.B(n_184),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_284),
.B(n_188),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g371 ( 
.A(n_302),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_315),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_315),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_293),
.B(n_223),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_315),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_286),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_279),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_309),
.B(n_238),
.Y(n_378)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_304),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_309),
.B(n_241),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_315),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_285),
.B(n_178),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_341),
.B(n_254),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_323),
.Y(n_384)
);

BUFx6f_ASAP7_75t_SL g385 ( 
.A(n_298),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_341),
.B(n_255),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_303),
.A2(n_292),
.B1(n_280),
.B2(n_324),
.Y(n_387)
);

OR2x6_ASAP7_75t_L g388 ( 
.A(n_280),
.B(n_221),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_323),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_294),
.B(n_226),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_323),
.Y(n_391)
);

INVx8_ASAP7_75t_L g392 ( 
.A(n_299),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_310),
.B(n_228),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_299),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_323),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_304),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_300),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_326),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_310),
.B(n_231),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_311),
.B(n_233),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_311),
.B(n_316),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_325),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_348),
.B(n_259),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_300),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_283),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_305),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_325),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_283),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_304),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_320),
.B(n_273),
.Y(n_411)
);

AO21x2_ASAP7_75t_L g412 ( 
.A1(n_317),
.A2(n_236),
.B(n_234),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_332),
.B(n_244),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_325),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_331),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_332),
.B(n_245),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_292),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_325),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_289),
.B(n_239),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_297),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_285),
.Y(n_421)
);

INVx5_ASAP7_75t_L g422 ( 
.A(n_306),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_291),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_290),
.B(n_253),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_296),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_301),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_297),
.Y(n_427)
);

NOR2x1p5_ASAP7_75t_L g428 ( 
.A(n_312),
.B(n_276),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_301),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_318),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_L g431 ( 
.A(n_350),
.B(n_209),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_339),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_333),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_333),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_333),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_333),
.Y(n_436)
);

BUFx4f_ASAP7_75t_L g437 ( 
.A(n_346),
.Y(n_437)
);

OR2x6_ASAP7_75t_L g438 ( 
.A(n_340),
.B(n_179),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_SL g439 ( 
.A(n_340),
.B(n_200),
.Y(n_439)
);

BUFx10_ASAP7_75t_L g440 ( 
.A(n_295),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_346),
.B(n_168),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_330),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_333),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_322),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_322),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_350),
.Y(n_446)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_330),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_334),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_334),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_342),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_349),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_349),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_337),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_349),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_339),
.Y(n_455)
);

BUFx6f_ASAP7_75t_SL g456 ( 
.A(n_288),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_349),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_349),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_342),
.B(n_250),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_344),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_398),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_354),
.B(n_345),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_437),
.B(n_163),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_405),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_L g465 ( 
.A1(n_360),
.A2(n_345),
.B1(n_343),
.B2(n_314),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_408),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_446),
.B(n_362),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_360),
.A2(n_328),
.B1(n_308),
.B2(n_287),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_362),
.B(n_287),
.Y(n_469)
);

AND2x6_ASAP7_75t_L g470 ( 
.A(n_351),
.B(n_251),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_371),
.B(n_200),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_408),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_425),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_368),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_437),
.B(n_174),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_367),
.B(n_176),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_392),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_371),
.B(n_202),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_367),
.B(n_177),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_378),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_385),
.B(n_202),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_430),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_366),
.B(n_252),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_410),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_428),
.B(n_329),
.Y(n_485)
);

INVx8_ASAP7_75t_L g486 ( 
.A(n_392),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_392),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_394),
.B(n_258),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_367),
.B(n_278),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_440),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_460),
.B(n_192),
.Y(n_491)
);

NOR3xp33_ASAP7_75t_L g492 ( 
.A(n_439),
.B(n_267),
.C(n_265),
.Y(n_492)
);

INVx8_ASAP7_75t_L g493 ( 
.A(n_456),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_415),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_450),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_397),
.B(n_270),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_404),
.B(n_272),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_351),
.B(n_220),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_441),
.B(n_229),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_370),
.B(n_274),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_411),
.B(n_383),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_388),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_386),
.B(n_235),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_403),
.B(n_237),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_370),
.B(n_164),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_456),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_385),
.A2(n_225),
.B1(n_204),
.B2(n_219),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_374),
.B(n_247),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_406),
.B(n_248),
.Y(n_509)
);

NAND3xp33_ASAP7_75t_L g510 ( 
.A(n_387),
.B(n_347),
.C(n_266),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_374),
.B(n_249),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_423),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_420),
.B(n_27),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_353),
.B(n_257),
.Y(n_514)
);

NOR3xp33_ASAP7_75t_L g515 ( 
.A(n_439),
.B(n_336),
.C(n_317),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_426),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_L g517 ( 
.A(n_376),
.B(n_260),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_355),
.B(n_262),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_357),
.B(n_263),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_364),
.B(n_264),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_429),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_364),
.B(n_269),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_380),
.B(n_377),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_388),
.B(n_219),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_444),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_445),
.Y(n_526)
);

OAI221xp5_ASAP7_75t_L g527 ( 
.A1(n_388),
.A2(n_187),
.B1(n_335),
.B2(n_307),
.C(n_321),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_448),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_401),
.B(n_336),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_363),
.B(n_165),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_449),
.Y(n_531)
);

AND3x1_ASAP7_75t_L g532 ( 
.A(n_356),
.B(n_225),
.C(n_242),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_401),
.B(n_307),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_453),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_419),
.B(n_347),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_424),
.B(n_347),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_399),
.B(n_307),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_379),
.B(n_209),
.Y(n_538)
);

OR2x6_ASAP7_75t_SL g539 ( 
.A(n_432),
.B(n_28),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_416),
.B(n_319),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_459),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_427),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_379),
.B(n_282),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_421),
.B(n_382),
.Y(n_544)
);

BUFx12f_ASAP7_75t_L g545 ( 
.A(n_369),
.Y(n_545)
);

NOR2x1p5_ASAP7_75t_L g546 ( 
.A(n_432),
.B(n_319),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_417),
.B(n_321),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_455),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_390),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_390),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_393),
.B(n_335),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_393),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_489),
.A2(n_412),
.B(n_409),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_467),
.B(n_417),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_525),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_523),
.A2(n_438),
.B1(n_369),
.B2(n_400),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_493),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_525),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_489),
.A2(n_412),
.B(n_409),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_487),
.Y(n_560)
);

NAND3xp33_ASAP7_75t_L g561 ( 
.A(n_542),
.B(n_413),
.C(n_409),
.Y(n_561)
);

O2A1O1Ixp33_ASAP7_75t_L g562 ( 
.A1(n_480),
.A2(n_469),
.B(n_501),
.C(n_542),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_465),
.B(n_468),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_SL g564 ( 
.A(n_486),
.B(n_438),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_486),
.A2(n_438),
.B1(n_396),
.B2(n_455),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_493),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_487),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_485),
.A2(n_431),
.B1(n_335),
.B2(n_313),
.Y(n_568)
);

AOI21x1_ASAP7_75t_L g569 ( 
.A1(n_529),
.A2(n_458),
.B(n_457),
.Y(n_569)
);

BUFx4f_ASAP7_75t_L g570 ( 
.A(n_486),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_484),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_543),
.A2(n_458),
.B(n_454),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_494),
.Y(n_573)
);

AOI21x1_ASAP7_75t_L g574 ( 
.A1(n_510),
.A2(n_454),
.B(n_452),
.Y(n_574)
);

INVxp67_ASAP7_75t_SL g575 ( 
.A(n_487),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_474),
.B(n_447),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_470),
.Y(n_577)
);

NAND3xp33_ASAP7_75t_L g578 ( 
.A(n_505),
.B(n_330),
.C(n_442),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_465),
.B(n_442),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_485),
.A2(n_470),
.B1(n_462),
.B2(n_500),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_471),
.B(n_478),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_524),
.A2(n_306),
.B1(n_313),
.B2(n_422),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_543),
.A2(n_452),
.B(n_451),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_535),
.A2(n_451),
.B(n_443),
.Y(n_584)
);

A2O1A1Ixp33_ASAP7_75t_L g585 ( 
.A1(n_536),
.A2(n_462),
.B(n_500),
.C(n_483),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_536),
.A2(n_436),
.B(n_435),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_524),
.B(n_29),
.Y(n_587)
);

AO22x1_ASAP7_75t_L g588 ( 
.A1(n_506),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_537),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_490),
.B(n_422),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_470),
.A2(n_306),
.B1(n_313),
.B2(n_422),
.Y(n_591)
);

AO21x1_ASAP7_75t_L g592 ( 
.A1(n_515),
.A2(n_434),
.B(n_433),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_468),
.A2(n_502),
.B1(n_477),
.B2(n_552),
.Y(n_593)
);

AND2x6_ASAP7_75t_SL g594 ( 
.A(n_539),
.B(n_31),
.Y(n_594)
);

O2A1O1Ixp33_ASAP7_75t_L g595 ( 
.A1(n_492),
.A2(n_527),
.B(n_496),
.C(n_497),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_502),
.A2(n_306),
.B1(n_313),
.B2(n_422),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_540),
.Y(n_597)
);

O2A1O1Ixp33_ASAP7_75t_L g598 ( 
.A1(n_492),
.A2(n_418),
.B(n_414),
.C(n_407),
.Y(n_598)
);

BUFx12f_ASAP7_75t_L g599 ( 
.A(n_545),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_493),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_547),
.Y(n_601)
);

O2A1O1Ixp33_ASAP7_75t_L g602 ( 
.A1(n_488),
.A2(n_497),
.B(n_496),
.C(n_513),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_470),
.Y(n_603)
);

OAI21xp33_ASAP7_75t_L g604 ( 
.A1(n_481),
.A2(n_505),
.B(n_483),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_550),
.A2(n_402),
.B(n_352),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_463),
.B(n_35),
.Y(n_606)
);

NOR3xp33_ASAP7_75t_L g607 ( 
.A(n_544),
.B(n_373),
.C(n_359),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_507),
.B(n_35),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_512),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_506),
.B(n_36),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_516),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_517),
.A2(n_375),
.B(n_391),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g613 ( 
.A1(n_515),
.A2(n_375),
.B(n_391),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_491),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_546),
.B(n_42),
.Y(n_615)
);

A2O1A1Ixp33_ASAP7_75t_L g616 ( 
.A1(n_549),
.A2(n_372),
.B(n_389),
.C(n_384),
.Y(n_616)
);

BUFx8_ASAP7_75t_SL g617 ( 
.A(n_548),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_521),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_L g619 ( 
.A1(n_541),
.A2(n_381),
.B(n_365),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_532),
.B(n_43),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_499),
.A2(n_508),
.B(n_511),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_509),
.B(n_48),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_526),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_528),
.B(n_531),
.Y(n_624)
);

O2A1O1Ixp5_ASAP7_75t_L g625 ( 
.A1(n_530),
.A2(n_361),
.B(n_358),
.C(n_395),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_534),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_464),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_466),
.Y(n_628)
);

A2O1A1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_461),
.A2(n_395),
.B(n_58),
.C(n_60),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_518),
.B(n_57),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_495),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_519),
.B(n_476),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_472),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_503),
.B(n_504),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_581),
.B(n_473),
.Y(n_635)
);

OAI21x1_ASAP7_75t_L g636 ( 
.A1(n_613),
.A2(n_533),
.B(n_538),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_585),
.A2(n_551),
.B(n_522),
.Y(n_637)
);

AOI221x1_ASAP7_75t_L g638 ( 
.A1(n_604),
.A2(n_520),
.B1(n_514),
.B2(n_395),
.C(n_482),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_580),
.B(n_498),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_SL g640 ( 
.A(n_595),
.B(n_479),
.C(n_475),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_570),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_580),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_571),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_570),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_632),
.B(n_65),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_634),
.A2(n_621),
.B(n_583),
.Y(n_646)
);

NOR2x1_ASAP7_75t_R g647 ( 
.A(n_599),
.B(n_67),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_573),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_557),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_572),
.A2(n_586),
.B(n_584),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_579),
.A2(n_597),
.B(n_589),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_614),
.B(n_72),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_602),
.B(n_73),
.Y(n_653)
);

AOI211x1_ASAP7_75t_L g654 ( 
.A1(n_563),
.A2(n_76),
.B(n_77),
.C(n_78),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_566),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_624),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_611),
.Y(n_657)
);

A2O1A1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_562),
.A2(n_103),
.B(n_105),
.C(n_106),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_618),
.Y(n_659)
);

OAI21xp5_ASAP7_75t_L g660 ( 
.A1(n_598),
.A2(n_116),
.B(n_118),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_560),
.Y(n_661)
);

CKINVDCx11_ASAP7_75t_R g662 ( 
.A(n_594),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_601),
.B(n_126),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_556),
.B(n_132),
.Y(n_664)
);

BUFx10_ASAP7_75t_L g665 ( 
.A(n_615),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_626),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_609),
.Y(n_667)
);

AO31x2_ASAP7_75t_L g668 ( 
.A1(n_629),
.A2(n_142),
.A3(n_145),
.B(n_146),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_593),
.B(n_587),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_631),
.B(n_632),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_623),
.Y(n_671)
);

BUFx12f_ASAP7_75t_L g672 ( 
.A(n_600),
.Y(n_672)
);

AO22x2_ASAP7_75t_L g673 ( 
.A1(n_565),
.A2(n_615),
.B1(n_608),
.B2(n_622),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_576),
.B(n_606),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_607),
.B(n_633),
.Y(n_675)
);

NOR4xp25_ASAP7_75t_L g676 ( 
.A(n_620),
.B(n_582),
.C(n_610),
.D(n_561),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_622),
.B(n_564),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_605),
.A2(n_619),
.B(n_558),
.Y(n_678)
);

AOI221xp5_ASAP7_75t_L g679 ( 
.A1(n_588),
.A2(n_568),
.B1(n_630),
.B2(n_555),
.C(n_627),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_577),
.B(n_603),
.Y(n_680)
);

O2A1O1Ixp33_ASAP7_75t_SL g681 ( 
.A1(n_616),
.A2(n_578),
.B(n_590),
.C(n_591),
.Y(n_681)
);

NAND3xp33_ASAP7_75t_L g682 ( 
.A(n_625),
.B(n_596),
.C(n_612),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_567),
.B(n_575),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_628),
.Y(n_684)
);

OAI22x1_ASAP7_75t_L g685 ( 
.A1(n_617),
.A2(n_297),
.B1(n_382),
.B2(n_507),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_553),
.A2(n_559),
.B(n_634),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_554),
.B(n_524),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_585),
.A2(n_602),
.B(n_595),
.C(n_621),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_571),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_569),
.A2(n_613),
.B(n_559),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_632),
.B(n_557),
.Y(n_691)
);

AOI21x1_ASAP7_75t_L g692 ( 
.A1(n_574),
.A2(n_569),
.B(n_559),
.Y(n_692)
);

INVx5_ASAP7_75t_L g693 ( 
.A(n_560),
.Y(n_693)
);

BUFx4_ASAP7_75t_SL g694 ( 
.A(n_594),
.Y(n_694)
);

OAI21x1_ASAP7_75t_L g695 ( 
.A1(n_569),
.A2(n_613),
.B(n_559),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_SL g696 ( 
.A1(n_580),
.A2(n_507),
.B(n_524),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_580),
.A2(n_524),
.B1(n_297),
.B2(n_474),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_585),
.A2(n_510),
.B(n_535),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_560),
.Y(n_699)
);

AOI221xp5_ASAP7_75t_SL g700 ( 
.A1(n_595),
.A2(n_602),
.B1(n_585),
.B2(n_562),
.C(n_604),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_560),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_554),
.B(n_474),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_617),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_570),
.Y(n_704)
);

AOI21x1_ASAP7_75t_L g705 ( 
.A1(n_574),
.A2(n_569),
.B(n_559),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_580),
.A2(n_524),
.B1(n_297),
.B2(n_474),
.Y(n_706)
);

AOI21xp33_ASAP7_75t_L g707 ( 
.A1(n_562),
.A2(n_420),
.B(n_371),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_585),
.A2(n_510),
.B(n_535),
.Y(n_708)
);

OAI21x1_ASAP7_75t_L g709 ( 
.A1(n_569),
.A2(n_613),
.B(n_559),
.Y(n_709)
);

OR2x6_ASAP7_75t_L g710 ( 
.A(n_557),
.B(n_486),
.Y(n_710)
);

NAND2x1p5_ASAP7_75t_L g711 ( 
.A(n_570),
.B(n_557),
.Y(n_711)
);

AO21x2_ASAP7_75t_L g712 ( 
.A1(n_592),
.A2(n_515),
.B(n_553),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_673),
.A2(n_669),
.B1(n_688),
.B2(n_656),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_696),
.B(n_687),
.Y(n_714)
);

AND2x2_ASAP7_75t_SL g715 ( 
.A(n_645),
.B(n_676),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_704),
.B(n_656),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_703),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_693),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_704),
.B(n_641),
.Y(n_719)
);

OAI21xp5_ASAP7_75t_L g720 ( 
.A1(n_698),
.A2(n_708),
.B(n_686),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_646),
.A2(n_650),
.B(n_678),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_643),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_707),
.A2(n_639),
.B(n_651),
.C(n_637),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_673),
.A2(n_640),
.B1(n_674),
.B2(n_697),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_648),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_702),
.B(n_706),
.Y(n_726)
);

AO21x2_ASAP7_75t_L g727 ( 
.A1(n_690),
.A2(n_709),
.B(n_695),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_635),
.B(n_657),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_648),
.Y(n_729)
);

OR2x6_ASAP7_75t_L g730 ( 
.A(n_710),
.B(n_711),
.Y(n_730)
);

OR3x4_ASAP7_75t_SL g731 ( 
.A(n_694),
.B(n_662),
.C(n_647),
.Y(n_731)
);

NOR2x1_ASAP7_75t_SL g732 ( 
.A(n_710),
.B(n_693),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_693),
.Y(n_733)
);

AO21x2_ASAP7_75t_L g734 ( 
.A1(n_712),
.A2(n_660),
.B(n_682),
.Y(n_734)
);

OAI21xp5_ASAP7_75t_L g735 ( 
.A1(n_653),
.A2(n_636),
.B(n_658),
.Y(n_735)
);

NAND3xp33_ASAP7_75t_L g736 ( 
.A(n_654),
.B(n_679),
.C(n_642),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_712),
.A2(n_681),
.B(n_663),
.Y(n_737)
);

NAND2x1p5_ASAP7_75t_L g738 ( 
.A(n_644),
.B(n_661),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_645),
.B(n_657),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_685),
.A2(n_677),
.B1(n_675),
.B2(n_670),
.Y(n_740)
);

OAI21x1_ASAP7_75t_SL g741 ( 
.A1(n_661),
.A2(n_664),
.B(n_680),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_689),
.B(n_667),
.Y(n_742)
);

OA21x2_ASAP7_75t_L g743 ( 
.A1(n_683),
.A2(n_666),
.B(n_659),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_672),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_691),
.B(n_684),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_671),
.Y(n_746)
);

BUFx2_ASAP7_75t_R g747 ( 
.A(n_655),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_652),
.B(n_665),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_665),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_649),
.B(n_701),
.Y(n_750)
);

INVx5_ASAP7_75t_L g751 ( 
.A(n_699),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_L g752 ( 
.A(n_699),
.B(n_654),
.C(n_700),
.Y(n_752)
);

NAND2x1p5_ASAP7_75t_L g753 ( 
.A(n_668),
.B(n_570),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_668),
.B(n_704),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_704),
.B(n_656),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_696),
.B(n_687),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_693),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_656),
.Y(n_758)
);

AO21x2_ASAP7_75t_L g759 ( 
.A1(n_692),
.A2(n_705),
.B(n_676),
.Y(n_759)
);

NAND2x1p5_ASAP7_75t_L g760 ( 
.A(n_704),
.B(n_570),
.Y(n_760)
);

OAI21xp5_ASAP7_75t_L g761 ( 
.A1(n_688),
.A2(n_585),
.B(n_708),
.Y(n_761)
);

AO21x2_ASAP7_75t_L g762 ( 
.A1(n_692),
.A2(n_705),
.B(n_676),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_672),
.Y(n_763)
);

AO21x2_ASAP7_75t_L g764 ( 
.A1(n_692),
.A2(n_705),
.B(n_676),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_702),
.B(n_480),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_656),
.Y(n_766)
);

BUFx2_ASAP7_75t_SL g767 ( 
.A(n_644),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_688),
.A2(n_585),
.B(n_708),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_656),
.Y(n_769)
);

OAI21xp5_ASAP7_75t_L g770 ( 
.A1(n_688),
.A2(n_585),
.B(n_708),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_673),
.A2(n_669),
.B1(n_688),
.B2(n_580),
.Y(n_771)
);

AO31x2_ASAP7_75t_L g772 ( 
.A1(n_688),
.A2(n_592),
.A3(n_638),
.B(n_686),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_725),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_739),
.B(n_758),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_758),
.B(n_766),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_729),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_751),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_766),
.B(n_769),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_751),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_765),
.B(n_728),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_751),
.Y(n_781)
);

INVx4_ASAP7_75t_L g782 ( 
.A(n_751),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_726),
.B(n_714),
.Y(n_783)
);

AO21x2_ASAP7_75t_L g784 ( 
.A1(n_721),
.A2(n_737),
.B(n_720),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_714),
.B(n_756),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_771),
.B(n_742),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_743),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_718),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_746),
.Y(n_789)
);

AO21x2_ASAP7_75t_L g790 ( 
.A1(n_735),
.A2(n_768),
.B(n_761),
.Y(n_790)
);

AO21x2_ASAP7_75t_L g791 ( 
.A1(n_735),
.A2(n_768),
.B(n_761),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_731),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_713),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_713),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_754),
.B(n_718),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_750),
.Y(n_796)
);

INVx4_ASAP7_75t_L g797 ( 
.A(n_730),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_722),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_754),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_733),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_716),
.Y(n_801)
);

AO21x2_ASAP7_75t_L g802 ( 
.A1(n_770),
.A2(n_752),
.B(n_759),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_723),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_716),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_755),
.Y(n_805)
);

INVx11_ASAP7_75t_L g806 ( 
.A(n_731),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_723),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_770),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_733),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_771),
.B(n_756),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_740),
.B(n_724),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_715),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_783),
.B(n_724),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_775),
.B(n_764),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_787),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_798),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_775),
.B(n_764),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_808),
.B(n_762),
.Y(n_818)
);

INVxp67_ASAP7_75t_SL g819 ( 
.A(n_778),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_778),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_785),
.B(n_745),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_780),
.B(n_745),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_773),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_810),
.A2(n_811),
.B1(n_786),
.B2(n_808),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_776),
.Y(n_825)
);

OR2x2_ASAP7_75t_L g826 ( 
.A(n_786),
.B(n_762),
.Y(n_826)
);

NAND3xp33_ASAP7_75t_L g827 ( 
.A(n_803),
.B(n_736),
.C(n_749),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_793),
.B(n_759),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_793),
.B(n_772),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_810),
.B(n_772),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_794),
.B(n_772),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_790),
.B(n_791),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_790),
.B(n_734),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_SL g834 ( 
.A1(n_797),
.A2(n_732),
.B1(n_753),
.B2(n_757),
.Y(n_834)
);

INVx4_ASAP7_75t_L g835 ( 
.A(n_774),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_791),
.B(n_727),
.Y(n_836)
);

OR2x6_ASAP7_75t_L g837 ( 
.A(n_774),
.B(n_741),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_777),
.Y(n_838)
);

AND2x2_ASAP7_75t_SL g839 ( 
.A(n_835),
.B(n_795),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_832),
.B(n_802),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_819),
.B(n_812),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_823),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_816),
.Y(n_843)
);

BUFx12f_ASAP7_75t_L g844 ( 
.A(n_838),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_824),
.B(n_807),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_815),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_832),
.B(n_828),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_823),
.B(n_807),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_828),
.B(n_802),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_829),
.B(n_802),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_829),
.B(n_799),
.Y(n_851)
);

INVxp33_ASAP7_75t_SL g852 ( 
.A(n_822),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_837),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_831),
.B(n_784),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_838),
.Y(n_855)
);

NOR2x1p5_ASAP7_75t_L g856 ( 
.A(n_853),
.B(n_792),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_843),
.B(n_820),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_847),
.B(n_813),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_847),
.B(n_836),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_853),
.B(n_837),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_853),
.B(n_837),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_854),
.B(n_836),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_842),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_854),
.B(n_818),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_850),
.B(n_814),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_851),
.B(n_814),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_846),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_850),
.B(n_818),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_845),
.B(n_825),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_840),
.B(n_833),
.Y(n_870)
);

OR2x6_ASAP7_75t_L g871 ( 
.A(n_844),
.B(n_837),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_840),
.B(n_817),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_863),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_857),
.Y(n_874)
);

AND2x2_ASAP7_75t_SL g875 ( 
.A(n_860),
.B(n_839),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_867),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_858),
.B(n_852),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_866),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_859),
.B(n_849),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_859),
.B(n_849),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_869),
.Y(n_881)
);

OR2x2_ASAP7_75t_L g882 ( 
.A(n_872),
.B(n_817),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_862),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_881),
.B(n_870),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_SL g885 ( 
.A1(n_875),
.A2(n_792),
.B1(n_871),
.B2(n_839),
.Y(n_885)
);

OAI322xp33_ASAP7_75t_L g886 ( 
.A1(n_874),
.A2(n_865),
.A3(n_872),
.B1(n_841),
.B2(n_830),
.C1(n_848),
.C2(n_826),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_876),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_877),
.Y(n_888)
);

AOI21xp33_ASAP7_75t_L g889 ( 
.A1(n_877),
.A2(n_827),
.B(n_848),
.Y(n_889)
);

O2A1O1Ixp33_ASAP7_75t_SL g890 ( 
.A1(n_875),
.A2(n_806),
.B(n_855),
.C(n_856),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_878),
.A2(n_883),
.B1(n_861),
.B2(n_860),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_873),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_879),
.B(n_864),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_890),
.A2(n_871),
.B(n_839),
.Y(n_894)
);

OR2x2_ASAP7_75t_L g895 ( 
.A(n_884),
.B(n_882),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_885),
.A2(n_860),
.B1(n_861),
.B2(n_882),
.Y(n_896)
);

AOI221xp5_ASAP7_75t_L g897 ( 
.A1(n_886),
.A2(n_880),
.B1(n_879),
.B2(n_864),
.C(n_868),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_896),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_897),
.B(n_887),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_895),
.B(n_888),
.Y(n_900)
);

OAI21xp33_ASAP7_75t_SL g901 ( 
.A1(n_899),
.A2(n_894),
.B(n_893),
.Y(n_901)
);

OAI211xp5_ASAP7_75t_L g902 ( 
.A1(n_898),
.A2(n_890),
.B(n_889),
.C(n_763),
.Y(n_902)
);

NOR2x1_ASAP7_75t_L g903 ( 
.A(n_902),
.B(n_763),
.Y(n_903)
);

NOR2x1_ASAP7_75t_L g904 ( 
.A(n_901),
.B(n_730),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_903),
.Y(n_905)
);

AO22x1_ASAP7_75t_SL g906 ( 
.A1(n_904),
.A2(n_806),
.B1(n_744),
.B2(n_717),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_905),
.A2(n_900),
.B1(n_891),
.B2(n_717),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_906),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_908),
.Y(n_909)
);

OAI211xp5_ASAP7_75t_L g910 ( 
.A1(n_907),
.A2(n_905),
.B(n_797),
.C(n_747),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_908),
.A2(n_827),
.B(n_760),
.Y(n_911)
);

OAI21x1_ASAP7_75t_L g912 ( 
.A1(n_909),
.A2(n_760),
.B(n_747),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_910),
.A2(n_911),
.B(n_797),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_909),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_909),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_909),
.A2(n_871),
.B1(n_861),
.B2(n_767),
.Y(n_916)
);

XOR2x2_ASAP7_75t_L g917 ( 
.A(n_913),
.B(n_719),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_915),
.B(n_892),
.Y(n_918)
);

NOR3xp33_ASAP7_75t_L g919 ( 
.A(n_912),
.B(n_782),
.C(n_748),
.Y(n_919)
);

OAI331xp33_ASAP7_75t_L g920 ( 
.A1(n_916),
.A2(n_789),
.A3(n_796),
.B1(n_821),
.B2(n_801),
.B3(n_804),
.C1(n_805),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_914),
.Y(n_921)
);

XNOR2x1_ASAP7_75t_L g922 ( 
.A(n_912),
.B(n_738),
.Y(n_922)
);

AO221x1_ASAP7_75t_L g923 ( 
.A1(n_921),
.A2(n_788),
.B1(n_800),
.B2(n_809),
.C(n_781),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_922),
.A2(n_738),
.B(n_834),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_918),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_923),
.A2(n_919),
.B1(n_917),
.B2(n_920),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_925),
.A2(n_871),
.B1(n_782),
.B2(n_781),
.Y(n_927)
);

XOR2xp5_ASAP7_75t_L g928 ( 
.A(n_926),
.B(n_924),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_928),
.A2(n_927),
.B1(n_781),
.B2(n_779),
.Y(n_929)
);


endmodule