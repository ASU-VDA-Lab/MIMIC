module fake_netlist_6_4788_n_1275 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_341, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_338, n_56, n_119, n_235, n_147, n_191, n_340, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_334, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1275);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_341;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_338;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1275;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_694;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_615;
wire n_1249;
wire n_1127;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_526;
wire n_1183;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_537;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_548;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_670;
wire n_1089;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_965;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_102),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_92),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_178),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_40),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_170),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_89),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_131),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_28),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_221),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_95),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_294),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_72),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_158),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_3),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_199),
.Y(n_356)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_164),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_166),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_143),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_332),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_160),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_140),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_248),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_93),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_20),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_308),
.Y(n_366)
);

BUFx5_ASAP7_75t_L g367 ( 
.A(n_338),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_2),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_47),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_159),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_161),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_58),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_289),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_202),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_188),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_245),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_325),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_11),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_210),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_147),
.Y(n_380)
);

INVxp67_ASAP7_75t_R g381 ( 
.A(n_184),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_284),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_241),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_25),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_57),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_209),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_112),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_273),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_78),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_187),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_100),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_230),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_192),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_341),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_198),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_287),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_326),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_141),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_201),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_286),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_204),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_105),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_86),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_181),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_265),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_171),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_116),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_68),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_3),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_253),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_73),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_274),
.Y(n_412)
);

BUFx5_ASAP7_75t_L g413 ( 
.A(n_271),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_63),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_45),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_31),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_148),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_125),
.Y(n_418)
);

BUFx10_ASAP7_75t_L g419 ( 
.A(n_303),
.Y(n_419)
);

BUFx10_ASAP7_75t_L g420 ( 
.A(n_121),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_239),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_9),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_312),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_152),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_214),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_279),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_35),
.Y(n_427)
);

BUFx10_ASAP7_75t_L g428 ( 
.A(n_57),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_114),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_89),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_224),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_306),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_200),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_216),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_231),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_156),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_222),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_28),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_219),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_247),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_68),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_56),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_142),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_269),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_328),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_75),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_0),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_R g448 ( 
.A(n_218),
.B(n_275),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_165),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_10),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_136),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_217),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_297),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_120),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_8),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_53),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_144),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_77),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_242),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_240),
.Y(n_460)
);

NOR2xp67_ASAP7_75t_L g461 ( 
.A(n_205),
.B(n_49),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_285),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_79),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_91),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_262),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_62),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_167),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_268),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_122),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_227),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_76),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_314),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_203),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_29),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_208),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_72),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_330),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_150),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_256),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_195),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_83),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_290),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_182),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_194),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_151),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_97),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_101),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_73),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_119),
.Y(n_489)
);

CKINVDCx14_ASAP7_75t_R g490 ( 
.A(n_329),
.Y(n_490)
);

BUFx5_ASAP7_75t_L g491 ( 
.A(n_139),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_229),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_197),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_322),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_137),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_7),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_135),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_333),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_115),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_132),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_189),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_104),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_98),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_26),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_145),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_276),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_146),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_311),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_153),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_254),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_433),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_433),
.Y(n_512)
);

BUFx8_ASAP7_75t_SL g513 ( 
.A(n_385),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_368),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_419),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_0),
.Y(n_516)
);

OAI22x1_ASAP7_75t_SL g517 ( 
.A1(n_456),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_368),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_442),
.Y(n_519)
);

BUFx12f_ASAP7_75t_L g520 ( 
.A(n_428),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_384),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_471),
.A2(n_5),
.B1(n_1),
.B2(n_4),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_384),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_384),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_463),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_463),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_345),
.Y(n_527)
);

OAI22x1_ASAP7_75t_SL g528 ( 
.A1(n_481),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_528)
);

AOI22x1_ASAP7_75t_SL g529 ( 
.A1(n_349),
.A2(n_9),
.B1(n_6),
.B2(n_8),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_357),
.B(n_10),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_343),
.B(n_11),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_463),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_448),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_433),
.Y(n_535)
);

BUFx12f_ASAP7_75t_L g536 ( 
.A(n_476),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_409),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_453),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_363),
.B(n_12),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_453),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_374),
.B(n_12),
.Y(n_541)
);

OAI22x1_ASAP7_75t_R g542 ( 
.A1(n_353),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_367),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_460),
.B(n_13),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_496),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_453),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_446),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_367),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_367),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_415),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_380),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_365),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_387),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_490),
.B(n_17),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_436),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_367),
.Y(n_556)
);

INVx5_ASAP7_75t_L g557 ( 
.A(n_420),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_367),
.Y(n_558)
);

BUFx8_ASAP7_75t_L g559 ( 
.A(n_347),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_500),
.B(n_19),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_355),
.Y(n_561)
);

BUFx8_ASAP7_75t_SL g562 ( 
.A(n_342),
.Y(n_562)
);

BUFx8_ASAP7_75t_L g563 ( 
.A(n_369),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_506),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_420),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_376),
.B(n_19),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_414),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_477),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_359),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_509),
.B(n_20),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_344),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_372),
.Y(n_572)
);

INVx5_ASAP7_75t_L g573 ( 
.A(n_362),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_378),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_370),
.Y(n_575)
);

CKINVDCx16_ASAP7_75t_R g576 ( 
.A(n_364),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_416),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_479),
.B(n_21),
.Y(n_578)
);

OAI22x1_ASAP7_75t_R g579 ( 
.A1(n_389),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_579)
);

BUFx12f_ASAP7_75t_L g580 ( 
.A(n_403),
.Y(n_580)
);

BUFx12f_ASAP7_75t_L g581 ( 
.A(n_408),
.Y(n_581)
);

INVx6_ASAP7_75t_L g582 ( 
.A(n_413),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_422),
.A2(n_450),
.B1(n_455),
.B2(n_438),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_458),
.Y(n_584)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_413),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_346),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_348),
.Y(n_587)
);

BUFx12f_ASAP7_75t_L g588 ( 
.A(n_411),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_354),
.Y(n_589)
);

AOI21x1_ASAP7_75t_L g590 ( 
.A1(n_543),
.A2(n_549),
.B(n_548),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_562),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_513),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_576),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_511),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_571),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_576),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_R g597 ( 
.A(n_572),
.B(n_427),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_R g598 ( 
.A(n_534),
.B(n_383),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_586),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_568),
.B(n_589),
.Y(n_600)
);

BUFx10_ASAP7_75t_L g601 ( 
.A(n_530),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_515),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_580),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_511),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_581),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_588),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_531),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_589),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_520),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_582),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_568),
.B(n_350),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_R g612 ( 
.A(n_527),
.B(n_430),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_574),
.B(n_454),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_R g614 ( 
.A(n_565),
.B(n_386),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_518),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_523),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_537),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_536),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_524),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_525),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_557),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_559),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_557),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_557),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_R g625 ( 
.A(n_565),
.B(n_390),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_559),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_519),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_533),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_568),
.B(n_351),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_551),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_512),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_512),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_512),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_R g634 ( 
.A(n_532),
.B(n_441),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_564),
.B(n_470),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_R g636 ( 
.A(n_541),
.B(n_435),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_551),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_564),
.B(n_352),
.Y(n_638)
);

NOR2xp67_ASAP7_75t_L g639 ( 
.A(n_585),
.B(n_371),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_590),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_613),
.B(n_556),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_594),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_627),
.Y(n_643)
);

NAND2xp33_ASAP7_75t_L g644 ( 
.A(n_636),
.B(n_554),
.Y(n_644)
);

BUFx5_ASAP7_75t_L g645 ( 
.A(n_632),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_635),
.B(n_558),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_610),
.B(n_573),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_610),
.B(n_573),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_610),
.B(n_573),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_610),
.B(n_566),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_594),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_608),
.B(n_544),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_595),
.B(n_553),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_604),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_633),
.B(n_566),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_602),
.B(n_553),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_615),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_620),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_599),
.B(n_555),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_628),
.B(n_569),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_616),
.Y(n_661)
);

INVxp67_ASAP7_75t_SL g662 ( 
.A(n_639),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_619),
.B(n_569),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_614),
.B(n_555),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_638),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_601),
.B(n_570),
.Y(n_666)
);

NOR3xp33_ASAP7_75t_L g667 ( 
.A(n_617),
.B(n_552),
.C(n_570),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_630),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_637),
.B(n_516),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_600),
.B(n_569),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_611),
.B(n_575),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_612),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_629),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_621),
.B(n_575),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_623),
.B(n_575),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_607),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_624),
.B(n_560),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_625),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_617),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_626),
.B(n_539),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_603),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_605),
.B(n_535),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_606),
.B(n_535),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_618),
.B(n_521),
.Y(n_684)
);

NOR3xp33_ASAP7_75t_L g685 ( 
.A(n_592),
.B(n_552),
.C(n_522),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_L g686 ( 
.A(n_634),
.B(n_578),
.C(n_545),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_598),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_609),
.Y(n_688)
);

BUFx5_ASAP7_75t_L g689 ( 
.A(n_634),
.Y(n_689)
);

OAI21xp33_ASAP7_75t_L g690 ( 
.A1(n_597),
.A2(n_578),
.B(n_545),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_622),
.B(n_457),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_597),
.B(n_538),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_593),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_596),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_591),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_612),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_613),
.B(n_538),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_631),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_613),
.B(n_521),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_627),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_613),
.B(n_538),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_590),
.Y(n_702)
);

AO221x1_ASAP7_75t_L g703 ( 
.A1(n_607),
.A2(n_583),
.B1(n_522),
.B2(n_379),
.C(n_366),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_613),
.B(n_526),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_676),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_676),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_676),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_689),
.B(n_445),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_687),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_666),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_657),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_656),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_698),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_652),
.B(n_462),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_658),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_679),
.B(n_561),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_699),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_661),
.Y(n_718)
);

NOR2x2_ASAP7_75t_L g719 ( 
.A(n_703),
.B(n_542),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_642),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_689),
.B(n_468),
.Y(n_721)
);

BUFx6f_ASAP7_75t_SL g722 ( 
.A(n_693),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_665),
.B(n_443),
.Y(n_723)
);

AND3x1_ASAP7_75t_L g724 ( 
.A(n_685),
.B(n_579),
.C(n_542),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_660),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_689),
.A2(n_449),
.B1(n_485),
.B2(n_461),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_640),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_654),
.Y(n_728)
);

OAI22xp33_ASAP7_75t_L g729 ( 
.A1(n_686),
.A2(n_381),
.B1(n_377),
.B2(n_360),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_669),
.B(n_391),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_663),
.Y(n_731)
);

CKINVDCx6p67_ASAP7_75t_R g732 ( 
.A(n_691),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_704),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_689),
.A2(n_358),
.B1(n_361),
.B2(n_356),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_SL g735 ( 
.A1(n_672),
.A2(n_694),
.B1(n_583),
.B2(n_643),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_646),
.B(n_394),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_668),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_702),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_663),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_692),
.B(n_447),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_SL g741 ( 
.A1(n_700),
.A2(n_579),
.B1(n_528),
.B2(n_517),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_651),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_686),
.A2(n_401),
.B1(n_405),
.B2(n_396),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_690),
.A2(n_375),
.B1(n_382),
.B2(n_373),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_667),
.A2(n_417),
.B1(n_421),
.B2(n_412),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_655),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_646),
.B(n_424),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_641),
.A2(n_429),
.B1(n_440),
.B2(n_432),
.Y(n_748)
);

AND3x1_ASAP7_75t_SL g749 ( 
.A(n_681),
.B(n_488),
.C(n_474),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_697),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_671),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_673),
.A2(n_469),
.B1(n_478),
.B2(n_472),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_644),
.A2(n_480),
.B1(n_483),
.B2(n_482),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_L g754 ( 
.A1(n_701),
.A2(n_484),
.B1(n_487),
.B2(n_486),
.Y(n_754)
);

BUFx2_ASAP7_75t_L g755 ( 
.A(n_684),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_674),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_670),
.B(n_492),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_645),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_653),
.B(n_659),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_664),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_645),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_R g762 ( 
.A(n_695),
.B(n_388),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_678),
.B(n_466),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_662),
.B(n_493),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_671),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_645),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_688),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_650),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_677),
.B(n_494),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_R g770 ( 
.A(n_682),
.B(n_392),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_675),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_680),
.A2(n_499),
.B1(n_502),
.B2(n_495),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_647),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_683),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_648),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_649),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_689),
.B(n_393),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_689),
.B(n_395),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_692),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_676),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_699),
.B(n_567),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_660),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_643),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_676),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_696),
.A2(n_398),
.B1(n_399),
.B2(n_397),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_676),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_667),
.A2(n_491),
.B1(n_413),
.B2(n_587),
.Y(n_787)
);

NOR2x2_ASAP7_75t_L g788 ( 
.A(n_679),
.B(n_517),
.Y(n_788)
);

OR2x2_ASAP7_75t_SL g789 ( 
.A(n_696),
.B(n_528),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_656),
.B(n_584),
.Y(n_790)
);

AOI22x1_ASAP7_75t_L g791 ( 
.A1(n_640),
.A2(n_547),
.B1(n_402),
.B2(n_404),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_699),
.B(n_567),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_667),
.A2(n_491),
.B1(n_413),
.B2(n_504),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_SL g794 ( 
.A1(n_652),
.A2(n_529),
.B1(n_547),
.B2(n_563),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_707),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_746),
.B(n_400),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_710),
.B(n_577),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_751),
.B(n_406),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_714),
.B(n_563),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_705),
.B(n_577),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_779),
.B(n_407),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_756),
.B(n_410),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_765),
.B(n_418),
.Y(n_803)
);

NOR2xp67_ASAP7_75t_L g804 ( 
.A(n_767),
.B(n_709),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_759),
.B(n_423),
.Y(n_805)
);

NOR3xp33_ASAP7_75t_L g806 ( 
.A(n_735),
.B(n_426),
.C(n_425),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_731),
.B(n_431),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_739),
.B(n_434),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_707),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_753),
.A2(n_437),
.B1(n_444),
.B2(n_439),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_715),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_727),
.A2(n_738),
.B1(n_730),
.B2(n_708),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_780),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_740),
.A2(n_451),
.B(n_459),
.C(n_452),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_766),
.A2(n_546),
.B(n_540),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_727),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_R g817 ( 
.A(n_783),
.B(n_464),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_738),
.A2(n_465),
.B1(n_473),
.B2(n_467),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_780),
.B(n_550),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_755),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_725),
.B(n_475),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_780),
.Y(n_822)
);

AO32x2_ASAP7_75t_L g823 ( 
.A1(n_743),
.A2(n_491),
.A3(n_413),
.B1(n_25),
.B2(n_23),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_767),
.B(n_489),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_784),
.Y(n_825)
);

HAxp5_ASAP7_75t_L g826 ( 
.A(n_724),
.B(n_24),
.CON(n_826),
.SN(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_722),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_777),
.A2(n_498),
.B(n_497),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_784),
.B(n_501),
.Y(n_829)
);

NAND3xp33_ASAP7_75t_SL g830 ( 
.A(n_794),
.B(n_505),
.C(n_503),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_782),
.B(n_507),
.Y(n_831)
);

XOR2x2_ASAP7_75t_L g832 ( 
.A(n_741),
.B(n_24),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_778),
.A2(n_510),
.B(n_508),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_763),
.B(n_26),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_723),
.A2(n_582),
.B1(n_514),
.B2(n_585),
.Y(n_835)
);

INVx4_ASAP7_75t_L g836 ( 
.A(n_786),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_706),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_712),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_750),
.B(n_27),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_726),
.A2(n_585),
.B1(n_94),
.B2(n_96),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_717),
.B(n_27),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_737),
.Y(n_842)
);

BUFx4f_ASAP7_75t_SL g843 ( 
.A(n_732),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_733),
.B(n_99),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_718),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_716),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_790),
.B(n_103),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_760),
.B(n_30),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_768),
.A2(n_771),
.B1(n_769),
.B2(n_773),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_774),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_781),
.B(n_792),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_729),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_758),
.A2(n_761),
.B(n_771),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_790),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_742),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_722),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_742),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_793),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_773),
.A2(n_107),
.B1(n_108),
.B2(n_106),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_736),
.A2(n_110),
.B(n_109),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_747),
.A2(n_113),
.B(n_111),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_776),
.A2(n_118),
.B(n_117),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_785),
.B(n_764),
.Y(n_863)
);

INVx5_ASAP7_75t_L g864 ( 
.A(n_775),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_757),
.A2(n_124),
.B(n_123),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_748),
.B(n_36),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_720),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_745),
.B(n_37),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_734),
.B(n_126),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_713),
.B(n_38),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_789),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_728),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_744),
.A2(n_128),
.B1(n_129),
.B2(n_127),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_754),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_762),
.B(n_41),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_770),
.B(n_42),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_787),
.B(n_43),
.Y(n_877)
);

OAI21x1_ASAP7_75t_L g878 ( 
.A1(n_752),
.A2(n_772),
.B(n_791),
.Y(n_878)
);

BUFx4f_ASAP7_75t_L g879 ( 
.A(n_749),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_719),
.A2(n_133),
.B(n_130),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_788),
.B(n_43),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_711),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_746),
.B(n_44),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_SL g884 ( 
.A(n_714),
.B(n_134),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_727),
.Y(n_885)
);

NOR3xp33_ASAP7_75t_SL g886 ( 
.A(n_741),
.B(n_46),
.C(n_47),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_721),
.A2(n_50),
.B(n_46),
.C(n_48),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_746),
.B(n_51),
.Y(n_888)
);

CKINVDCx6p67_ASAP7_75t_R g889 ( 
.A(n_722),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_707),
.B(n_138),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_746),
.B(n_51),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_707),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_710),
.B(n_52),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_746),
.B(n_54),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_707),
.Y(n_895)
);

OA22x2_ASAP7_75t_L g896 ( 
.A1(n_741),
.A2(n_58),
.B1(n_55),
.B2(n_56),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_710),
.B(n_55),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_746),
.B(n_59),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_710),
.B(n_59),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_711),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_R g901 ( 
.A(n_709),
.B(n_149),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_711),
.Y(n_902)
);

O2A1O1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_721),
.A2(n_63),
.B(n_60),
.C(n_61),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_707),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_707),
.B(n_154),
.Y(n_905)
);

NAND2x1p5_ASAP7_75t_L g906 ( 
.A(n_707),
.B(n_155),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_710),
.B(n_60),
.Y(n_907)
);

BUFx12f_ASAP7_75t_L g908 ( 
.A(n_707),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_714),
.A2(n_65),
.B(n_61),
.C(n_64),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_710),
.B(n_64),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_711),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_851),
.B(n_157),
.Y(n_912)
);

AOI22x1_ASAP7_75t_L g913 ( 
.A1(n_853),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_913)
);

BUFx12f_ASAP7_75t_L g914 ( 
.A(n_837),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_816),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_908),
.Y(n_916)
);

INVxp67_ASAP7_75t_SL g917 ( 
.A(n_855),
.Y(n_917)
);

INVxp67_ASAP7_75t_SL g918 ( 
.A(n_855),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_885),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_812),
.A2(n_163),
.B(n_162),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_820),
.Y(n_921)
);

BUFx12f_ASAP7_75t_L g922 ( 
.A(n_837),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_843),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_842),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_836),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_813),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_813),
.Y(n_927)
);

BUFx12f_ASAP7_75t_L g928 ( 
.A(n_827),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_850),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_838),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_863),
.A2(n_169),
.B(n_168),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_904),
.Y(n_932)
);

INVx6_ASAP7_75t_SL g933 ( 
.A(n_890),
.Y(n_933)
);

OA21x2_ASAP7_75t_L g934 ( 
.A1(n_878),
.A2(n_173),
.B(n_172),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_819),
.Y(n_935)
);

NAND2x1p5_ASAP7_75t_L g936 ( 
.A(n_857),
.B(n_174),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_846),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_817),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_889),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_795),
.B(n_175),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_797),
.B(n_800),
.Y(n_941)
);

OR2x6_ASAP7_75t_L g942 ( 
.A(n_804),
.B(n_66),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_856),
.Y(n_943)
);

INVx6_ASAP7_75t_L g944 ( 
.A(n_904),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_854),
.B(n_176),
.Y(n_945)
);

OAI21x1_ASAP7_75t_SL g946 ( 
.A1(n_887),
.A2(n_179),
.B(n_177),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_844),
.B(n_180),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_799),
.B(n_67),
.Y(n_948)
);

BUFx2_ASAP7_75t_R g949 ( 
.A(n_822),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_844),
.B(n_183),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_811),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_805),
.B(n_69),
.Y(n_952)
);

NAND3xp33_ASAP7_75t_L g953 ( 
.A(n_834),
.B(n_806),
.C(n_801),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_882),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_825),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_796),
.B(n_70),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_849),
.A2(n_186),
.B(n_185),
.Y(n_957)
);

AO21x2_ASAP7_75t_L g958 ( 
.A1(n_869),
.A2(n_191),
.B(n_190),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_825),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_841),
.B(n_70),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_883),
.B(n_71),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_895),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_884),
.A2(n_264),
.B1(n_340),
.B2(n_339),
.Y(n_963)
);

BUFx3_ASAP7_75t_L g964 ( 
.A(n_825),
.Y(n_964)
);

NAND2x1p5_ASAP7_75t_L g965 ( 
.A(n_892),
.B(n_193),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_L g966 ( 
.A1(n_868),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_892),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_900),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_892),
.Y(n_969)
);

INVx8_ASAP7_75t_L g970 ( 
.A(n_905),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_902),
.Y(n_971)
);

AND2x6_ASAP7_75t_L g972 ( 
.A(n_905),
.B(n_196),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_888),
.B(n_74),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_911),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_802),
.A2(n_267),
.B1(n_337),
.B2(n_336),
.Y(n_975)
);

CKINVDCx6p67_ASAP7_75t_R g976 ( 
.A(n_871),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_893),
.B(n_77),
.Y(n_977)
);

OR3x4_ASAP7_75t_SL g978 ( 
.A(n_826),
.B(n_78),
.C(n_79),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_845),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_891),
.B(n_80),
.Y(n_980)
);

INVx3_ASAP7_75t_SL g981 ( 
.A(n_847),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_894),
.B(n_80),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_867),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_870),
.Y(n_984)
);

INVx6_ASAP7_75t_SL g985 ( 
.A(n_879),
.Y(n_985)
);

NAND3xp33_ASAP7_75t_L g986 ( 
.A(n_858),
.B(n_81),
.C(n_82),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_898),
.B(n_81),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_798),
.B(n_82),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_872),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_897),
.B(n_83),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_899),
.B(n_84),
.Y(n_991)
);

OR2x6_ASAP7_75t_L g992 ( 
.A(n_880),
.B(n_84),
.Y(n_992)
);

OAI21x1_ASAP7_75t_SL g993 ( 
.A1(n_903),
.A2(n_277),
.B(n_335),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_907),
.B(n_85),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_809),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_876),
.Y(n_996)
);

BUFx2_ASAP7_75t_R g997 ( 
.A(n_877),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_803),
.A2(n_272),
.B(n_334),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_875),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_829),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_906),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_910),
.Y(n_1002)
);

BUFx4f_ASAP7_75t_L g1003 ( 
.A(n_901),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_864),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_848),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_821),
.Y(n_1006)
);

BUFx4_ASAP7_75t_SL g1007 ( 
.A(n_896),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_SL g1008 ( 
.A1(n_862),
.A2(n_270),
.B(n_331),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_866),
.Y(n_1009)
);

INVxp33_ASAP7_75t_L g1010 ( 
.A(n_839),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_807),
.B(n_85),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_808),
.B(n_86),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_831),
.Y(n_1013)
);

BUFx12f_ASAP7_75t_L g1014 ( 
.A(n_886),
.Y(n_1014)
);

OA21x2_ASAP7_75t_L g1015 ( 
.A1(n_815),
.A2(n_266),
.B(n_327),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_832),
.Y(n_1016)
);

AOI22x1_ASAP7_75t_L g1017 ( 
.A1(n_860),
.A2(n_87),
.B1(n_88),
.B2(n_90),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_823),
.Y(n_1018)
);

AO21x2_ASAP7_75t_L g1019 ( 
.A1(n_814),
.A2(n_278),
.B(n_324),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_824),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_823),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_823),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_830),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_881),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_818),
.B(n_87),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_859),
.Y(n_1026)
);

INVxp33_ASAP7_75t_L g1027 ( 
.A(n_921),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_914),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_919),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_915),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_R g1031 ( 
.A(n_943),
.B(n_206),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_1004),
.Y(n_1032)
);

INVx4_ASAP7_75t_L g1033 ( 
.A(n_922),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_926),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_929),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_941),
.B(n_909),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_953),
.A2(n_810),
.B1(n_840),
.B2(n_873),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_1013),
.A2(n_828),
.B(n_833),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_983),
.Y(n_1039)
);

OAI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_1010),
.A2(n_835),
.B1(n_861),
.B2(n_865),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_SL g1041 ( 
.A1(n_948),
.A2(n_852),
.B1(n_874),
.B2(n_90),
.Y(n_1041)
);

CKINVDCx6p67_ASAP7_75t_R g1042 ( 
.A(n_928),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_952),
.A2(n_207),
.B1(n_211),
.B2(n_212),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1006),
.B(n_213),
.Y(n_1044)
);

BUFx8_ASAP7_75t_L g1045 ( 
.A(n_996),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_1025),
.A2(n_215),
.B1(n_220),
.B2(n_223),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_990),
.A2(n_225),
.B1(n_226),
.B2(n_228),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_930),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1009),
.B(n_935),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_924),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_956),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_1051)
);

OAI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_1023),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_SL g1053 ( 
.A1(n_1016),
.A2(n_238),
.B1(n_243),
.B2(n_244),
.Y(n_1053)
);

INVx5_ASAP7_75t_L g1054 ( 
.A(n_959),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_971),
.Y(n_1055)
);

OA21x2_ASAP7_75t_L g1056 ( 
.A1(n_957),
.A2(n_246),
.B(n_249),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_923),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_971),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_927),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_SL g1060 ( 
.A1(n_1002),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_1060)
);

INVx8_ASAP7_75t_L g1061 ( 
.A(n_970),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_979),
.Y(n_1062)
);

OAI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_1005),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_1063)
);

NAND2xp33_ASAP7_75t_SL g1064 ( 
.A(n_981),
.B(n_259),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_970),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_986),
.A2(n_260),
.B1(n_261),
.B2(n_263),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_962),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_951),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_960),
.B(n_937),
.Y(n_1069)
);

BUFx4f_ASAP7_75t_SL g1070 ( 
.A(n_985),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_954),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_977),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_968),
.Y(n_1073)
);

OAI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_938),
.A2(n_283),
.B1(n_288),
.B2(n_291),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_974),
.Y(n_1075)
);

BUFx4f_ASAP7_75t_SL g1076 ( 
.A(n_985),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_984),
.B(n_292),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_991),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.Y(n_1078)
);

BUFx4f_ASAP7_75t_SL g1079 ( 
.A(n_933),
.Y(n_1079)
);

AO21x2_ASAP7_75t_L g1080 ( 
.A1(n_920),
.A2(n_298),
.B(n_299),
.Y(n_1080)
);

AOI21x1_ASAP7_75t_L g1081 ( 
.A1(n_984),
.A2(n_323),
.B(n_300),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_916),
.Y(n_1082)
);

AOI222xp33_ASAP7_75t_L g1083 ( 
.A1(n_966),
.A2(n_301),
.B1(n_302),
.B2(n_304),
.C1(n_305),
.C2(n_307),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_933),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_912),
.A2(n_309),
.B1(n_310),
.B2(n_313),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_944),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_SL g1087 ( 
.A(n_949),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1026),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_995),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_994),
.B(n_999),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_947),
.B(n_318),
.Y(n_1091)
);

BUFx2_ASAP7_75t_R g1092 ( 
.A(n_1024),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_912),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_932),
.Y(n_1094)
);

OAI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_999),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_989),
.Y(n_1096)
);

CKINVDCx11_ASAP7_75t_R g1097 ( 
.A(n_939),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_976),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_967),
.Y(n_1099)
);

OAI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_992),
.A2(n_942),
.B1(n_1003),
.B2(n_1011),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_1007),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_950),
.A2(n_1012),
.B1(n_988),
.B2(n_945),
.Y(n_1102)
);

OR2x2_ASAP7_75t_L g1103 ( 
.A(n_961),
.B(n_982),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_969),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_997),
.B(n_992),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_913),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_SL g1107 ( 
.A1(n_972),
.A2(n_1020),
.B1(n_1000),
.B2(n_1014),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_964),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_955),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_944),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_913),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1029),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_SL g1113 ( 
.A1(n_1083),
.A2(n_1041),
.B(n_1100),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1038),
.A2(n_998),
.B(n_931),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_1097),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_1035),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_1049),
.B(n_973),
.Y(n_1117)
);

NAND2xp33_ASAP7_75t_R g1118 ( 
.A(n_1057),
.B(n_1031),
.Y(n_1118)
);

NAND2xp33_ASAP7_75t_R g1119 ( 
.A(n_1084),
.B(n_925),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1102),
.A2(n_1036),
.B1(n_1090),
.B2(n_1037),
.Y(n_1120)
);

CKINVDCx16_ASAP7_75t_R g1121 ( 
.A(n_1087),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1030),
.Y(n_1122)
);

AO31x2_ASAP7_75t_L g1123 ( 
.A1(n_1106),
.A2(n_1022),
.A3(n_1018),
.B(n_980),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1069),
.B(n_987),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_1108),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_R g1126 ( 
.A(n_1070),
.B(n_1076),
.Y(n_1126)
);

OR2x6_ASAP7_75t_L g1127 ( 
.A(n_1061),
.B(n_942),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1103),
.B(n_1020),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1030),
.Y(n_1129)
);

CKINVDCx20_ASAP7_75t_R g1130 ( 
.A(n_1098),
.Y(n_1130)
);

INVxp33_ASAP7_75t_SL g1131 ( 
.A(n_1101),
.Y(n_1131)
);

CKINVDCx16_ASAP7_75t_R g1132 ( 
.A(n_1028),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_1089),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1093),
.B(n_1001),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_SL g1135 ( 
.A(n_1107),
.B(n_963),
.C(n_975),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1039),
.Y(n_1136)
);

NAND3xp33_ASAP7_75t_SL g1137 ( 
.A(n_1053),
.B(n_936),
.C(n_965),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1027),
.B(n_917),
.Y(n_1138)
);

NOR3xp33_ASAP7_75t_SL g1139 ( 
.A(n_1064),
.B(n_978),
.C(n_918),
.Y(n_1139)
);

INVx4_ASAP7_75t_SL g1140 ( 
.A(n_1079),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_1067),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_1045),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1066),
.A2(n_1017),
.B1(n_993),
.B2(n_946),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_1042),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_1094),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1058),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_SL g1147 ( 
.A1(n_1105),
.A2(n_1021),
.B1(n_1008),
.B2(n_958),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1045),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1075),
.Y(n_1149)
);

AND2x2_ASAP7_75t_SL g1150 ( 
.A(n_1056),
.B(n_934),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_1048),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1104),
.Y(n_1152)
);

CKINVDCx20_ASAP7_75t_R g1153 ( 
.A(n_1033),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1062),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1099),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_R g1156 ( 
.A(n_1065),
.B(n_940),
.Y(n_1156)
);

CKINVDCx14_ASAP7_75t_R g1157 ( 
.A(n_1033),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_1092),
.Y(n_1158)
);

CKINVDCx16_ASAP7_75t_R g1159 ( 
.A(n_1082),
.Y(n_1159)
);

BUFx12f_ASAP7_75t_L g1160 ( 
.A(n_1034),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1050),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1099),
.Y(n_1162)
);

NOR3xp33_ASAP7_75t_SL g1163 ( 
.A(n_1052),
.B(n_1019),
.C(n_1015),
.Y(n_1163)
);

CKINVDCx8_ASAP7_75t_R g1164 ( 
.A(n_1054),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_SL g1165 ( 
.A1(n_1085),
.A2(n_1051),
.B(n_1043),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1059),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1040),
.A2(n_1044),
.B(n_1077),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_1059),
.Y(n_1168)
);

INVxp67_ASAP7_75t_L g1169 ( 
.A(n_1086),
.Y(n_1169)
);

INVxp67_ASAP7_75t_SL g1170 ( 
.A(n_1146),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1122),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1129),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1152),
.B(n_1096),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1113),
.B(n_1120),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1112),
.Y(n_1175)
);

OR2x2_ASAP7_75t_L g1176 ( 
.A(n_1124),
.B(n_1068),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1135),
.A2(n_1080),
.B1(n_1046),
.B2(n_1047),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1145),
.Y(n_1178)
);

BUFx4f_ASAP7_75t_L g1179 ( 
.A(n_1160),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1154),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1114),
.A2(n_1060),
.B1(n_1111),
.B2(n_1078),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_1116),
.B(n_1071),
.Y(n_1182)
);

BUFx2_ASAP7_75t_SL g1183 ( 
.A(n_1125),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1123),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1123),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1136),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1149),
.Y(n_1187)
);

OR2x2_ASAP7_75t_L g1188 ( 
.A(n_1128),
.B(n_1073),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1117),
.B(n_1055),
.Y(n_1189)
);

OAI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1165),
.A2(n_1072),
.B1(n_1091),
.B2(n_1088),
.C(n_1032),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_1133),
.B(n_1109),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1138),
.B(n_1139),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_1161),
.Y(n_1193)
);

INVxp67_ASAP7_75t_L g1194 ( 
.A(n_1155),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1150),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1137),
.A2(n_1063),
.B1(n_1074),
.B2(n_1095),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1147),
.B(n_1081),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1184),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1195),
.B(n_1167),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1186),
.B(n_1132),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1170),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1175),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1189),
.B(n_1162),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1180),
.B(n_1143),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1171),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1172),
.B(n_1163),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1196),
.A2(n_1127),
.B1(n_1164),
.B2(n_1121),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1188),
.B(n_1134),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1182),
.B(n_1159),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1187),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1174),
.B(n_1156),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1202),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1198),
.Y(n_1213)
);

OR2x2_ASAP7_75t_L g1214 ( 
.A(n_1200),
.B(n_1185),
.Y(n_1214)
);

NOR2x1_ASAP7_75t_L g1215 ( 
.A(n_1209),
.B(n_1178),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1199),
.B(n_1174),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1198),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1199),
.B(n_1192),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1203),
.B(n_1173),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1201),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1205),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1208),
.B(n_1176),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1215),
.Y(n_1223)
);

AOI322xp5_ASAP7_75t_L g1224 ( 
.A1(n_1216),
.A2(n_1211),
.A3(n_1196),
.B1(n_1206),
.B2(n_1177),
.C1(n_1181),
.C2(n_1204),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1220),
.B(n_1206),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1220),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1213),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1213),
.Y(n_1228)
);

NOR4xp25_ASAP7_75t_L g1229 ( 
.A(n_1218),
.B(n_1211),
.C(n_1207),
.D(n_1181),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1222),
.B(n_1210),
.Y(n_1230)
);

OAI321xp33_ASAP7_75t_L g1231 ( 
.A1(n_1214),
.A2(n_1177),
.A3(n_1190),
.B1(n_1197),
.B2(n_1204),
.C(n_1127),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1217),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1212),
.Y(n_1233)
);

O2A1O1Ixp33_ASAP7_75t_SL g1234 ( 
.A1(n_1224),
.A2(n_1219),
.B(n_1193),
.C(n_1221),
.Y(n_1234)
);

OAI22xp33_ASAP7_75t_R g1235 ( 
.A1(n_1229),
.A2(n_1118),
.B1(n_1119),
.B2(n_1191),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1233),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1226),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_SL g1238 ( 
.A1(n_1223),
.A2(n_1157),
.B(n_1197),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1230),
.B(n_1115),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1227),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1228),
.Y(n_1241)
);

INVxp67_ASAP7_75t_SL g1242 ( 
.A(n_1235),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1236),
.B(n_1225),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1237),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1240),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1234),
.A2(n_1229),
.B(n_1231),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1242),
.B(n_1225),
.Y(n_1247)
);

AOI221xp5_ASAP7_75t_L g1248 ( 
.A1(n_1246),
.A2(n_1231),
.B1(n_1241),
.B2(n_1238),
.C(n_1239),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1243),
.B(n_1144),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1244),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1244),
.Y(n_1251)
);

O2A1O1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1245),
.A2(n_1194),
.B(n_1169),
.C(n_1232),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1250),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1251),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1252),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1255),
.B(n_1248),
.Y(n_1256)
);

XNOR2x1_ASAP7_75t_L g1257 ( 
.A(n_1253),
.B(n_1158),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1257),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1258),
.B(n_1256),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_1259),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_1259),
.Y(n_1261)
);

OR3x1_ASAP7_75t_L g1262 ( 
.A(n_1260),
.B(n_1254),
.C(n_1249),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1261),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1263),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1262),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_1264),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1265),
.A2(n_1247),
.B1(n_1130),
.B2(n_1153),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1266),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1267),
.B(n_1183),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1268),
.B(n_1131),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1269),
.A2(n_1148),
.B1(n_1140),
.B2(n_1142),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1270),
.A2(n_1140),
.B1(n_1151),
.B2(n_1179),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_SL g1273 ( 
.A1(n_1271),
.A2(n_1126),
.B1(n_1179),
.B2(n_1141),
.Y(n_1273)
);

OR2x6_ASAP7_75t_L g1274 ( 
.A(n_1273),
.B(n_1110),
.Y(n_1274)
);

AOI211xp5_ASAP7_75t_L g1275 ( 
.A1(n_1274),
.A2(n_1272),
.B(n_1168),
.C(n_1166),
.Y(n_1275)
);


endmodule