module fake_jpeg_19599_n_255 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_6),
.B(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_38),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NAND2xp33_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_40),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_3),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_22),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_20),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_49),
.B(n_30),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_22),
.B1(n_27),
.B2(n_26),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_34),
.B1(n_55),
.B2(n_44),
.Y(n_57)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_28),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_57),
.A2(n_76),
.B1(n_87),
.B2(n_88),
.Y(n_96)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_37),
.C(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_70),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_37),
.C(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_65),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_26),
.B1(n_40),
.B2(n_35),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_37),
.C(n_33),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_33),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_69),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_20),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_68),
.B(n_77),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_33),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_72),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_47),
.B1(n_27),
.B2(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_21),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_79),
.B(n_80),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_21),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_82),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_53),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_41),
.Y(n_85)
);

NAND2x1_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_19),
.Y(n_99)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_37),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_38),
.B1(n_26),
.B2(n_37),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_50),
.A2(n_37),
.B1(n_16),
.B2(n_24),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_81),
.B1(n_57),
.B2(n_38),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_101),
.B1(n_87),
.B2(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_60),
.A2(n_40),
.B1(n_35),
.B2(n_37),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_98),
.A2(n_74),
.B1(n_59),
.B2(n_86),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_106),
.B(n_112),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_60),
.A2(n_38),
.B1(n_40),
.B2(n_35),
.Y(n_101)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_17),
.A3(n_31),
.B1(n_32),
.B2(n_29),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_28),
.Y(n_133)
);

AND2x4_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_29),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_67),
.A2(n_17),
.B(n_31),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_115),
.A2(n_133),
.B1(n_111),
.B2(n_114),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_118),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_62),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_122),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_125),
.B1(n_89),
.B2(n_102),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_139),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_24),
.Y(n_122)
);

NOR2x1_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_103),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_136),
.B(n_28),
.Y(n_158)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_96),
.A2(n_105),
.B1(n_95),
.B2(n_92),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_35),
.B1(n_59),
.B2(n_64),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_127),
.A2(n_135),
.B1(n_104),
.B2(n_99),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_128),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_30),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_131),
.B(n_137),
.Y(n_144)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_66),
.B(n_17),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_138),
.B(n_89),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_58),
.B1(n_72),
.B2(n_31),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_92),
.A2(n_29),
.B(n_32),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_25),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_112),
.A2(n_32),
.B1(n_29),
.B2(n_25),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_102),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_99),
.C(n_108),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_56),
.C(n_93),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_147),
.B1(n_123),
.B2(n_120),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_132),
.B1(n_127),
.B2(n_115),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_158),
.B(n_133),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_148),
.B(n_154),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_166),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_15),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_124),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_157),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_32),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_156),
.B(n_164),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_130),
.B(n_110),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_32),
.B(n_28),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_134),
.B(n_138),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_93),
.C(n_114),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_163),
.C(n_135),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_56),
.C(n_73),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_28),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_28),
.Y(n_165)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_107),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_142),
.B1(n_160),
.B2(n_151),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_168),
.A2(n_143),
.B1(n_163),
.B2(n_159),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_182),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_170),
.A2(n_169),
.B1(n_183),
.B2(n_185),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_171),
.A2(n_158),
.B(n_161),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_145),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_174),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_149),
.Y(n_177)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_153),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_181),
.A2(n_187),
.B1(n_165),
.B2(n_18),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_116),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_116),
.C(n_123),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_185),
.C(n_186),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_184),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_139),
.C(n_107),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_110),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_153),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_198),
.B1(n_193),
.B2(n_202),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_184),
.A3(n_179),
.B1(n_168),
.B2(n_170),
.C1(n_146),
.C2(n_178),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_SL g214 ( 
.A(n_190),
.B(n_18),
.C(n_4),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_182),
.B(n_176),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_164),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_196),
.C(n_194),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_159),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_179),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_199),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_SL g200 ( 
.A(n_173),
.B(n_144),
.C(n_152),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_200),
.B(n_176),
.Y(n_212)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_203),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_211),
.Y(n_221)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_212),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_186),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_25),
.C(n_4),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_216),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_215),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_3),
.C(n_4),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_200),
.B(n_5),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_13),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_217),
.A2(n_218),
.B1(n_5),
.B2(n_6),
.Y(n_220)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_203),
.B1(n_195),
.B2(n_194),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_226),
.Y(n_230)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_204),
.A2(n_191),
.B1(n_7),
.B2(n_8),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_205),
.B(n_5),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_215),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_218),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_229)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_229),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_211),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_233),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_223),
.A2(n_210),
.B(n_206),
.Y(n_232)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_229),
.Y(n_236)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

AOI221xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_209),
.B1(n_214),
.B2(n_217),
.C(n_12),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_227),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_224),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_9),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_240),
.A2(n_235),
.B1(n_226),
.B2(n_225),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_221),
.C(n_228),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_221),
.C(n_10),
.Y(n_246)
);

AOI21x1_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_237),
.B(n_231),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_244),
.A2(n_247),
.B(n_242),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_246),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_9),
.C(n_10),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_243),
.B(n_12),
.C(n_13),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_251),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_249),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_252),
.A2(n_248),
.B(n_12),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_254),
.B(n_253),
.Y(n_255)
);


endmodule