module real_aes_1447_n_4 (n_0, n_3, n_2, n_1, n_4);
input n_0;
input n_3;
input n_2;
input n_1;
output n_4;
wire n_16;
wire n_17;
wire n_13;
wire n_18;
wire n_5;
wire n_15;
wire n_7;
wire n_8;
wire n_9;
wire n_6;
wire n_12;
wire n_14;
wire n_10;
wire n_11;
AOI32xp33_ASAP7_75t_L g4 ( .A1(n_0), .A2(n_5), .A3(n_8), .B1(n_9), .B2(n_16), .Y(n_4) );
INVx2_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_0), .B(n_15), .Y(n_14) );
INVx1_ASAP7_75t_L g7 ( .A(n_1), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_2), .Y(n_8) );
NAND2xp5_ASAP7_75t_SL g12 ( .A(n_2), .B(n_13), .Y(n_12) );
AND2x4_ASAP7_75t_L g18 ( .A(n_2), .B(n_7), .Y(n_18) );
INVxp67_ASAP7_75t_L g11 ( .A(n_3), .Y(n_11) );
INVx1_ASAP7_75t_L g15 ( .A(n_3), .Y(n_15) );
INVx1_ASAP7_75t_L g5 ( .A(n_6), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_7), .Y(n_6) );
OR2x2_ASAP7_75t_L g9 ( .A(n_10), .B(n_14), .Y(n_9) );
NOR2xp33_ASAP7_75t_L g10 ( .A(n_11), .B(n_12), .Y(n_10) );
INVx1_ASAP7_75t_L g16 ( .A(n_17), .Y(n_16) );
INVxp67_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
endmodule