module fake_jpeg_21152_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_23),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_65),
.C(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_69),
.Y(n_77)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_70),
.B(n_55),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_81),
.Y(n_90)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_78),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_63),
.B1(n_51),
.B2(n_42),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_84),
.B1(n_66),
.B2(n_40),
.Y(n_91)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_1),
.B(n_2),
.Y(n_81)
);

HAxp5_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_49),
.CON(n_84),
.SN(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_86),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_64),
.B1(n_53),
.B2(n_62),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_94),
.B1(n_87),
.B2(n_52),
.Y(n_99)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_52),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_2),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_59),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_57),
.Y(n_103)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_56),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_54),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_106),
.A2(n_112),
.B(n_44),
.Y(n_124)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_61),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_45),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_46),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_115),
.A2(n_105),
.B1(n_6),
.B2(n_9),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_118),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_50),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_119),
.B(n_123),
.Y(n_125)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_121),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_124),
.B(n_43),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_116),
.B(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_127),
.B(n_128),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_10),
.Y(n_137)
);

NAND2xp33_ASAP7_75t_SL g130 ( 
.A(n_118),
.B(n_3),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_122),
.C(n_113),
.Y(n_135)
);

AO22x1_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_38),
.B1(n_18),
.B2(n_20),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_137),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_132),
.C(n_133),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_134),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_138),
.B(n_125),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_128),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_126),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_145),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_21),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_22),
.Y(n_148)
);

BUFx24_ASAP7_75t_SL g149 ( 
.A(n_148),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_27),
.Y(n_150)
);


endmodule