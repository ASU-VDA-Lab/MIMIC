module fake_jpeg_1562_n_487 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_487);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_487;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_52),
.Y(n_141)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_53),
.Y(n_119)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_64),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_69),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_30),
.B(n_0),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_30),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_92),
.Y(n_124)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

BUFx2_ASAP7_75t_SL g101 ( 
.A(n_85),
.Y(n_101)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_17),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_47),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_98),
.B(n_103),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_38),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_52),
.A2(n_46),
.B1(n_43),
.B2(n_45),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g174 ( 
.A1(n_104),
.A2(n_90),
.B1(n_87),
.B2(n_81),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_48),
.A2(n_35),
.B1(n_45),
.B2(n_39),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_107),
.A2(n_145),
.B1(n_150),
.B2(n_44),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_66),
.A2(n_46),
.B1(n_45),
.B2(n_39),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_109),
.A2(n_138),
.B1(n_44),
.B2(n_80),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_33),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_110),
.B(n_130),
.Y(n_161)
);

INVx5_ASAP7_75t_SL g118 ( 
.A(n_68),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_118),
.B(n_142),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_79),
.B(n_33),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_50),
.B(n_23),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_56),
.A2(n_46),
.B1(n_45),
.B2(n_39),
.Y(n_138)
);

INVx5_ASAP7_75t_SL g142 ( 
.A(n_59),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_61),
.B(n_24),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_64),
.A2(n_39),
.B1(n_46),
.B2(n_43),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_65),
.Y(n_148)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_71),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_24),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_157),
.B(n_159),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_SL g238 ( 
.A1(n_158),
.A2(n_174),
.B(n_208),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_28),
.Y(n_159)
);

BUFx2_ASAP7_75t_SL g160 ( 
.A(n_118),
.Y(n_160)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_160),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_100),
.B(n_44),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_162),
.B(n_191),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_107),
.A2(n_40),
.B1(n_36),
.B2(n_82),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_164),
.A2(n_165),
.B1(n_128),
.B2(n_149),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_97),
.A2(n_112),
.B1(n_125),
.B2(n_132),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_166),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_167),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_94),
.B(n_41),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_168),
.B(n_171),
.Y(n_217)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_169),
.Y(n_245)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_99),
.Y(n_170)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_115),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_172),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_115),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_173),
.B(n_175),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_105),
.B(n_41),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_197),
.B1(n_200),
.B2(n_141),
.Y(n_211)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_183),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_119),
.Y(n_184)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_185),
.Y(n_254)
);

AOI32xp33_ASAP7_75t_L g186 ( 
.A1(n_113),
.A2(n_37),
.A3(n_28),
.B1(n_29),
.B2(n_42),
.Y(n_186)
);

AOI32xp33_ASAP7_75t_L g230 ( 
.A1(n_186),
.A2(n_1),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_230)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_127),
.Y(n_187)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_187),
.Y(n_255)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_108),
.Y(n_188)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_188),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_189),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_102),
.B(n_37),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_192),
.Y(n_213)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_135),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_95),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_193),
.B(n_195),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_SL g194 ( 
.A(n_144),
.B(n_42),
.C(n_29),
.Y(n_194)
);

NOR2x1_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_204),
.Y(n_239)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_95),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_196),
.B(n_198),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_138),
.A2(n_78),
.B1(n_42),
.B2(n_29),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_123),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_123),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_199),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_104),
.A2(n_25),
.B1(n_1),
.B2(n_3),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_207),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_119),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_111),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_129),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_206),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_140),
.B(n_0),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_101),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_146),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_142),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_146),
.B(n_3),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_114),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_117),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_211),
.A2(n_212),
.B1(n_224),
.B2(n_231),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_L g212 ( 
.A1(n_158),
.A2(n_128),
.B1(n_147),
.B2(n_129),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_218),
.A2(n_210),
.B1(n_189),
.B2(n_156),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_221),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_147),
.B1(n_121),
.B2(n_139),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_222),
.A2(n_227),
.B1(n_246),
.B2(n_252),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_162),
.A2(n_149),
.B1(n_139),
.B2(n_122),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_223),
.A2(n_260),
.B(n_257),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_163),
.A2(n_162),
.B1(n_174),
.B2(n_177),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_200),
.A2(n_121),
.B1(n_122),
.B2(n_117),
.Y(n_227)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_228),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_161),
.B(n_114),
.C(n_4),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_235),
.C(n_184),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_154),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_174),
.A2(n_17),
.B1(n_7),
.B2(n_8),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_177),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_251),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_155),
.B(n_6),
.C(n_8),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_174),
.A2(n_16),
.B1(n_8),
.B2(n_9),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_244),
.B1(n_247),
.B2(n_180),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_165),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_179),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_192),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_11),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_196),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_207),
.A2(n_12),
.B(n_13),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_208),
.B(n_167),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_169),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_211),
.A2(n_199),
.B1(n_191),
.B2(n_187),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_262),
.A2(n_274),
.B1(n_283),
.B2(n_286),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_263),
.B(n_267),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_265),
.B(n_270),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_268),
.A2(n_275),
.B(n_281),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_254),
.Y(n_269)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_269),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_170),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_224),
.B(n_201),
.Y(n_271)
);

NAND2x1_ASAP7_75t_SL g317 ( 
.A(n_271),
.B(n_278),
.Y(n_317)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_272),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_238),
.A2(n_188),
.B1(n_195),
.B2(n_172),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_239),
.A2(n_221),
.B(n_251),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_231),
.A2(n_166),
.B1(n_203),
.B2(n_185),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_276),
.A2(n_296),
.B1(n_274),
.B2(n_278),
.Y(n_339)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_249),
.Y(n_277)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_277),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_225),
.B(n_178),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_236),
.A2(n_14),
.B1(n_183),
.B2(n_212),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_279),
.A2(n_291),
.B1(n_301),
.B2(n_305),
.Y(n_307)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_280),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g281 ( 
.A(n_226),
.B(n_237),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_219),
.B(n_217),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_282),
.B(n_289),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_222),
.A2(n_227),
.B1(n_223),
.B2(n_225),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_284),
.Y(n_324)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_285),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_225),
.A2(n_226),
.B1(n_213),
.B2(n_239),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_287),
.B(n_290),
.Y(n_320)
);

XOR2x2_ASAP7_75t_L g288 ( 
.A(n_226),
.B(n_230),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_250),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_248),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_229),
.B(n_228),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_218),
.A2(n_244),
.B1(n_247),
.B2(n_233),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_233),
.B(n_259),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_292),
.B(n_295),
.Y(n_332)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_214),
.Y(n_294)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_294),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_232),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_232),
.B(n_214),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_235),
.C(n_256),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_220),
.B(n_254),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_298),
.B(n_300),
.Y(n_340)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_215),
.Y(n_299)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_243),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_300),
.B(n_278),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_258),
.A2(n_245),
.B1(n_215),
.B2(n_252),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_216),
.A2(n_260),
.B(n_242),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_302),
.A2(n_266),
.B(n_268),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_258),
.A2(n_245),
.B1(n_255),
.B2(n_253),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_303),
.A2(n_296),
.B1(n_283),
.B2(n_262),
.Y(n_326)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_255),
.Y(n_304)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_243),
.A2(n_220),
.B1(n_242),
.B2(n_253),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_280),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_306),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_261),
.A2(n_240),
.B1(n_256),
.B2(n_250),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_308),
.A2(n_328),
.B1(n_343),
.B2(n_279),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_310),
.B(n_314),
.C(n_330),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_312),
.B(n_304),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_240),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_298),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_319),
.B(n_331),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_326),
.A2(n_339),
.B1(n_318),
.B2(n_313),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_261),
.A2(n_271),
.B1(n_291),
.B2(n_273),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_297),
.B(n_263),
.C(n_281),
.Y(n_330)
);

AND2x6_ASAP7_75t_L g331 ( 
.A(n_288),
.B(n_286),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_340),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_270),
.B(n_292),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_334),
.B(n_336),
.C(n_338),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_335),
.A2(n_289),
.B(n_301),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_281),
.B(n_271),
.C(n_288),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_281),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_337),
.B(n_344),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_264),
.B(n_281),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_273),
.A2(n_265),
.B1(n_264),
.B2(n_275),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_303),
.Y(n_344)
);

OAI211xp5_ASAP7_75t_L g345 ( 
.A1(n_332),
.A2(n_267),
.B(n_336),
.C(n_322),
.Y(n_345)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_345),
.Y(n_379)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_315),
.Y(n_348)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_348),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_335),
.A2(n_302),
.B(n_287),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_349),
.A2(n_351),
.B(n_376),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_325),
.B(n_295),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_350),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_359),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_320),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_353),
.B(n_372),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_326),
.A2(n_277),
.B1(n_284),
.B2(n_293),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_354),
.A2(n_369),
.B1(n_371),
.B2(n_373),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_355),
.B(n_357),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_285),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_364),
.C(n_311),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_332),
.B(n_299),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_367),
.Y(n_387)
);

OAI21x1_ASAP7_75t_SL g359 ( 
.A1(n_323),
.A2(n_305),
.B(n_294),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_317),
.B(n_282),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_360),
.Y(n_388)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_315),
.Y(n_363)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_314),
.B(n_312),
.C(n_338),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_321),
.Y(n_365)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_365),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_340),
.Y(n_366)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_366),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_309),
.B(n_334),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_309),
.B(n_328),
.Y(n_368)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_368),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_318),
.A2(n_323),
.B1(n_343),
.B2(n_331),
.Y(n_369)
);

INVx11_ASAP7_75t_L g370 ( 
.A(n_329),
.Y(n_370)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_370),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_310),
.B(n_317),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_321),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_316),
.B(n_324),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_327),
.Y(n_384)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_341),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_368),
.A2(n_307),
.B1(n_313),
.B2(n_308),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_378),
.A2(n_393),
.B1(n_395),
.B2(n_401),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_383),
.B(n_384),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_361),
.B(n_311),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_385),
.B(n_390),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_361),
.B(n_341),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_352),
.A2(n_307),
.B1(n_342),
.B2(n_329),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_353),
.B(n_342),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_396),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_346),
.A2(n_306),
.B1(n_329),
.B2(n_349),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_362),
.B(n_372),
.C(n_364),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_399),
.B(n_403),
.C(n_390),
.Y(n_404)
);

AOI21x1_ASAP7_75t_SL g400 ( 
.A1(n_374),
.A2(n_351),
.B(n_360),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_400),
.A2(n_376),
.B(n_356),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_367),
.A2(n_347),
.B1(n_360),
.B2(n_358),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_362),
.B(n_355),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_404),
.B(n_424),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_401),
.B(n_375),
.Y(n_405)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_405),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_377),
.A2(n_347),
.B1(n_348),
.B2(n_365),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_406),
.A2(n_408),
.B1(n_409),
.B2(n_413),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_387),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_393),
.A2(n_369),
.B1(n_354),
.B2(n_359),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_389),
.Y(n_411)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_411),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_379),
.B(n_363),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_398),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_414),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_387),
.B(n_373),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_415),
.Y(n_429)
);

AOI21x1_ASAP7_75t_SL g433 ( 
.A1(n_416),
.A2(n_381),
.B(n_380),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_385),
.B(n_370),
.C(n_382),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_417),
.B(n_418),
.C(n_421),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_382),
.B(n_399),
.C(n_403),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_392),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_419),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_383),
.B(n_394),
.C(n_396),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_397),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_422),
.A2(n_425),
.B1(n_426),
.B2(n_391),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_384),
.B(n_388),
.C(n_386),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_420),
.C(n_404),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_386),
.B(n_402),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_378),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_381),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_407),
.A2(n_391),
.B1(n_381),
.B2(n_400),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_427),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_412),
.B(n_421),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_439),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_433),
.A2(n_438),
.B(n_429),
.Y(n_449)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_436),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_425),
.A2(n_380),
.B1(n_407),
.B2(n_405),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_437),
.A2(n_415),
.B1(n_411),
.B2(n_419),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_409),
.A2(n_424),
.B(n_416),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_412),
.B(n_417),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_418),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_442),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_423),
.B(n_410),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_444),
.A2(n_440),
.B1(n_428),
.B2(n_442),
.Y(n_453)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_446),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_434),
.A2(n_410),
.B1(n_435),
.B2(n_438),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_448),
.B(n_458),
.Y(n_463)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_449),
.Y(n_462)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_432),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_452),
.Y(n_459)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_430),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_453),
.B(n_454),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_429),
.A2(n_433),
.B1(n_430),
.B2(n_443),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_428),
.C(n_441),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_445),
.C(n_451),
.Y(n_466)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_444),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_457),
.B(n_445),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_431),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_455),
.B(n_458),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_466),
.Y(n_472)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_465),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_451),
.B(n_456),
.C(n_448),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_467),
.B(n_449),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_447),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_468),
.Y(n_473)
);

XNOR2x1_ASAP7_75t_L g470 ( 
.A(n_463),
.B(n_453),
.Y(n_470)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_470),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_462),
.B(n_456),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_471),
.B(n_467),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_474),
.B(n_461),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_476),
.B(n_477),
.Y(n_480)
);

NOR2xp67_ASAP7_75t_L g478 ( 
.A(n_472),
.B(n_466),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_478),
.A2(n_463),
.B(n_473),
.Y(n_479)
);

AOI221xp5_ASAP7_75t_SL g482 ( 
.A1(n_479),
.A2(n_473),
.B1(n_475),
.B2(n_460),
.C(n_469),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_480),
.Y(n_481)
);

NOR3xp33_ASAP7_75t_L g483 ( 
.A(n_481),
.B(n_482),
.C(n_459),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_483),
.A2(n_450),
.B(n_468),
.Y(n_484)
);

BUFx24_ASAP7_75t_SL g485 ( 
.A(n_484),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_485),
.B(n_470),
.Y(n_486)
);

BUFx2_ASAP7_75t_SL g487 ( 
.A(n_486),
.Y(n_487)
);


endmodule