module fake_jpeg_22193_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_9),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_44),
.B(n_22),
.Y(n_69)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_46),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_48),
.Y(n_79)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_32),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_59),
.Y(n_91)
);

CKINVDCx6p67_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_54),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_32),
.B1(n_37),
.B2(n_36),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_70),
.B1(n_73),
.B2(n_31),
.Y(n_102)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_21),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_67),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_32),
.B1(n_29),
.B2(n_28),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_68),
.A2(n_74),
.B1(n_31),
.B2(n_25),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_84),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_37),
.B1(n_36),
.B2(n_33),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_17),
.B1(n_29),
.B2(n_28),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_38),
.B1(n_22),
.B2(n_17),
.Y(n_74)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_76),
.Y(n_99)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

CKINVDCx6p67_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_35),
.B1(n_20),
.B2(n_23),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_23),
.B1(n_38),
.B2(n_43),
.Y(n_95)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_42),
.B(n_35),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_20),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_26),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_87),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_90),
.B(n_94),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_19),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_107),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_63),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_95),
.A2(n_18),
.B(n_34),
.C(n_30),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_18),
.B(n_19),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_100),
.B(n_53),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_109),
.Y(n_137)
);

AND2x4_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_19),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_105),
.B1(n_65),
.B2(n_81),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_54),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_119),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_31),
.B1(n_11),
.B2(n_13),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_19),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_19),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_65),
.B1(n_81),
.B2(n_56),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_19),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_116),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_57),
.A2(n_31),
.B1(n_18),
.B2(n_30),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_30),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_60),
.A2(n_34),
.B1(n_30),
.B2(n_25),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_82),
.B1(n_77),
.B2(n_79),
.Y(n_135)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_60),
.B(n_18),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_0),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_124),
.A2(n_24),
.B(n_103),
.Y(n_174)
);

OAI22x1_ASAP7_75t_L g186 ( 
.A1(n_126),
.A2(n_9),
.B1(n_4),
.B2(n_6),
.Y(n_186)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_130),
.B(n_138),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_97),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_131),
.B(n_133),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_56),
.B1(n_76),
.B2(n_72),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_79),
.B1(n_66),
.B2(n_71),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_139),
.B(n_144),
.Y(n_191)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_141),
.Y(n_189)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_100),
.A2(n_64),
.B1(n_62),
.B2(n_59),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_92),
.B1(n_114),
.B2(n_89),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_52),
.C(n_51),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_149),
.C(n_89),
.Y(n_169)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_157),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_13),
.Y(n_148)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_52),
.C(n_18),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_97),
.B(n_12),
.Y(n_153)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_155),
.A2(n_156),
.B1(n_92),
.B2(n_99),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_98),
.A2(n_34),
.B1(n_25),
.B2(n_24),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_178),
.Y(n_204)
);

AO22x1_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_115),
.B1(n_98),
.B2(n_108),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_159),
.A2(n_166),
.B(n_174),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_128),
.B(n_88),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_162),
.B(n_164),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_85),
.B1(n_114),
.B2(n_86),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_165),
.B(n_137),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_154),
.B(n_149),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_108),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_172),
.C(n_127),
.Y(n_197)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_34),
.B(n_18),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_168),
.A2(n_146),
.B(n_125),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_152),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_131),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_170),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_86),
.B1(n_106),
.B2(n_110),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_171),
.A2(n_180),
.B1(n_182),
.B2(n_135),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_52),
.C(n_117),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g178 ( 
.A(n_127),
.B(n_87),
.C(n_110),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_136),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_181),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_117),
.B1(n_24),
.B2(n_3),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_145),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_129),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_187),
.Y(n_219)
);

OAI22x1_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_16),
.B1(n_4),
.B2(n_6),
.Y(n_195)
);

BUFx24_ASAP7_75t_SL g187 ( 
.A(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_188),
.B(n_190),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_152),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_166),
.A2(n_130),
.B(n_138),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_213),
.B(n_218),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_193),
.B(n_197),
.C(n_221),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_195),
.A2(n_196),
.B1(n_212),
.B2(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_198),
.B(n_200),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_186),
.A2(n_151),
.B1(n_141),
.B2(n_150),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_202),
.B(n_168),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_203),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_174),
.A2(n_137),
.B(n_140),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_208),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_137),
.Y(n_207)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_146),
.Y(n_209)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_159),
.B1(n_158),
.B2(n_191),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_159),
.A2(n_123),
.B1(n_1),
.B2(n_7),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_169),
.A2(n_172),
.B1(n_180),
.B2(n_160),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_177),
.B1(n_175),
.B2(n_183),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g217 ( 
.A1(n_167),
.A2(n_4),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_182),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_162),
.B(n_123),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_123),
.C(n_10),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_210),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_224),
.B(n_225),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_211),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_226),
.A2(n_232),
.B(n_242),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_230),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_209),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_168),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_238),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_185),
.B(n_173),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_245),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_185),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_173),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_241),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_214),
.A2(n_177),
.B(n_175),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_222),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_244),
.B(n_208),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_195),
.Y(n_245)
);

OA22x2_ASAP7_75t_L g248 ( 
.A1(n_226),
.A2(n_202),
.B1(n_215),
.B2(n_212),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_248),
.A2(n_257),
.B1(n_260),
.B2(n_266),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_234),
.A2(n_241),
.B1(n_245),
.B2(n_235),
.Y(n_249)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_216),
.B1(n_206),
.B2(n_201),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_254),
.A2(n_259),
.B1(n_261),
.B2(n_267),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_237),
.Y(n_256)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_223),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_258),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_196),
.B1(n_204),
.B2(n_203),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_227),
.A2(n_194),
.B1(n_217),
.B2(n_218),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_234),
.A2(n_205),
.B1(n_192),
.B2(n_198),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_218),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_231),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_229),
.Y(n_269)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_233),
.A2(n_200),
.B1(n_221),
.B2(n_161),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_268),
.B(n_271),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_269),
.A2(n_278),
.B(n_248),
.Y(n_291)
);

XNOR2x1_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_229),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_254),
.B(n_238),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_273),
.C(n_274),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_243),
.C(n_233),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_243),
.C(n_232),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_236),
.Y(n_276)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

INVxp33_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_247),
.B(n_228),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_255),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_280),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_247),
.C(n_246),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_282),
.B(n_277),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_246),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_248),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_255),
.A2(n_161),
.B1(n_12),
.B2(n_14),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_285),
.A2(n_260),
.B1(n_267),
.B2(n_262),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_287),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_282),
.C(n_276),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_279),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_291),
.A2(n_297),
.B(n_269),
.Y(n_301)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_295),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_278),
.Y(n_295)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_263),
.C(n_251),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_284),
.B(n_281),
.Y(n_307)
);

INVx13_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_302),
.C(n_307),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_301),
.A2(n_287),
.B1(n_297),
.B2(n_292),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_273),
.C(n_274),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_283),
.B(n_272),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_248),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_268),
.C(n_275),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_288),
.C(n_293),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_303),
.A2(n_293),
.B(n_298),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_316),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_312),
.C(n_314),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_SL g312 ( 
.A(n_305),
.B(n_304),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_304),
.A2(n_294),
.B1(n_292),
.B2(n_305),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_261),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_306),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_285),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_319),
.B(n_321),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_311),
.B(n_253),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_299),
.Y(n_323)
);

AOI31xp33_ASAP7_75t_L g327 ( 
.A1(n_323),
.A2(n_299),
.A3(n_313),
.B(n_219),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_320),
.A2(n_318),
.B(n_315),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_321),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_326),
.Y(n_328)
);

AO221x1_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_327),
.B1(n_325),
.B2(n_15),
.C(n_14),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_8),
.B(n_14),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_8),
.B(n_15),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_15),
.Y(n_332)
);


endmodule