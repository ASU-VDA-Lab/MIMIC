module fake_jpeg_12533_n_452 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_452);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_452;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_18;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_56),
.Y(n_138)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_17),
.B(n_15),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_60),
.B(n_65),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_61),
.Y(n_154)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_64),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_17),
.B(n_15),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_67),
.Y(n_173)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_72),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_75),
.Y(n_177)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_77),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_26),
.B(n_13),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_78),
.B(n_95),
.Y(n_153)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_79),
.Y(n_157)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_51),
.Y(n_82)
);

CKINVDCx12_ASAP7_75t_R g156 ( 
.A(n_82),
.Y(n_156)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_84),
.Y(n_185)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_85),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_34),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_SL g160 ( 
.A(n_86),
.B(n_94),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_26),
.B(n_13),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_99),
.Y(n_128)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_88),
.Y(n_179)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_39),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_101),
.Y(n_127)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_90),
.Y(n_184)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_53),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_33),
.B(n_0),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_33),
.A2(n_1),
.B(n_3),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_96),
.B(n_4),
.Y(n_182)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_31),
.B(n_11),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_100),
.Y(n_176)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_51),
.Y(n_102)
);

INVx2_ASAP7_75t_R g174 ( 
.A(n_102),
.Y(n_174)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_38),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_107),
.Y(n_130)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_108),
.Y(n_134)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_28),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_34),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_34),
.B1(n_37),
.B2(n_29),
.Y(n_129)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_48),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_111),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_28),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_28),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_113),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_28),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_114),
.B(n_40),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_47),
.B1(n_53),
.B2(n_50),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_116),
.A2(n_122),
.B1(n_131),
.B2(n_145),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_118),
.B(n_132),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_37),
.B1(n_44),
.B2(n_43),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_119),
.A2(n_143),
.B1(n_159),
.B2(n_162),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_38),
.B1(n_44),
.B2(n_43),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_129),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_95),
.A2(n_113),
.B1(n_112),
.B2(n_84),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_61),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_86),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_135),
.B(n_140),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_102),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_54),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_142),
.B(n_171),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_59),
.A2(n_21),
.B1(n_42),
.B2(n_32),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_144),
.B(n_10),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_58),
.A2(n_21),
.B1(n_42),
.B2(n_19),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_98),
.A2(n_54),
.B1(n_46),
.B2(n_40),
.Y(n_159)
);

AO22x1_ASAP7_75t_SL g162 ( 
.A1(n_56),
.A2(n_32),
.B1(n_29),
.B2(n_27),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_64),
.A2(n_18),
.B1(n_27),
.B2(n_23),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_163),
.A2(n_167),
.B1(n_119),
.B2(n_143),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_72),
.A2(n_23),
.B1(n_20),
.B2(n_19),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_164),
.A2(n_41),
.B1(n_5),
.B2(n_6),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_67),
.A2(n_20),
.B1(n_18),
.B2(n_31),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_73),
.B(n_46),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_172),
.B(n_152),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_69),
.B(n_1),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_181),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_70),
.B(n_3),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_182),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_211)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_186),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_187),
.Y(n_249)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_189),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_134),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_190),
.B(n_209),
.Y(n_248)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_192),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_182),
.A2(n_160),
.B1(n_162),
.B2(n_122),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_193),
.A2(n_231),
.B1(n_245),
.B2(n_117),
.Y(n_250)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_194),
.Y(n_247)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_195),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_129),
.A2(n_66),
.B(n_57),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_198),
.A2(n_242),
.B(n_240),
.Y(n_277)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_199),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_200),
.A2(n_233),
.B1(n_235),
.B2(n_238),
.Y(n_280)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_138),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_201),
.Y(n_270)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_136),
.Y(n_202)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_202),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_121),
.A2(n_103),
.B1(n_76),
.B2(n_109),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_203),
.Y(n_260)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_204),
.Y(n_279)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_205),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_41),
.C(n_5),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_210),
.C(n_225),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_207),
.A2(n_189),
.B1(n_201),
.B2(n_213),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_156),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_41),
.C(n_5),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_211),
.B(n_243),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_121),
.A2(n_41),
.B1(n_8),
.B2(n_10),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_212),
.A2(n_228),
.B1(n_229),
.B2(n_241),
.Y(n_288)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_138),
.Y(n_213)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_213),
.Y(n_253)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_214),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_117),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_215),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_128),
.B(n_8),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_216),
.B(n_217),
.Y(n_263)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_219),
.B(n_220),
.Y(n_272)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_167),
.A2(n_10),
.B1(n_41),
.B2(n_145),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_221),
.A2(n_239),
.B1(n_207),
.B2(n_215),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_125),
.B(n_10),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_222),
.B(n_223),
.Y(n_282)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_153),
.B(n_174),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_224),
.B(n_226),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_130),
.B(n_149),
.C(n_148),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_163),
.B(n_141),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_166),
.A2(n_158),
.B1(n_141),
.B2(n_152),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_120),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_124),
.B(n_127),
.C(n_169),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_232),
.B(n_154),
.C(n_220),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g233 ( 
.A1(n_137),
.A2(n_146),
.B1(n_133),
.B2(n_120),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_133),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_234),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_137),
.A2(n_146),
.B1(n_155),
.B2(n_165),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_155),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_236),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_139),
.B(n_115),
.Y(n_237)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_237),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_165),
.A2(n_173),
.B1(n_170),
.B2(n_123),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_173),
.A2(n_158),
.B1(n_179),
.B2(n_147),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_126),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_240),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_126),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_244),
.Y(n_262)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_139),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_115),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_166),
.A2(n_123),
.B1(n_117),
.B2(n_175),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_250),
.A2(n_277),
.B(n_290),
.Y(n_304)
);

OA21x2_ASAP7_75t_L g251 ( 
.A1(n_227),
.A2(n_147),
.B(n_179),
.Y(n_251)
);

O2A1O1Ixp33_ASAP7_75t_SL g321 ( 
.A1(n_251),
.A2(n_269),
.B(n_271),
.C(n_284),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_218),
.A2(n_175),
.B1(n_227),
.B2(n_226),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_255),
.A2(n_257),
.B1(n_265),
.B2(n_268),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_218),
.A2(n_225),
.B1(n_198),
.B2(n_197),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_211),
.B(n_232),
.C(n_230),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_L g319 ( 
.A1(n_259),
.A2(n_267),
.B(n_291),
.C(n_279),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_266),
.A2(n_276),
.B1(n_251),
.B2(n_281),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_231),
.A2(n_208),
.B(n_196),
.C(n_191),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_200),
.A2(n_210),
.B1(n_206),
.B2(n_223),
.Y(n_268)
);

OA22x2_ASAP7_75t_L g269 ( 
.A1(n_233),
.A2(n_236),
.B1(n_214),
.B2(n_217),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_234),
.A2(n_186),
.B1(n_205),
.B2(n_199),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_274),
.A2(n_281),
.B1(n_285),
.B2(n_283),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_192),
.A2(n_194),
.B1(n_195),
.B2(n_229),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_188),
.A2(n_235),
.B1(n_238),
.B2(n_241),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_187),
.A2(n_227),
.B(n_160),
.Y(n_290)
);

XNOR2x1_ASAP7_75t_SL g325 ( 
.A(n_291),
.B(n_251),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_289),
.Y(n_292)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_292),
.Y(n_327)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_293),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_268),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_295),
.B(n_299),
.Y(n_339)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_262),
.Y(n_296)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_296),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_282),
.B(n_286),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_297),
.B(n_298),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_263),
.B(n_252),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_252),
.B(n_259),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_271),
.Y(n_300)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_300),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_274),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_301),
.B(n_302),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_256),
.B(n_267),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_247),
.Y(n_303)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_303),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_272),
.B(n_258),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_305),
.B(n_307),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_260),
.A2(n_255),
.B1(n_254),
.B2(n_251),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_306),
.A2(n_311),
.B1(n_317),
.B2(n_320),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_248),
.B(n_275),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_256),
.B(n_287),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_310),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_279),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_309),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_256),
.B(n_287),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_280),
.A2(n_250),
.B1(n_277),
.B2(n_260),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_270),
.Y(n_312)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_312),
.Y(n_351)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_253),
.Y(n_313)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_313),
.Y(n_353)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_247),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_314),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_278),
.B(n_254),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_324),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_265),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_316),
.A2(n_318),
.B(n_319),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_280),
.A2(n_288),
.B1(n_291),
.B2(n_285),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_261),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_321),
.A2(n_322),
.B1(n_326),
.B2(n_246),
.Y(n_341)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_261),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_323),
.A2(n_269),
.B1(n_273),
.B2(n_284),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_273),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_299),
.Y(n_336)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_304),
.A2(n_283),
.B(n_264),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_330),
.A2(n_341),
.B(n_344),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_304),
.A2(n_249),
.B(n_289),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_331),
.A2(n_334),
.B(n_338),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_332),
.A2(n_301),
.B1(n_324),
.B2(n_315),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_308),
.A2(n_310),
.B(n_302),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_336),
.B(n_316),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_311),
.A2(n_246),
.B(n_269),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_325),
.A2(n_269),
.B(n_249),
.Y(n_344)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_313),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_346),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_298),
.B(n_295),
.C(n_294),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_348),
.B(n_317),
.C(n_316),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_343),
.B(n_305),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_365),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_294),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_359),
.C(n_361),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_321),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_368),
.Y(n_392)
);

XNOR2x1_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_342),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_348),
.B(n_293),
.C(n_296),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_362),
.A2(n_367),
.B1(n_335),
.B2(n_334),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_319),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_347),
.C(n_375),
.Y(n_385)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_340),
.Y(n_364)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_364),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_350),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_332),
.A2(n_350),
.B1(n_335),
.B2(n_328),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_340),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_349),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_371),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_333),
.A2(n_297),
.B1(n_318),
.B2(n_323),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_370),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_349),
.Y(n_371)
);

NOR2x1_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_303),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_372),
.B(n_373),
.Y(n_391)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_329),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_328),
.B(n_314),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_374),
.B(n_375),
.Y(n_377)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_329),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_339),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_381),
.C(n_383),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_358),
.B(n_361),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_360),
.A2(n_333),
.B(n_345),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_382),
.B(n_384),
.Y(n_395)
);

MAJx2_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_356),
.C(n_357),
.Y(n_401)
);

AOI211xp5_ASAP7_75t_L g386 ( 
.A1(n_365),
.A2(n_345),
.B(n_331),
.C(n_341),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_386),
.A2(n_394),
.B1(n_371),
.B2(n_369),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_344),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_359),
.C(n_373),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_356),
.A2(n_338),
.B(n_321),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_390),
.B(n_393),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_360),
.A2(n_327),
.B(n_337),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_357),
.A2(n_352),
.B1(n_351),
.B2(n_353),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_379),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_389),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_399),
.B(n_407),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_381),
.B(n_367),
.C(n_374),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_400),
.B(n_402),
.C(n_406),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_388),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_376),
.B(n_362),
.C(n_364),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_380),
.Y(n_403)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_403),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_352),
.C(n_366),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_409),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_405),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_368),
.C(n_372),
.Y(n_406)
);

BUFx5_ASAP7_75t_L g407 ( 
.A(n_387),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_378),
.A2(n_343),
.B1(n_351),
.B2(n_327),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_384),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_353),
.C(n_337),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_410),
.B(n_419),
.C(n_398),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_395),
.A2(n_378),
.B1(n_390),
.B2(n_377),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_411),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_396),
.A2(n_377),
.B1(n_394),
.B2(n_391),
.Y(n_412)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_412),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_415),
.B(n_397),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_402),
.B(n_397),
.C(n_400),
.Y(n_419)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_420),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_423),
.B(n_425),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_419),
.B(n_401),
.C(n_406),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_426),
.B(n_427),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_417),
.B(n_393),
.C(n_382),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_414),
.B(n_407),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_428),
.B(n_429),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_392),
.C(n_377),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_422),
.A2(n_416),
.B1(n_413),
.B2(n_418),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_326),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_428),
.B(n_416),
.Y(n_432)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_432),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_421),
.A2(n_411),
.B1(n_386),
.B2(n_387),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_434),
.A2(n_392),
.B(n_346),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_424),
.A2(n_392),
.B(n_415),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_435),
.B(n_320),
.Y(n_440)
);

XNOR2x1_ASAP7_75t_SL g437 ( 
.A(n_433),
.B(n_410),
.Y(n_437)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_437),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_438),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_439),
.B(n_440),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_436),
.B(n_322),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_442),
.B(n_431),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_446),
.B(n_440),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_443),
.B(n_441),
.Y(n_447)
);

AOI321xp33_ASAP7_75t_L g449 ( 
.A1(n_447),
.A2(n_448),
.A3(n_444),
.B1(n_445),
.B2(n_435),
.C(n_434),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_449),
.B(n_312),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_450),
.B(n_292),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_451),
.B(n_312),
.Y(n_452)
);


endmodule