module fake_jpeg_7213_n_343 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_9),
.B(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_10),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_0),
.C(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_38),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_51),
.B(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_27),
.B1(n_24),
.B2(n_21),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_53),
.A2(n_26),
.B1(n_23),
.B2(n_17),
.Y(n_95)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_63),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_27),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_70),
.A2(n_73),
.B1(n_86),
.B2(n_89),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_76),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_64),
.A2(n_27),
.B1(n_24),
.B2(n_21),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

BUFx4f_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_49),
.B1(n_46),
.B2(n_42),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_90),
.B1(n_52),
.B2(n_50),
.Y(n_103)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_49),
.B1(n_46),
.B2(n_42),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_77),
.A2(n_57),
.B1(n_23),
.B2(n_33),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_80),
.Y(n_117)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_62),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_81),
.B(n_91),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

CKINVDCx9p33_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_57),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_22),
.Y(n_131)
);

NAND2x1_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_22),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_23),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_51),
.A2(n_24),
.B1(n_21),
.B2(n_26),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_24),
.B1(n_26),
.B2(n_36),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_28),
.B1(n_17),
.B2(n_35),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_96),
.B(n_97),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_44),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_32),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_98),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_100),
.B(n_95),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_32),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_41),
.C(n_62),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_104),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_103),
.A2(n_109),
.B1(n_86),
.B2(n_72),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_41),
.C(n_66),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_114),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_112),
.A2(n_118),
.B1(n_35),
.B2(n_33),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_100),
.A2(n_88),
.B1(n_77),
.B2(n_91),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_120),
.B1(n_79),
.B2(n_70),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g115 ( 
.A(n_77),
.B(n_0),
.Y(n_115)
);

AOI32xp33_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_85),
.A3(n_22),
.B1(n_20),
.B2(n_30),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_60),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_116),
.B(n_131),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_55),
.B1(n_28),
.B2(n_33),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_94),
.A2(n_55),
.B1(n_28),
.B2(n_35),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_123),
.Y(n_137)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_115),
.B1(n_103),
.B2(n_113),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_139),
.B1(n_149),
.B2(n_80),
.Y(n_176)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_133),
.B(n_134),
.Y(n_192)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_15),
.Y(n_136)
);

XNOR2x1_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_140),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_93),
.Y(n_138)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_70),
.B1(n_71),
.B2(n_81),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_13),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_142),
.A2(n_156),
.B1(n_19),
.B2(n_76),
.Y(n_186)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_144),
.A2(n_129),
.B(n_18),
.Y(n_183)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_146),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_14),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_151),
.Y(n_172)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_60),
.B1(n_72),
.B2(n_41),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_9),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_153),
.Y(n_193)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_106),
.Y(n_181)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_122),
.B1(n_84),
.B2(n_121),
.Y(n_162)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_162),
.A2(n_176),
.B1(n_186),
.B2(n_160),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_104),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_168),
.C(n_178),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_102),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_166),
.B(n_182),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_135),
.C(n_159),
.Y(n_168)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_147),
.A2(n_116),
.A3(n_127),
.B1(n_120),
.B2(n_126),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_30),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_151),
.A2(n_119),
.B1(n_126),
.B2(n_105),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_184),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_132),
.A2(n_105),
.B1(n_19),
.B2(n_18),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_175),
.Y(n_223)
);

O2A1O1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_129),
.B(n_20),
.C(n_130),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_179),
.B1(n_122),
.B2(n_154),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_39),
.Y(n_178)
);

OAI22x1_ASAP7_75t_SL g179 ( 
.A1(n_132),
.A2(n_30),
.B1(n_34),
.B2(n_20),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_39),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_189),
.C(n_178),
.Y(n_211)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

AOI21x1_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_22),
.B(n_34),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_183),
.B(n_155),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_78),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_139),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_30),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_135),
.B(n_45),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_140),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_15),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_195),
.B(n_198),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_141),
.Y(n_197)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

AND2x6_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_136),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_205),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_132),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_211),
.C(n_221),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_201),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_176),
.A2(n_150),
.B1(n_149),
.B2(n_158),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_202),
.A2(n_212),
.B1(n_217),
.B2(n_223),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_193),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_203),
.B(n_214),
.Y(n_244)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_206),
.Y(n_247)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_163),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_210),
.Y(n_251)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_179),
.A2(n_122),
.B1(n_143),
.B2(n_157),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_153),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_222),
.Y(n_231)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_190),
.B(n_175),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_168),
.B(n_45),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_187),
.Y(n_224)
);

NOR3xp33_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_82),
.C(n_74),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_78),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

OAI221xp5_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_188),
.B1(n_166),
.B2(n_189),
.C(n_180),
.Y(n_230)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_213),
.B1(n_220),
.B2(n_199),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_161),
.Y(n_233)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_215),
.Y(n_235)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_237),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_191),
.Y(n_238)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_238),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_202),
.A2(n_191),
.B1(n_167),
.B2(n_106),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_240),
.A2(n_223),
.B1(n_213),
.B2(n_212),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g241 ( 
.A1(n_217),
.A2(n_78),
.B(n_99),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_250),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_34),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_242),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_209),
.A2(n_69),
.B1(n_99),
.B2(n_74),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_82),
.B1(n_69),
.B2(n_34),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_196),
.B(n_69),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_196),
.Y(n_254)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_249),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_271),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_244),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_253),
.A2(n_272),
.B(n_226),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_243),
.Y(n_275)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_208),
.Y(n_261)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_229),
.B(n_236),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_262),
.B(n_229),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_221),
.C(n_213),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_270),
.C(n_242),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_246),
.B(n_195),
.Y(n_266)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_228),
.A2(n_6),
.B1(n_14),
.B2(n_11),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_269),
.A2(n_251),
.B1(n_231),
.B2(n_232),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_22),
.C(n_1),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_246),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_234),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_276),
.C(n_277),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_238),
.B(n_241),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_280),
.A2(n_239),
.B1(n_241),
.B2(n_263),
.Y(n_298)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_238),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_284),
.C(n_286),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_240),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_237),
.Y(n_286)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_227),
.Y(n_289)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_258),
.A2(n_247),
.B1(n_231),
.B2(n_239),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_263),
.B1(n_245),
.B2(n_233),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_274),
.A2(n_260),
.B1(n_269),
.B2(n_259),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_291),
.A2(n_292),
.B1(n_8),
.B2(n_6),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_273),
.A2(n_259),
.B1(n_264),
.B2(n_255),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_285),
.A2(n_271),
.B1(n_272),
.B2(n_253),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_293),
.A2(n_278),
.B(n_284),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_233),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_305),
.C(n_0),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_286),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_300),
.A2(n_306),
.B1(n_2),
.B2(n_3),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_11),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_277),
.B(n_252),
.C(n_268),
.Y(n_305)
);

OAI321xp33_ASAP7_75t_L g306 ( 
.A1(n_280),
.A2(n_11),
.A3(n_8),
.B1(n_7),
.B2(n_6),
.C(n_4),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_287),
.B(n_282),
.Y(n_307)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_308),
.B(n_309),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_303),
.B(n_290),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_311),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_275),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_314),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_8),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_316),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_1),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_2),
.Y(n_324)
);

A2O1A1Ixp33_ASAP7_75t_SL g320 ( 
.A1(n_318),
.A2(n_295),
.B(n_294),
.C(n_4),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_320),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_310),
.A2(n_300),
.B(n_305),
.Y(n_322)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_322),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_324),
.B(n_2),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_297),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_308),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_328),
.Y(n_334)
);

AOI31xp67_ASAP7_75t_L g330 ( 
.A1(n_320),
.A2(n_302),
.A3(n_316),
.B(n_313),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_R g335 ( 
.A(n_330),
.B(n_331),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_311),
.C(n_296),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_332),
.A2(n_333),
.B1(n_321),
.B2(n_326),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_329),
.B(n_319),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_335),
.Y(n_338)
);

AOI21x1_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_320),
.B(n_296),
.Y(n_339)
);

NAND3xp33_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_327),
.C(n_334),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_3),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_3),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_5),
.Y(n_343)
);


endmodule