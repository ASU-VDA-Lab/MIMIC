module fake_aes_4638_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx16_ASAP7_75t_R g11 ( .A(n_10), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
CKINVDCx8_ASAP7_75t_R g15 ( .A(n_4), .Y(n_15) );
BUFx2_ASAP7_75t_L g16 ( .A(n_11), .Y(n_16) );
BUFx3_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_18), .B(n_13), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
OR2x2_ASAP7_75t_L g24 ( .A(n_22), .B(n_16), .Y(n_24) );
OAI322xp33_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_18), .A3(n_21), .B1(n_20), .B2(n_13), .C1(n_15), .C2(n_19), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
AOI221xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_13), .B1(n_15), .B2(n_2), .C(n_3), .Y(n_27) );
NAND2xp33_ASAP7_75t_SL g28 ( .A(n_26), .B(n_13), .Y(n_28) );
BUFx2_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
NOR2xp33_ASAP7_75t_R g30 ( .A(n_27), .B(n_0), .Y(n_30) );
OAI22x1_ASAP7_75t_SL g31 ( .A1(n_30), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
AOI22xp5_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_1), .B1(n_3), .B2(n_5), .Y(n_33) );
AOI322xp5_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_5), .A3(n_6), .B1(n_9), .B2(n_32), .C1(n_12), .C2(n_27), .Y(n_34) );
endmodule