module fake_netlist_1_2512_n_1160 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1160);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1160;
wire n_791;
wire n_707;
wire n_663;
wire n_513;
wire n_361;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_1122;
wire n_779;
wire n_993;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_345;
wire n_360;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_638;
wire n_563;
wire n_830;
wire n_517;
wire n_560;
wire n_955;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1011;
wire n_1025;
wire n_1132;
wire n_1155;
wire n_1101;
wire n_1159;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_844;
wire n_818;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_1138;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_1154;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_771;
wire n_696;
wire n_735;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_1046;
wire n_935;
wire n_460;
wire n_950;
wire n_478;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_880;
wire n_799;
wire n_1089;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_1157;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_1125;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_1060;
wire n_1133;
wire n_908;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_1042;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_912;
wire n_947;
wire n_924;
wire n_1043;
wire n_378;
wire n_582;
wire n_1141;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_994;
wire n_930;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_919;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_1146;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_257;
wire n_992;
wire n_1127;
wire n_269;
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_66), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_139), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_8), .Y(n_251) );
CKINVDCx16_ASAP7_75t_R g252 ( .A(n_232), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_159), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_228), .Y(n_254) );
NOR2xp67_ASAP7_75t_L g255 ( .A(n_39), .B(n_127), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_192), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_35), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_121), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_73), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_236), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_209), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_9), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_208), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_12), .Y(n_264) );
OR2x2_ASAP7_75t_L g265 ( .A(n_96), .B(n_166), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_78), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_229), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_92), .Y(n_268) );
NOR2xp67_ASAP7_75t_L g269 ( .A(n_22), .B(n_155), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_49), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_43), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_84), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_21), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_239), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_194), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_221), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_11), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_74), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_212), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_191), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_72), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_108), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_225), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_226), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g285 ( .A(n_149), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_144), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_126), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_97), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_136), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_214), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_147), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_113), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_248), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g294 ( .A(n_243), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_26), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g296 ( .A(n_160), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_211), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_227), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_98), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_151), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_138), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_235), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_40), .Y(n_303) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_182), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_242), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_128), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_150), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_137), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_76), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_247), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_176), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_86), .Y(n_312) );
CKINVDCx16_ASAP7_75t_R g313 ( .A(n_237), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_201), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_153), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_219), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_50), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_195), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_115), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_188), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_60), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_106), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_104), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_154), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_241), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_123), .Y(n_326) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_133), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_53), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_167), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_103), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_132), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_67), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_102), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_37), .Y(n_334) );
BUFx10_ASAP7_75t_L g335 ( .A(n_63), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_131), .Y(n_336) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_69), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_100), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_56), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_55), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_179), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_183), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_10), .Y(n_343) );
BUFx2_ASAP7_75t_SL g344 ( .A(n_173), .Y(n_344) );
CKINVDCx16_ASAP7_75t_R g345 ( .A(n_99), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_218), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_68), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_78), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_105), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_118), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_184), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_0), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_31), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_120), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_20), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_2), .Y(n_356) );
INVxp67_ASAP7_75t_L g357 ( .A(n_119), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_246), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_80), .B(n_206), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_145), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_217), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_204), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_171), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_7), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_117), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_77), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_186), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_111), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_101), .Y(n_369) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_88), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_107), .Y(n_371) );
NOR2xp67_ASAP7_75t_L g372 ( .A(n_180), .B(n_12), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_234), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_172), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_134), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_222), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_87), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_33), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_202), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_233), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_36), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_143), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_57), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_112), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_156), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_177), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_276), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_316), .Y(n_388) );
AND2x2_ASAP7_75t_SL g389 ( .A(n_265), .B(n_245), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_328), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_276), .B(n_1), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_276), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_328), .Y(n_393) );
INVx3_ASAP7_75t_L g394 ( .A(n_370), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_343), .B(n_1), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_250), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_396) );
BUFx3_ASAP7_75t_L g397 ( .A(n_316), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_331), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_283), .B(n_3), .Y(n_399) );
INVx3_ASAP7_75t_L g400 ( .A(n_370), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_343), .Y(n_401) );
INVx5_ASAP7_75t_L g402 ( .A(n_331), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_250), .A2(n_6), .B1(n_4), .B2(n_5), .Y(n_403) );
AND2x4_ASAP7_75t_L g404 ( .A(n_352), .B(n_5), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_352), .Y(n_405) );
BUFx2_ASAP7_75t_L g406 ( .A(n_268), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_252), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_313), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_264), .A2(n_8), .B1(n_6), .B2(n_7), .Y(n_409) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_331), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_295), .B(n_9), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_331), .Y(n_412) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_333), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_345), .B(n_10), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_300), .B(n_11), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_342), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_261), .B(n_13), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_275), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_333), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_253), .Y(n_420) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_333), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_264), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_275), .A2(n_15), .B1(n_13), .B2(n_14), .Y(n_423) );
INVx6_ASAP7_75t_L g424 ( .A(n_402), .Y(n_424) );
BUFx3_ASAP7_75t_L g425 ( .A(n_388), .Y(n_425) );
AND2x6_ASAP7_75t_L g426 ( .A(n_417), .B(n_258), .Y(n_426) );
BUFx8_ASAP7_75t_SL g427 ( .A(n_406), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_416), .B(n_323), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_420), .B(n_261), .Y(n_429) );
INVx3_ASAP7_75t_L g430 ( .A(n_417), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_395), .A2(n_259), .B1(n_262), .B2(n_257), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_417), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_410), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_417), .B(n_270), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_422), .Y(n_435) );
NAND3xp33_ASAP7_75t_L g436 ( .A(n_417), .B(n_386), .C(n_263), .Y(n_436) );
INVx4_ASAP7_75t_L g437 ( .A(n_395), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_420), .B(n_280), .Y(n_438) );
BUFx10_ASAP7_75t_L g439 ( .A(n_389), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_416), .B(n_280), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_389), .B(n_290), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_409), .A2(n_251), .B1(n_317), .B2(n_249), .Y(n_442) );
INVx5_ASAP7_75t_L g443 ( .A(n_410), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_422), .B(n_335), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_389), .B(n_290), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_410), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_395), .A2(n_272), .B1(n_273), .B2(n_271), .Y(n_447) );
INVx2_ASAP7_75t_SL g448 ( .A(n_388), .Y(n_448) );
INVx2_ASAP7_75t_SL g449 ( .A(n_388), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_395), .A2(n_278), .B1(n_281), .B2(n_277), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_395), .Y(n_451) );
AND2x2_ASAP7_75t_SL g452 ( .A(n_404), .B(n_359), .Y(n_452) );
OAI22xp33_ASAP7_75t_SL g453 ( .A1(n_396), .A2(n_266), .B1(n_377), .B2(n_309), .Y(n_453) );
BUFx3_ASAP7_75t_L g454 ( .A(n_397), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_404), .B(n_291), .Y(n_455) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_410), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_404), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_412), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_404), .Y(n_459) );
AND3x2_ASAP7_75t_L g460 ( .A(n_406), .B(n_357), .C(n_312), .Y(n_460) );
AND2x6_ASAP7_75t_L g461 ( .A(n_411), .B(n_260), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_414), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_394), .Y(n_463) );
INVxp33_ASAP7_75t_SL g464 ( .A(n_407), .Y(n_464) );
INVxp33_ASAP7_75t_L g465 ( .A(n_414), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_412), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_412), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_411), .B(n_335), .Y(n_468) );
INVxp33_ASAP7_75t_L g469 ( .A(n_414), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_394), .Y(n_470) );
OAI22xp33_ASAP7_75t_L g471 ( .A1(n_462), .A2(n_409), .B1(n_403), .B2(n_396), .Y(n_471) );
OR2x6_ASAP7_75t_L g472 ( .A(n_444), .B(n_403), .Y(n_472) );
NAND2x1p5_ASAP7_75t_L g473 ( .A(n_435), .B(n_411), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_428), .B(n_468), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_425), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_435), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_425), .Y(n_477) );
BUFx5_ASAP7_75t_L g478 ( .A(n_426), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_455), .A2(n_397), .B(n_391), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_441), .A2(n_445), .B1(n_468), .B2(n_461), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_462), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_430), .A2(n_399), .B(n_415), .C(n_393), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_428), .B(n_415), .Y(n_483) );
INVx4_ASAP7_75t_L g484 ( .A(n_437), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_452), .B(n_267), .Y(n_485) );
BUFx3_ASAP7_75t_L g486 ( .A(n_427), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_437), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_444), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_440), .B(n_444), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_437), .B(n_408), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_465), .B(n_418), .Y(n_491) );
AND2x2_ASAP7_75t_SL g492 ( .A(n_452), .B(n_370), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_426), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_441), .A2(n_393), .B1(n_401), .B2(n_390), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_445), .A2(n_401), .B1(n_405), .B2(n_390), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_434), .B(n_405), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_452), .B(n_308), .Y(n_497) );
NOR2xp67_ASAP7_75t_L g498 ( .A(n_442), .B(n_423), .Y(n_498) );
NOR2x1p5_ASAP7_75t_L g499 ( .A(n_464), .B(n_266), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_426), .B(n_308), .Y(n_500) );
OR2x6_ASAP7_75t_L g501 ( .A(n_442), .B(n_423), .Y(n_501) );
AND2x2_ASAP7_75t_SL g502 ( .A(n_434), .B(n_370), .Y(n_502) );
NAND2x1p5_ASAP7_75t_L g503 ( .A(n_451), .B(n_303), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_457), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_439), .A2(n_251), .B1(n_317), .B2(n_249), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_426), .B(n_375), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_426), .B(n_379), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_426), .B(n_380), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_426), .B(n_380), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_426), .B(n_385), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_434), .B(n_385), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_457), .A2(n_334), .B1(n_339), .B2(n_332), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_434), .B(n_254), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_469), .B(n_335), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_434), .B(n_256), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_461), .A2(n_294), .B1(n_296), .B2(n_285), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_461), .B(n_286), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_461), .B(n_432), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_461), .B(n_288), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_461), .B(n_289), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_430), .B(n_451), .Y(n_521) );
AND2x6_ASAP7_75t_SL g522 ( .A(n_453), .B(n_340), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_451), .Y(n_523) );
INVx8_ASAP7_75t_L g524 ( .A(n_461), .Y(n_524) );
BUFx3_ASAP7_75t_L g525 ( .A(n_451), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_431), .B(n_299), .Y(n_526) );
NOR2xp67_ASAP7_75t_L g527 ( .A(n_436), .B(n_377), .Y(n_527) );
INVx2_ASAP7_75t_SL g528 ( .A(n_460), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_453), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_430), .B(n_310), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_451), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_430), .B(n_311), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_448), .A2(n_307), .B(n_297), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_447), .B(n_322), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_459), .A2(n_355), .B1(n_364), .B2(n_348), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_447), .B(n_329), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_459), .A2(n_378), .B1(n_381), .B2(n_366), .Y(n_537) );
INVxp67_ASAP7_75t_L g538 ( .A(n_429), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_450), .B(n_338), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_439), .A2(n_296), .B1(n_304), .B2(n_294), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_454), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_459), .A2(n_383), .B1(n_282), .B2(n_284), .Y(n_542) );
BUFx3_ASAP7_75t_L g543 ( .A(n_454), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_438), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_436), .B(n_354), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_439), .A2(n_318), .B1(n_319), .B2(n_304), .Y(n_546) );
NOR2x2_ASAP7_75t_L g547 ( .A(n_460), .B(n_337), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_449), .B(n_358), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_449), .B(n_362), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_439), .B(n_365), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_488), .B(n_439), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_476), .A2(n_319), .B1(n_327), .B2(n_318), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_521), .A2(n_470), .B(n_463), .Y(n_553) );
O2A1O1Ixp33_ASAP7_75t_L g554 ( .A1(n_471), .A2(n_337), .B(n_279), .C(n_292), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_538), .B(n_327), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_516), .A2(n_330), .B1(n_369), .B2(n_336), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_481), .Y(n_557) );
OAI21xp33_ASAP7_75t_SL g558 ( .A1(n_502), .A2(n_269), .B(n_255), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_492), .A2(n_336), .B1(n_369), .B2(n_330), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_487), .Y(n_560) );
INVx3_ASAP7_75t_L g561 ( .A(n_484), .Y(n_561) );
INVx5_ASAP7_75t_L g562 ( .A(n_524), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_481), .B(n_321), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_523), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_483), .B(n_489), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_531), .Y(n_566) );
AO32x1_ASAP7_75t_L g567 ( .A1(n_475), .A2(n_398), .A3(n_392), .B1(n_387), .B2(n_298), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_502), .A2(n_353), .B1(n_356), .B2(n_347), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_530), .A2(n_532), .B(n_485), .Y(n_569) );
A2O1A1Ixp33_ASAP7_75t_L g570 ( .A1(n_504), .A2(n_496), .B(n_482), .C(n_498), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_474), .A2(n_446), .B(n_433), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_501), .B(n_14), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_488), .B(n_274), .Y(n_573) );
INVx4_ASAP7_75t_L g574 ( .A(n_524), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_472), .B(n_372), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_492), .A2(n_293), .B1(n_301), .B2(n_287), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_473), .B(n_374), .Y(n_577) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_524), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_518), .A2(n_466), .B(n_458), .Y(n_579) );
O2A1O1Ixp33_ASAP7_75t_L g580 ( .A1(n_471), .A2(n_306), .B(n_314), .C(n_302), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_514), .B(n_305), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_491), .B(n_367), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_533), .A2(n_467), .B(n_320), .Y(n_583) );
NOR2xp67_ASAP7_75t_L g584 ( .A(n_528), .B(n_15), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_497), .B(n_315), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_513), .A2(n_467), .B(n_325), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g587 ( .A1(n_479), .A2(n_326), .B(n_324), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_478), .B(n_341), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_515), .A2(n_467), .B(n_351), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_480), .A2(n_472), .B1(n_503), .B2(n_540), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_472), .A2(n_360), .B1(n_363), .B2(n_349), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_511), .A2(n_371), .B(n_368), .Y(n_592) );
AO22x1_ASAP7_75t_L g593 ( .A1(n_486), .A2(n_376), .B1(n_382), .B2(n_373), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_499), .B(n_384), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_505), .B(n_16), .Y(n_595) );
O2A1O1Ixp33_ASAP7_75t_L g596 ( .A1(n_526), .A2(n_346), .B(n_350), .C(n_307), .Y(n_596) );
A2O1A1Ixp33_ASAP7_75t_L g597 ( .A1(n_496), .A2(n_350), .B(n_346), .C(n_394), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_544), .Y(n_598) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_484), .Y(n_599) );
A2O1A1Ixp33_ASAP7_75t_L g600 ( .A1(n_527), .A2(n_400), .B(n_344), .C(n_361), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_546), .B(n_16), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_493), .A2(n_400), .B1(n_361), .B2(n_333), .Y(n_602) );
BUFx12f_ASAP7_75t_L g603 ( .A(n_522), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_490), .B(n_17), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_512), .B(n_400), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_529), .B(n_17), .Y(n_606) );
A2O1A1Ixp33_ASAP7_75t_L g607 ( .A1(n_494), .A2(n_412), .B(n_419), .C(n_413), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_512), .B(n_18), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_534), .B(n_18), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_535), .B(n_19), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_493), .B(n_402), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_537), .B(n_19), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_542), .A2(n_402), .B1(n_424), .B2(n_413), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_536), .B(n_20), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_539), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_537), .B(n_21), .Y(n_616) );
BUFx8_ASAP7_75t_L g617 ( .A(n_547), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_500), .B(n_412), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_L g619 ( .A1(n_494), .A2(n_419), .B(n_421), .C(n_413), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_517), .A2(n_443), .B(n_456), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_SL g621 ( .A1(n_495), .A2(n_424), .B(n_456), .C(n_419), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_495), .A2(n_424), .B1(n_419), .B2(n_421), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_519), .A2(n_443), .B(n_456), .Y(n_623) );
INVx5_ASAP7_75t_L g624 ( .A(n_543), .Y(n_624) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_477), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g626 ( .A1(n_545), .A2(n_421), .B(n_419), .C(n_443), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_520), .B(n_23), .Y(n_627) );
INVx4_ASAP7_75t_L g628 ( .A(n_541), .Y(n_628) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_506), .A2(n_443), .B(n_421), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_507), .B(n_456), .Y(n_630) );
NOR2xp33_ASAP7_75t_SL g631 ( .A(n_508), .B(n_24), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_548), .A2(n_456), .B(n_94), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_549), .Y(n_633) );
NAND2x1p5_ASAP7_75t_L g634 ( .A(n_509), .B(n_25), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_510), .B(n_25), .Y(n_635) );
AOI21x1_ASAP7_75t_L g636 ( .A1(n_550), .A2(n_456), .B(n_95), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_525), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_538), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_538), .B(n_26), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_476), .B(n_27), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_488), .B(n_28), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_538), .B(n_28), .Y(n_642) );
OAI321xp33_ASAP7_75t_L g643 ( .A1(n_471), .A2(n_29), .A3(n_30), .B1(n_31), .B2(n_32), .C(n_33), .Y(n_643) );
INVx1_ASAP7_75t_SL g644 ( .A(n_476), .Y(n_644) );
AOI21xp33_ASAP7_75t_L g645 ( .A1(n_476), .A2(n_30), .B(n_32), .Y(n_645) );
CKINVDCx5p33_ASAP7_75t_R g646 ( .A(n_486), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_488), .B(n_34), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_476), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_488), .B(n_35), .Y(n_649) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_476), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_488), .B(n_37), .Y(n_651) );
BUFx2_ASAP7_75t_L g652 ( .A(n_476), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_538), .B(n_38), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_538), .B(n_38), .Y(n_654) );
OR2x6_ASAP7_75t_L g655 ( .A(n_524), .B(n_41), .Y(n_655) );
BUFx10_ASAP7_75t_L g656 ( .A(n_476), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_L g657 ( .A1(n_471), .A2(n_41), .B(n_42), .C(n_43), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_538), .B(n_42), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_488), .B(n_44), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_SL g660 ( .A1(n_482), .A2(n_152), .B(n_244), .C(n_240), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_538), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_565), .A2(n_110), .B(n_109), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_638), .B(n_44), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_569), .A2(n_116), .B(n_114), .Y(n_664) );
NAND3xp33_ASAP7_75t_L g665 ( .A(n_558), .B(n_45), .C(n_46), .Y(n_665) );
OAI21x1_ASAP7_75t_SL g666 ( .A1(n_590), .A2(n_45), .B(n_46), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_570), .A2(n_47), .B(n_48), .C(n_49), .Y(n_667) );
BUFx3_ASAP7_75t_L g668 ( .A(n_656), .Y(n_668) );
OAI21x1_ASAP7_75t_L g669 ( .A1(n_632), .A2(n_124), .B(n_122), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_557), .B(n_47), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_615), .B(n_48), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_572), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_555), .B(n_50), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_652), .Y(n_674) );
INVx2_ASAP7_75t_SL g675 ( .A(n_656), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_630), .A2(n_165), .B(n_238), .Y(n_676) );
INVx1_ASAP7_75t_SL g677 ( .A(n_644), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g678 ( .A1(n_580), .A2(n_51), .B(n_52), .Y(n_678) );
AO31x2_ASAP7_75t_L g679 ( .A1(n_607), .A2(n_52), .A3(n_53), .B(n_54), .Y(n_679) );
NAND2xp33_ASAP7_75t_SL g680 ( .A(n_574), .B(n_54), .Y(n_680) );
A2O1A1Ixp33_ASAP7_75t_L g681 ( .A1(n_609), .A2(n_55), .B(n_56), .C(n_57), .Y(n_681) );
AOI221x1_ASAP7_75t_L g682 ( .A1(n_575), .A2(n_58), .B1(n_59), .B2(n_60), .C(n_61), .Y(n_682) );
A2O1A1Ixp33_ASAP7_75t_L g683 ( .A1(n_614), .A2(n_62), .B(n_63), .C(n_64), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_633), .B(n_62), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_564), .Y(n_685) );
AO31x2_ASAP7_75t_L g686 ( .A1(n_619), .A2(n_64), .A3(n_65), .B(n_66), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_563), .B(n_65), .Y(n_687) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_648), .Y(n_688) );
INVx3_ASAP7_75t_L g689 ( .A(n_599), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_566), .Y(n_690) );
A2O1A1Ixp33_ASAP7_75t_L g691 ( .A1(n_604), .A2(n_68), .B(n_69), .C(n_70), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_650), .B(n_70), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_646), .Y(n_693) );
OAI22x1_ASAP7_75t_L g694 ( .A1(n_552), .A2(n_71), .B1(n_72), .B2(n_73), .Y(n_694) );
AO31x2_ASAP7_75t_L g695 ( .A1(n_626), .A2(n_74), .A3(n_75), .B(n_76), .Y(n_695) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_620), .A2(n_175), .B(n_231), .Y(n_696) );
AO31x2_ASAP7_75t_L g697 ( .A1(n_597), .A2(n_622), .A3(n_591), .B(n_627), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_623), .A2(n_174), .B(n_230), .Y(n_698) );
OAI21xp5_ASAP7_75t_L g699 ( .A1(n_587), .A2(n_75), .B(n_77), .Y(n_699) );
AND2x4_ASAP7_75t_L g700 ( .A(n_562), .B(n_79), .Y(n_700) );
NOR2xp67_ASAP7_75t_SL g701 ( .A(n_562), .B(n_79), .Y(n_701) );
AO31x2_ASAP7_75t_L g702 ( .A1(n_583), .A2(n_80), .A3(n_81), .B(n_82), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_655), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_703) );
BUFx3_ASAP7_75t_L g704 ( .A(n_617), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_601), .B(n_83), .Y(n_705) );
OAI21xp5_ASAP7_75t_L g706 ( .A1(n_586), .A2(n_84), .B(n_85), .Y(n_706) );
AND2x4_ASAP7_75t_L g707 ( .A(n_562), .B(n_85), .Y(n_707) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_655), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_559), .B(n_89), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_574), .B(n_90), .Y(n_710) );
AND2x4_ASAP7_75t_L g711 ( .A(n_578), .B(n_90), .Y(n_711) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_655), .Y(n_712) );
AO31x2_ASAP7_75t_L g713 ( .A1(n_635), .A2(n_91), .A3(n_93), .B(n_125), .Y(n_713) );
INVxp67_ASAP7_75t_L g714 ( .A(n_640), .Y(n_714) );
O2A1O1Ixp33_ASAP7_75t_L g715 ( .A1(n_554), .A2(n_129), .B(n_130), .C(n_135), .Y(n_715) );
OAI21xp5_ASAP7_75t_L g716 ( .A1(n_589), .A2(n_140), .B(n_141), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_575), .A2(n_142), .B1(n_146), .B2(n_148), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_598), .B(n_551), .Y(n_718) );
CKINVDCx11_ASAP7_75t_R g719 ( .A(n_603), .Y(n_719) );
BUFx10_ASAP7_75t_L g720 ( .A(n_641), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_618), .A2(n_157), .B(n_158), .Y(n_721) );
O2A1O1Ixp33_ASAP7_75t_L g722 ( .A1(n_657), .A2(n_161), .B(n_162), .C(n_163), .Y(n_722) );
O2A1O1Ixp33_ASAP7_75t_SL g723 ( .A1(n_621), .A2(n_164), .B(n_168), .C(n_169), .Y(n_723) );
AOI222xp33_ASAP7_75t_L g724 ( .A1(n_617), .A2(n_170), .B1(n_178), .B2(n_181), .C1(n_185), .C2(n_187), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_634), .A2(n_189), .B1(n_190), .B2(n_193), .Y(n_725) );
CKINVDCx16_ASAP7_75t_R g726 ( .A(n_595), .Y(n_726) );
OAI21x1_ASAP7_75t_SL g727 ( .A1(n_639), .A2(n_196), .B(n_197), .Y(n_727) );
OAI21x1_ASAP7_75t_L g728 ( .A1(n_579), .A2(n_198), .B(n_199), .Y(n_728) );
NAND2x1p5_ASAP7_75t_L g729 ( .A(n_578), .B(n_200), .Y(n_729) );
AOI221xp5_ASAP7_75t_SL g730 ( .A1(n_592), .A2(n_203), .B1(n_205), .B2(n_207), .C(n_210), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_585), .B(n_213), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_573), .B(n_215), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g733 ( .A1(n_629), .A2(n_216), .B(n_220), .Y(n_733) );
BUFx3_ASAP7_75t_L g734 ( .A(n_624), .Y(n_734) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_553), .A2(n_223), .B(n_224), .Y(n_735) );
INVx2_ASAP7_75t_SL g736 ( .A(n_594), .Y(n_736) );
INVxp67_ASAP7_75t_L g737 ( .A(n_647), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_582), .B(n_581), .Y(n_738) );
BUFx4f_ASAP7_75t_SL g739 ( .A(n_594), .Y(n_739) );
AND2x6_ASAP7_75t_L g740 ( .A(n_561), .B(n_637), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_642), .Y(n_741) );
AOI21xp33_ASAP7_75t_SL g742 ( .A1(n_606), .A2(n_593), .B(n_659), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_588), .A2(n_611), .B(n_660), .Y(n_743) );
INVx2_ASAP7_75t_SL g744 ( .A(n_624), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_653), .Y(n_745) );
AO31x2_ASAP7_75t_L g746 ( .A1(n_576), .A2(n_651), .A3(n_649), .B(n_613), .Y(n_746) );
A2O1A1Ixp33_ASAP7_75t_L g747 ( .A1(n_596), .A2(n_616), .B(n_612), .C(n_610), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_654), .Y(n_748) );
AO32x2_ASAP7_75t_L g749 ( .A1(n_628), .A2(n_567), .A3(n_602), .B1(n_643), .B2(n_568), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_608), .B(n_658), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_605), .Y(n_751) );
A2O1A1Ixp33_ASAP7_75t_L g752 ( .A1(n_645), .A2(n_631), .B(n_584), .C(n_577), .Y(n_752) );
INVx5_ASAP7_75t_L g753 ( .A(n_625), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_567), .A2(n_625), .B(n_628), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_625), .A2(n_498), .B1(n_501), .B2(n_471), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_565), .B(n_538), .Y(n_756) );
OAI22x1_ASAP7_75t_L g757 ( .A1(n_552), .A2(n_540), .B1(n_546), .B2(n_516), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_646), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_565), .B(n_538), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_555), .B(n_472), .Y(n_760) );
INVxp67_ASAP7_75t_SL g761 ( .A(n_552), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_638), .Y(n_762) );
A2O1A1Ixp33_ASAP7_75t_L g763 ( .A1(n_570), .A2(n_614), .B(n_609), .C(n_569), .Y(n_763) );
INVx3_ASAP7_75t_SL g764 ( .A(n_646), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_565), .B(n_538), .Y(n_765) );
INVx3_ASAP7_75t_L g766 ( .A(n_599), .Y(n_766) );
OR2x2_ASAP7_75t_L g767 ( .A(n_552), .B(n_476), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_646), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_565), .B(n_538), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_555), .B(n_472), .Y(n_770) );
O2A1O1Ixp33_ASAP7_75t_SL g771 ( .A1(n_570), .A2(n_626), .B(n_600), .C(n_619), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g772 ( .A(n_646), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_638), .Y(n_773) );
AO31x2_ASAP7_75t_L g774 ( .A1(n_607), .A2(n_619), .A3(n_570), .B(n_626), .Y(n_774) );
AND2x4_ASAP7_75t_L g775 ( .A(n_638), .B(n_661), .Y(n_775) );
AO21x2_ASAP7_75t_L g776 ( .A1(n_621), .A2(n_636), .B(n_619), .Y(n_776) );
OAI21xp33_ASAP7_75t_SL g777 ( .A1(n_655), .A2(n_445), .B(n_441), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_565), .A2(n_569), .B(n_571), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_638), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_556), .A2(n_501), .B1(n_498), .B2(n_472), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_565), .B(n_538), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_638), .B(n_462), .Y(n_782) );
OAI21xp5_ASAP7_75t_L g783 ( .A1(n_570), .A2(n_569), .B(n_480), .Y(n_783) );
AOI221x1_ASAP7_75t_L g784 ( .A1(n_575), .A2(n_619), .B1(n_607), .B2(n_591), .C(n_600), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_555), .B(n_472), .Y(n_785) );
A2O1A1Ixp33_ASAP7_75t_L g786 ( .A1(n_570), .A2(n_614), .B(n_609), .C(n_569), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_565), .A2(n_569), .B(n_571), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_560), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_560), .Y(n_789) );
OA22x2_ASAP7_75t_L g790 ( .A1(n_552), .A2(n_501), .B1(n_546), .B2(n_540), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_638), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g792 ( .A1(n_763), .A2(n_786), .B(n_778), .Y(n_792) );
INVx2_ASAP7_75t_SL g793 ( .A(n_668), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g794 ( .A1(n_750), .A2(n_783), .B(n_771), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_756), .Y(n_795) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_677), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_783), .A2(n_731), .B(n_747), .Y(n_797) );
INVx1_ASAP7_75t_SL g798 ( .A(n_677), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_759), .Y(n_799) );
BUFx2_ASAP7_75t_L g800 ( .A(n_674), .Y(n_800) );
INVx4_ASAP7_75t_L g801 ( .A(n_764), .Y(n_801) );
AO31x2_ASAP7_75t_L g802 ( .A1(n_784), .A2(n_667), .A3(n_682), .B(n_751), .Y(n_802) );
BUFx6f_ASAP7_75t_L g803 ( .A(n_753), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_726), .B(n_761), .Y(n_804) );
OAI221xp5_ASAP7_75t_L g805 ( .A1(n_780), .A2(n_755), .B1(n_765), .B2(n_769), .C(n_781), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_755), .B(n_718), .Y(n_806) );
AOI21xp33_ASAP7_75t_L g807 ( .A1(n_777), .A2(n_715), .B(n_722), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_718), .B(n_788), .Y(n_808) );
AO31x2_ASAP7_75t_L g809 ( .A1(n_743), .A2(n_664), .A3(n_752), .B(n_725), .Y(n_809) );
A2O1A1Ixp33_ASAP7_75t_L g810 ( .A1(n_777), .A2(n_748), .B(n_741), .C(n_745), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_762), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_773), .Y(n_812) );
AO21x2_ASAP7_75t_L g813 ( .A1(n_776), .A2(n_727), .B(n_733), .Y(n_813) );
NAND2x1p5_ASAP7_75t_L g814 ( .A(n_700), .B(n_707), .Y(n_814) );
OA21x2_ASAP7_75t_L g815 ( .A1(n_730), .A2(n_733), .B(n_716), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_779), .Y(n_816) );
OA21x2_ASAP7_75t_L g817 ( .A1(n_716), .A2(n_728), .B(n_669), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_791), .Y(n_818) );
BUFx2_ASAP7_75t_L g819 ( .A(n_693), .Y(n_819) );
AOI21xp5_ASAP7_75t_L g820 ( .A1(n_731), .A2(n_776), .B(n_723), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_684), .Y(n_821) );
AND2x4_ASAP7_75t_L g822 ( .A(n_775), .B(n_675), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_775), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_685), .Y(n_824) );
A2O1A1Ixp33_ASAP7_75t_L g825 ( .A1(n_678), .A2(n_699), .B(n_680), .C(n_742), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_782), .B(n_790), .Y(n_826) );
BUFx5_ASAP7_75t_L g827 ( .A(n_740), .Y(n_827) );
NAND2x1p5_ASAP7_75t_L g828 ( .A(n_700), .B(n_707), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_690), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_789), .B(n_672), .Y(n_830) );
OAI21xp5_ASAP7_75t_L g831 ( .A1(n_671), .A2(n_699), .B(n_678), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_671), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_663), .Y(n_833) );
AO31x2_ASAP7_75t_L g834 ( .A1(n_725), .A2(n_681), .A3(n_683), .B(n_691), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_767), .B(n_705), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_670), .Y(n_836) );
BUFx6f_ASAP7_75t_L g837 ( .A(n_753), .Y(n_837) );
INVx4_ASAP7_75t_L g838 ( .A(n_739), .Y(n_838) );
AND2x4_ASAP7_75t_L g839 ( .A(n_710), .B(n_753), .Y(n_839) );
INVx3_ASAP7_75t_L g840 ( .A(n_734), .Y(n_840) );
OAI21xp5_ASAP7_75t_L g841 ( .A1(n_706), .A2(n_737), .B(n_665), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_738), .B(n_770), .Y(n_842) );
BUFx4f_ASAP7_75t_SL g843 ( .A(n_704), .Y(n_843) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_688), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_703), .Y(n_845) );
OAI21xp5_ASAP7_75t_L g846 ( .A1(n_706), .A2(n_665), .B(n_676), .Y(n_846) );
AND2x2_ASAP7_75t_L g847 ( .A(n_760), .B(n_785), .Y(n_847) );
OA21x2_ASAP7_75t_L g848 ( .A1(n_696), .A2(n_698), .B(n_735), .Y(n_848) );
CKINVDCx5p33_ASAP7_75t_R g849 ( .A(n_719), .Y(n_849) );
INVx1_ASAP7_75t_SL g850 ( .A(n_710), .Y(n_850) );
OAI21xp5_ASAP7_75t_L g851 ( .A1(n_662), .A2(n_721), .B(n_687), .Y(n_851) );
OA21x2_ASAP7_75t_L g852 ( .A1(n_666), .A2(n_717), .B(n_732), .Y(n_852) );
BUFx2_ASAP7_75t_L g853 ( .A(n_758), .Y(n_853) );
OAI21x1_ASAP7_75t_L g854 ( .A1(n_729), .A2(n_766), .B(n_689), .Y(n_854) );
BUFx8_ASAP7_75t_L g855 ( .A(n_736), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g856 ( .A(n_742), .B(n_714), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_757), .B(n_709), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_746), .B(n_712), .Y(n_858) );
OR2x6_ASAP7_75t_L g859 ( .A(n_708), .B(n_711), .Y(n_859) );
INVx2_ASAP7_75t_SL g860 ( .A(n_772), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_692), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_694), .Y(n_862) );
AOI22xp33_ASAP7_75t_SL g863 ( .A1(n_711), .A2(n_673), .B1(n_720), .B2(n_768), .Y(n_863) );
AOI21xp5_ASAP7_75t_L g864 ( .A1(n_744), .A2(n_724), .B(n_774), .Y(n_864) );
CKINVDCx12_ASAP7_75t_R g865 ( .A(n_701), .Y(n_865) );
AO21x2_ASAP7_75t_L g866 ( .A1(n_749), .A2(n_697), .B(n_713), .Y(n_866) );
OAI21x1_ASAP7_75t_L g867 ( .A1(n_697), .A2(n_740), .B(n_749), .Y(n_867) );
AOI21xp5_ASAP7_75t_L g868 ( .A1(n_746), .A2(n_679), .B(n_686), .Y(n_868) );
AOI21x1_ASAP7_75t_L g869 ( .A1(n_713), .A2(n_695), .B(n_686), .Y(n_869) );
OAI21x1_ASAP7_75t_SL g870 ( .A1(n_695), .A2(n_699), .B(n_733), .Y(n_870) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_695), .Y(n_871) );
OR2x2_ASAP7_75t_L g872 ( .A(n_702), .B(n_756), .Y(n_872) );
BUFx2_ASAP7_75t_L g873 ( .A(n_677), .Y(n_873) );
AOI21xp33_ASAP7_75t_SL g874 ( .A1(n_764), .A2(n_471), .B(n_442), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_756), .B(n_759), .Y(n_875) );
INVxp67_ASAP7_75t_SL g876 ( .A(n_756), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_756), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_756), .Y(n_878) );
AOI21xp5_ASAP7_75t_L g879 ( .A1(n_763), .A2(n_786), .B(n_778), .Y(n_879) );
A2O1A1Ixp33_ASAP7_75t_L g880 ( .A1(n_777), .A2(n_750), .B(n_715), .C(n_558), .Y(n_880) );
AOI21xp5_ASAP7_75t_L g881 ( .A1(n_763), .A2(n_786), .B(n_778), .Y(n_881) );
OR3x4_ASAP7_75t_SL g882 ( .A(n_719), .B(n_617), .C(n_761), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g883 ( .A(n_726), .B(n_761), .Y(n_883) );
OAI21xp5_ASAP7_75t_L g884 ( .A1(n_778), .A2(n_570), .B(n_787), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_756), .B(n_759), .Y(n_885) );
INVx3_ASAP7_75t_L g886 ( .A(n_734), .Y(n_886) );
AND2x4_ASAP7_75t_L g887 ( .A(n_756), .B(n_759), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_756), .B(n_759), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_756), .B(n_759), .Y(n_889) );
INVx2_ASAP7_75t_L g890 ( .A(n_756), .Y(n_890) );
INVxp33_ASAP7_75t_L g891 ( .A(n_756), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_756), .B(n_759), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_756), .B(n_759), .Y(n_893) );
AOI21xp5_ASAP7_75t_L g894 ( .A1(n_763), .A2(n_786), .B(n_778), .Y(n_894) );
AO31x2_ASAP7_75t_L g895 ( .A1(n_763), .A2(n_786), .A3(n_784), .B(n_754), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_756), .B(n_759), .Y(n_896) );
AO21x2_ASAP7_75t_L g897 ( .A1(n_820), .A2(n_870), .B(n_879), .Y(n_897) );
AOI222xp33_ASAP7_75t_L g898 ( .A1(n_887), .A2(n_893), .B1(n_888), .B2(n_896), .C1(n_875), .C2(n_889), .Y(n_898) );
INVx2_ASAP7_75t_SL g899 ( .A(n_855), .Y(n_899) );
BUFx3_ASAP7_75t_L g900 ( .A(n_803), .Y(n_900) );
OAI21xp5_ASAP7_75t_L g901 ( .A1(n_825), .A2(n_810), .B(n_880), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_876), .B(n_877), .Y(n_902) );
AND2x2_ASAP7_75t_L g903 ( .A(n_878), .B(n_890), .Y(n_903) );
AND2x4_ASAP7_75t_L g904 ( .A(n_806), .B(n_884), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_887), .B(n_795), .Y(n_905) );
INVx3_ASAP7_75t_L g906 ( .A(n_803), .Y(n_906) );
INVx3_ASAP7_75t_L g907 ( .A(n_837), .Y(n_907) );
INVx3_ASAP7_75t_L g908 ( .A(n_837), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_872), .Y(n_909) );
HB1xp67_ASAP7_75t_L g910 ( .A(n_844), .Y(n_910) );
AO21x2_ASAP7_75t_L g911 ( .A1(n_881), .A2(n_894), .B(n_792), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_871), .Y(n_912) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_796), .Y(n_913) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_843), .Y(n_914) );
BUFx6f_ASAP7_75t_L g915 ( .A(n_837), .Y(n_915) );
AND2x4_ASAP7_75t_L g916 ( .A(n_806), .B(n_884), .Y(n_916) );
OR2x2_ASAP7_75t_L g917 ( .A(n_875), .B(n_885), .Y(n_917) );
INVx1_ASAP7_75t_SL g918 ( .A(n_819), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_832), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_891), .B(n_874), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_808), .Y(n_921) );
INVx2_ASAP7_75t_SL g922 ( .A(n_855), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_885), .B(n_889), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_808), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_821), .Y(n_925) );
AND2x2_ASAP7_75t_L g926 ( .A(n_892), .B(n_896), .Y(n_926) );
OR2x6_ASAP7_75t_L g927 ( .A(n_864), .B(n_814), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_845), .Y(n_928) );
BUFx3_ASAP7_75t_L g929 ( .A(n_839), .Y(n_929) );
NAND2x1p5_ASAP7_75t_L g930 ( .A(n_839), .B(n_850), .Y(n_930) );
BUFx2_ASAP7_75t_L g931 ( .A(n_814), .Y(n_931) );
INVx5_ASAP7_75t_L g932 ( .A(n_859), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_869), .Y(n_933) );
OA21x2_ASAP7_75t_L g934 ( .A1(n_868), .A2(n_867), .B(n_797), .Y(n_934) );
BUFx2_ASAP7_75t_L g935 ( .A(n_828), .Y(n_935) );
BUFx2_ASAP7_75t_L g936 ( .A(n_859), .Y(n_936) );
HB1xp67_ASAP7_75t_L g937 ( .A(n_873), .Y(n_937) );
INVxp67_ASAP7_75t_L g938 ( .A(n_892), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_850), .A2(n_805), .B1(n_859), .B2(n_863), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_805), .A2(n_826), .B1(n_883), .B2(n_804), .Y(n_940) );
OR2x2_ASAP7_75t_L g941 ( .A(n_857), .B(n_858), .Y(n_941) );
AND3x1_ASAP7_75t_L g942 ( .A(n_856), .B(n_862), .C(n_857), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_858), .Y(n_943) );
HB1xp67_ASAP7_75t_L g944 ( .A(n_800), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_847), .B(n_835), .Y(n_945) );
INVx1_ASAP7_75t_SL g946 ( .A(n_853), .Y(n_946) );
INVx3_ASAP7_75t_L g947 ( .A(n_827), .Y(n_947) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_798), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_824), .B(n_829), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_811), .Y(n_950) );
OA21x2_ASAP7_75t_L g951 ( .A1(n_846), .A2(n_831), .B(n_794), .Y(n_951) );
INVxp67_ASAP7_75t_SL g952 ( .A(n_830), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_812), .Y(n_953) );
OR2x2_ASAP7_75t_L g954 ( .A(n_842), .B(n_798), .Y(n_954) );
HB1xp67_ASAP7_75t_L g955 ( .A(n_799), .Y(n_955) );
AO21x2_ASAP7_75t_L g956 ( .A1(n_831), .A2(n_807), .B(n_866), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_842), .B(n_816), .Y(n_957) );
BUFx3_ASAP7_75t_L g958 ( .A(n_822), .Y(n_958) );
INVx2_ASAP7_75t_SL g959 ( .A(n_793), .Y(n_959) );
OR2x6_ASAP7_75t_L g960 ( .A(n_841), .B(n_854), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_818), .B(n_833), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_841), .B(n_830), .Y(n_962) );
OR2x2_ASAP7_75t_L g963 ( .A(n_836), .B(n_866), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_895), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_823), .B(n_861), .Y(n_965) );
INVxp67_ASAP7_75t_L g966 ( .A(n_860), .Y(n_966) );
AND2x2_ASAP7_75t_L g967 ( .A(n_904), .B(n_813), .Y(n_967) );
OR2x2_ASAP7_75t_L g968 ( .A(n_941), .B(n_802), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_928), .B(n_802), .Y(n_969) );
OR2x2_ASAP7_75t_L g970 ( .A(n_941), .B(n_802), .Y(n_970) );
INVx1_ASAP7_75t_SL g971 ( .A(n_902), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_904), .B(n_809), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_904), .B(n_809), .Y(n_973) );
AND2x4_ASAP7_75t_L g974 ( .A(n_927), .B(n_809), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_962), .B(n_834), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_904), .B(n_815), .Y(n_976) );
INVx4_ASAP7_75t_L g977 ( .A(n_932), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_928), .B(n_834), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_916), .B(n_815), .Y(n_979) );
AND2x4_ASAP7_75t_SL g980 ( .A(n_902), .B(n_886), .Y(n_980) );
BUFx2_ASAP7_75t_L g981 ( .A(n_927), .Y(n_981) );
HB1xp67_ASAP7_75t_L g982 ( .A(n_948), .Y(n_982) );
NOR2xp67_ASAP7_75t_R g983 ( .A(n_932), .B(n_801), .Y(n_983) );
HB1xp67_ASAP7_75t_L g984 ( .A(n_912), .Y(n_984) );
HB1xp67_ASAP7_75t_L g985 ( .A(n_912), .Y(n_985) );
INVx4_ASAP7_75t_R g986 ( .A(n_899), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_963), .Y(n_987) );
HB1xp67_ASAP7_75t_L g988 ( .A(n_909), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_916), .B(n_817), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_964), .B(n_852), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_909), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_943), .Y(n_992) );
OR2x2_ASAP7_75t_L g993 ( .A(n_954), .B(n_886), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_933), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_926), .B(n_840), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_926), .B(n_840), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_898), .A2(n_851), .B1(n_801), .B2(n_827), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_939), .A2(n_838), .B1(n_848), .B2(n_882), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_921), .B(n_865), .Y(n_999) );
AND2x4_ASAP7_75t_L g1000 ( .A(n_927), .B(n_947), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_924), .B(n_849), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_957), .B(n_903), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_957), .B(n_903), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_925), .Y(n_1004) );
INVx2_ASAP7_75t_SL g1005 ( .A(n_932), .Y(n_1005) );
INVx2_ASAP7_75t_SL g1006 ( .A(n_932), .Y(n_1006) );
NOR2xp33_ASAP7_75t_L g1007 ( .A(n_966), .B(n_918), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_994), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_972), .B(n_973), .Y(n_1009) );
NOR2xp33_ASAP7_75t_L g1010 ( .A(n_1001), .B(n_899), .Y(n_1010) );
INVxp67_ASAP7_75t_SL g1011 ( .A(n_982), .Y(n_1011) );
NAND2xp5_ASAP7_75t_SL g1012 ( .A(n_998), .B(n_932), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1004), .Y(n_1013) );
AND2x6_ASAP7_75t_SL g1014 ( .A(n_1007), .B(n_914), .Y(n_1014) );
INVxp67_ASAP7_75t_SL g1015 ( .A(n_982), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_1002), .B(n_952), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_978), .B(n_956), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_1002), .B(n_955), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_978), .B(n_956), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_969), .B(n_956), .Y(n_1020) );
OR2x2_ASAP7_75t_L g1021 ( .A(n_971), .B(n_913), .Y(n_1021) );
NAND2x1p5_ASAP7_75t_L g1022 ( .A(n_977), .B(n_932), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_969), .B(n_951), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_976), .B(n_951), .Y(n_1024) );
INVxp67_ASAP7_75t_L g1025 ( .A(n_1001), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_976), .B(n_951), .Y(n_1026) );
HB1xp67_ASAP7_75t_L g1027 ( .A(n_971), .Y(n_1027) );
OR2x2_ASAP7_75t_L g1028 ( .A(n_968), .B(n_951), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_997), .A2(n_940), .B1(n_920), .B2(n_945), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_1003), .B(n_938), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_976), .B(n_897), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_968), .B(n_917), .Y(n_1032) );
INVx4_ASAP7_75t_L g1033 ( .A(n_977), .Y(n_1033) );
OR2x2_ASAP7_75t_L g1034 ( .A(n_970), .B(n_917), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_979), .B(n_897), .Y(n_1035) );
INVx5_ASAP7_75t_SL g1036 ( .A(n_983), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_979), .B(n_897), .Y(n_1037) );
OR2x2_ASAP7_75t_L g1038 ( .A(n_975), .B(n_937), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_988), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1003), .Y(n_1040) );
INVx1_ASAP7_75t_SL g1041 ( .A(n_980), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_967), .B(n_934), .Y(n_1042) );
AND2x4_ASAP7_75t_L g1043 ( .A(n_1000), .B(n_960), .Y(n_1043) );
AND2x4_ASAP7_75t_L g1044 ( .A(n_1000), .B(n_960), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_995), .B(n_953), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_995), .B(n_953), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1040), .B(n_991), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_1045), .B(n_991), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1011), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_1009), .B(n_967), .Y(n_1050) );
INVx4_ASAP7_75t_L g1051 ( .A(n_1033), .Y(n_1051) );
INVx2_ASAP7_75t_SL g1052 ( .A(n_1033), .Y(n_1052) );
AND2x4_ASAP7_75t_L g1053 ( .A(n_1043), .B(n_974), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1009), .B(n_989), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1008), .Y(n_1055) );
AOI22xp5_ASAP7_75t_L g1056 ( .A1(n_1029), .A2(n_942), .B1(n_999), .B2(n_905), .Y(n_1056) );
OR2x2_ASAP7_75t_L g1057 ( .A(n_1038), .B(n_987), .Y(n_1057) );
INVxp67_ASAP7_75t_L g1058 ( .A(n_1027), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_1031), .B(n_989), .Y(n_1059) );
HB1xp67_ASAP7_75t_L g1060 ( .A(n_1021), .Y(n_1060) );
OR2x2_ASAP7_75t_L g1061 ( .A(n_1038), .B(n_987), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1008), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1046), .B(n_984), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_1018), .B(n_984), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_1030), .B(n_985), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1015), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1016), .B(n_985), .Y(n_1067) );
AOI221xp5_ASAP7_75t_L g1068 ( .A1(n_1025), .A2(n_942), .B1(n_910), .B2(n_901), .C(n_945), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_1031), .B(n_989), .Y(n_1069) );
BUFx2_ASAP7_75t_L g1070 ( .A(n_1033), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_1035), .B(n_1037), .Y(n_1071) );
NAND2x1p5_ASAP7_75t_L g1072 ( .A(n_1041), .B(n_977), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_1039), .B(n_992), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1035), .B(n_990), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1037), .B(n_1024), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1024), .B(n_990), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1013), .Y(n_1077) );
INVx1_ASAP7_75t_SL g1078 ( .A(n_1014), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1075), .B(n_1042), .Y(n_1079) );
INVxp67_ASAP7_75t_L g1080 ( .A(n_1060), .Y(n_1080) );
NAND2xp5_ASAP7_75t_SL g1081 ( .A(n_1051), .B(n_1036), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1057), .Y(n_1082) );
HB1xp67_ASAP7_75t_L g1083 ( .A(n_1058), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1057), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1071), .B(n_1026), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1071), .B(n_1023), .Y(n_1086) );
INVxp33_ASAP7_75t_L g1087 ( .A(n_1070), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1061), .Y(n_1088) );
OAI22xp33_ASAP7_75t_R g1089 ( .A1(n_1078), .A2(n_946), .B1(n_1010), .B2(n_922), .Y(n_1089) );
AOI21xp5_ASAP7_75t_L g1090 ( .A1(n_1051), .A2(n_1012), .B(n_983), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1054), .B(n_1026), .Y(n_1091) );
OR2x6_ASAP7_75t_L g1092 ( .A(n_1051), .B(n_1022), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1074), .B(n_1017), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1061), .Y(n_1094) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_1056), .A2(n_1036), .B1(n_980), .B2(n_1022), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1049), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1066), .Y(n_1097) );
OR2x2_ASAP7_75t_L g1098 ( .A(n_1076), .B(n_1028), .Y(n_1098) );
NAND2x1p5_ASAP7_75t_L g1099 ( .A(n_1052), .B(n_977), .Y(n_1099) );
INVxp67_ASAP7_75t_L g1100 ( .A(n_1064), .Y(n_1100) );
INVxp67_ASAP7_75t_L g1101 ( .A(n_1065), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1055), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1054), .B(n_1020), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_1067), .B(n_1019), .Y(n_1104) );
INVx1_ASAP7_75t_SL g1105 ( .A(n_1063), .Y(n_1105) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1098), .Y(n_1106) );
NAND2xp5_ASAP7_75t_SL g1107 ( .A(n_1090), .B(n_1036), .Y(n_1107) );
OAI21xp33_ASAP7_75t_SL g1108 ( .A1(n_1081), .A2(n_1068), .B(n_1050), .Y(n_1108) );
NAND3xp33_ASAP7_75t_SL g1109 ( .A(n_1087), .B(n_1022), .C(n_1072), .Y(n_1109) );
AOI21xp33_ASAP7_75t_SL g1110 ( .A1(n_1081), .A2(n_1072), .B(n_922), .Y(n_1110) );
OAI22xp33_ASAP7_75t_L g1111 ( .A1(n_1092), .A2(n_1034), .B1(n_1032), .B2(n_981), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1102), .Y(n_1112) );
AOI22xp5_ASAP7_75t_L g1113 ( .A1(n_1089), .A2(n_1053), .B1(n_1059), .B2(n_1069), .Y(n_1113) );
NOR2xp33_ASAP7_75t_L g1114 ( .A(n_1101), .B(n_1047), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_1092), .A2(n_1036), .B1(n_1053), .B2(n_980), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_1100), .A2(n_996), .B1(n_905), .B2(n_1032), .Y(n_1116) );
O2A1O1Ixp33_ASAP7_75t_SL g1117 ( .A1(n_1087), .A2(n_986), .B(n_944), .C(n_1006), .Y(n_1117) );
OAI221xp5_ASAP7_75t_L g1118 ( .A1(n_1095), .A2(n_1048), .B1(n_959), .B2(n_1073), .C(n_1077), .Y(n_1118) );
HB1xp67_ASAP7_75t_L g1119 ( .A(n_1080), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1096), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1079), .B(n_1050), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_1108), .A2(n_1044), .B1(n_1043), .B2(n_1105), .Y(n_1122) );
AOI21xp5_ASAP7_75t_L g1123 ( .A1(n_1107), .A2(n_1099), .B(n_1104), .Y(n_1123) );
O2A1O1Ixp33_ASAP7_75t_L g1124 ( .A1(n_1107), .A2(n_1083), .B(n_1097), .C(n_959), .Y(n_1124) );
AOI22xp5_ASAP7_75t_L g1125 ( .A1(n_1113), .A2(n_1118), .B1(n_1111), .B2(n_1114), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_1111), .A2(n_1044), .B1(n_1043), .B2(n_1084), .Y(n_1126) );
AOI221xp5_ASAP7_75t_L g1127 ( .A1(n_1114), .A2(n_1082), .B1(n_1094), .B2(n_1088), .C(n_1103), .Y(n_1127) );
NOR3xp33_ASAP7_75t_L g1128 ( .A(n_1109), .B(n_923), .C(n_961), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1119), .B(n_1103), .Y(n_1129) );
AOI21xp5_ASAP7_75t_L g1130 ( .A1(n_1117), .A2(n_1099), .B(n_1086), .Y(n_1130) );
AOI211xp5_ASAP7_75t_L g1131 ( .A1(n_1110), .A2(n_1028), .B(n_1034), .C(n_1044), .Y(n_1131) );
NOR3x1_ASAP7_75t_L g1132 ( .A(n_1115), .B(n_986), .C(n_1093), .Y(n_1132) );
AOI221xp5_ASAP7_75t_L g1133 ( .A1(n_1116), .A2(n_1085), .B1(n_1091), .B2(n_1059), .C(n_1069), .Y(n_1133) );
OAI21xp5_ASAP7_75t_L g1134 ( .A1(n_1120), .A2(n_1091), .B(n_1006), .Y(n_1134) );
NAND3xp33_ASAP7_75t_SL g1135 ( .A(n_1106), .B(n_931), .C(n_935), .Y(n_1135) );
NOR2xp67_ASAP7_75t_SL g1136 ( .A(n_1121), .B(n_915), .Y(n_1136) );
NAND3xp33_ASAP7_75t_SL g1137 ( .A(n_1112), .B(n_931), .C(n_935), .Y(n_1137) );
AOI21xp5_ASAP7_75t_L g1138 ( .A1(n_1107), .A2(n_1005), .B(n_1006), .Y(n_1138) );
AND4x1_ASAP7_75t_L g1139 ( .A(n_1132), .B(n_1122), .C(n_1124), .D(n_1125), .Y(n_1139) );
NAND3x1_ASAP7_75t_L g1140 ( .A(n_1128), .B(n_1130), .C(n_1123), .Y(n_1140) );
NAND3xp33_ASAP7_75t_L g1141 ( .A(n_1128), .B(n_1131), .C(n_1126), .Y(n_1141) );
NAND4xp25_ASAP7_75t_L g1142 ( .A(n_1127), .B(n_1133), .C(n_1138), .D(n_1137), .Y(n_1142) );
NOR3xp33_ASAP7_75t_L g1143 ( .A(n_1135), .B(n_1134), .C(n_1129), .Y(n_1143) );
NOR2x1_ASAP7_75t_L g1144 ( .A(n_1142), .B(n_900), .Y(n_1144) );
NAND2x1p5_ASAP7_75t_L g1145 ( .A(n_1139), .B(n_1136), .Y(n_1145) );
NOR3xp33_ASAP7_75t_L g1146 ( .A(n_1141), .B(n_907), .C(n_906), .Y(n_1146) );
NAND4xp25_ASAP7_75t_L g1147 ( .A(n_1144), .B(n_1143), .C(n_1140), .D(n_958), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1146), .B(n_1062), .Y(n_1148) );
NAND3x2_ASAP7_75t_L g1149 ( .A(n_1145), .B(n_936), .C(n_993), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1148), .Y(n_1150) );
OAI22xp5_ASAP7_75t_SL g1151 ( .A1(n_1147), .A2(n_929), .B1(n_958), .B2(n_936), .Y(n_1151) );
AO22x2_ASAP7_75t_L g1152 ( .A1(n_1150), .A2(n_1149), .B1(n_950), .B2(n_961), .Y(n_1152) );
AO22x2_ASAP7_75t_L g1153 ( .A1(n_1151), .A2(n_965), .B1(n_908), .B2(n_906), .Y(n_1153) );
NAND3xp33_ASAP7_75t_L g1154 ( .A(n_1152), .B(n_915), .C(n_900), .Y(n_1154) );
AOI21xp5_ASAP7_75t_L g1155 ( .A1(n_1152), .A2(n_919), .B(n_949), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1154), .Y(n_1156) );
OAI222xp33_ASAP7_75t_L g1157 ( .A1(n_1155), .A2(n_1153), .B1(n_930), .B2(n_919), .C1(n_1005), .C2(n_907), .Y(n_1157) );
OAI22xp33_ASAP7_75t_L g1158 ( .A1(n_1156), .A2(n_929), .B1(n_900), .B2(n_1005), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_1158), .B(n_1157), .Y(n_1159) );
AOI22xp5_ASAP7_75t_L g1160 ( .A1(n_1159), .A2(n_996), .B1(n_911), .B2(n_908), .Y(n_1160) );
endmodule