module fake_jpeg_28323_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_19),
.B1(n_27),
.B2(n_26),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_56),
.B1(n_57),
.B2(n_64),
.Y(n_68)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_19),
.B1(n_25),
.B2(n_34),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_19),
.B1(n_34),
.B2(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_44),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_27),
.B1(n_26),
.B2(n_16),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_26),
.B1(n_27),
.B2(n_16),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_18),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_16),
.B1(n_21),
.B2(n_30),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_69),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_32),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_75),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_81),
.Y(n_115)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_52),
.A2(n_20),
.B1(n_24),
.B2(n_30),
.Y(n_78)
);

OAI22x1_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_28),
.B1(n_22),
.B2(n_90),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_29),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_33),
.C(n_41),
.Y(n_120)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_20),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_83),
.Y(n_117)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_86),
.A2(n_37),
.B1(n_35),
.B2(n_59),
.Y(n_124)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_88),
.Y(n_121)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_46),
.A2(n_28),
.B1(n_24),
.B2(n_33),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_90),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_48),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_42),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_54),
.Y(n_108)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_94),
.B1(n_50),
.B2(n_40),
.Y(n_119)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_98),
.B(n_112),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_69),
.B1(n_68),
.B2(n_56),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_114),
.B1(n_118),
.B2(n_95),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_103),
.B(n_105),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_68),
.A2(n_54),
.B1(n_43),
.B2(n_57),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_107),
.B1(n_124),
.B2(n_74),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_54),
.B1(n_43),
.B2(n_42),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_70),
.B(n_53),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_32),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_70),
.B(n_58),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_39),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_43),
.B1(n_50),
.B2(n_37),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_50),
.B1(n_37),
.B2(n_62),
.Y(n_118)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_23),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_36),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_114),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_129),
.B1(n_142),
.B2(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_72),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_131),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_127),
.A2(n_131),
.B1(n_146),
.B2(n_154),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_99),
.A2(n_81),
.B1(n_80),
.B2(n_77),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_130),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_67),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_133),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_87),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_84),
.Y(n_134)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_122),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_135),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_148),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_39),
.C(n_36),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_143),
.C(n_152),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_89),
.Y(n_138)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_139),
.A2(n_140),
.B1(n_144),
.B2(n_154),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_88),
.B1(n_91),
.B2(n_94),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_137),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_35),
.B1(n_74),
.B2(n_93),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_36),
.C(n_41),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_83),
.B1(n_35),
.B2(n_49),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_36),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_145),
.B(n_118),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_151),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_85),
.B1(n_48),
.B2(n_41),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_123),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_41),
.C(n_39),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_124),
.C(n_105),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_110),
.C(n_103),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_104),
.A2(n_48),
.B1(n_39),
.B2(n_18),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_104),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_155),
.A2(n_164),
.B(n_174),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_167),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_146),
.A2(n_110),
.B1(n_97),
.B2(n_102),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_121),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_168),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_121),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_127),
.A2(n_112),
.B(n_102),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_171),
.B(n_184),
.Y(n_198)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_176),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_109),
.B(n_100),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_119),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_177),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_119),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_122),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_183),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_18),
.B1(n_31),
.B2(n_23),
.Y(n_206)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_119),
.B1(n_97),
.B2(n_100),
.Y(n_181)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_126),
.B(n_119),
.Y(n_182)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

NAND2x1_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_22),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_187),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_152),
.C(n_139),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_186),
.B(n_142),
.Y(n_192)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_125),
.A2(n_109),
.B1(n_97),
.B2(n_48),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_149),
.B1(n_18),
.B2(n_23),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_156),
.C(n_1),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_159),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_204),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_150),
.B1(n_130),
.B2(n_147),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_202),
.B1(n_203),
.B2(n_206),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_197),
.A2(n_209),
.B1(n_214),
.B2(n_216),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_175),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_201),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_171),
.A2(n_149),
.B1(n_18),
.B2(n_31),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_172),
.A2(n_186),
.B1(n_157),
.B2(n_182),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_31),
.Y(n_204)
);

AOI22x1_ASAP7_75t_SL g205 ( 
.A1(n_184),
.A2(n_174),
.B1(n_181),
.B2(n_155),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_205),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_180),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_207),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_174),
.A2(n_166),
.B1(n_188),
.B2(n_155),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_180),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_210),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_22),
.Y(n_211)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_213),
.B(n_217),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_166),
.A2(n_23),
.B1(n_15),
.B2(n_14),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_161),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_215),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_23),
.B1(n_15),
.B2(n_14),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_2),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_168),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_222),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_177),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_169),
.B(n_183),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_194),
.B(n_198),
.Y(n_251)
);

OAI21x1_ASAP7_75t_SL g226 ( 
.A1(n_205),
.A2(n_167),
.B(n_158),
.Y(n_226)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_218),
.A2(n_156),
.B1(n_160),
.B2(n_2),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_206),
.B1(n_202),
.B2(n_213),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_239),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_198),
.C(n_201),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_234),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_238),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_216),
.B1(n_214),
.B2(n_217),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_191),
.B(n_11),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_237),
.B(n_189),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_13),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_13),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_196),
.Y(n_248)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_189),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_195),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_244),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_248),
.B(n_253),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_219),
.A2(n_215),
.B1(n_209),
.B2(n_200),
.Y(n_250)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_250),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_256),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_259),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_211),
.Y(n_255)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_208),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_263),
.B1(n_190),
.B2(n_236),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_195),
.C(n_199),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_261),
.C(n_237),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_240),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_199),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_233),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_221),
.A2(n_190),
.B1(n_207),
.B2(n_210),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_267),
.C(n_4),
.Y(n_293)
);

XNOR2x1_ASAP7_75t_SL g267 ( 
.A(n_251),
.B(n_225),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_222),
.C(n_227),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_271),
.C(n_274),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_241),
.C(n_219),
.Y(n_271)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_273),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_242),
.C(n_238),
.Y(n_274)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_230),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_279),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_223),
.C(n_221),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_261),
.C(n_256),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_247),
.A2(n_235),
.B1(n_197),
.B2(n_11),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_260),
.B(n_254),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_265),
.B(n_281),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_269),
.A2(n_263),
.B1(n_264),
.B2(n_249),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_270),
.A2(n_248),
.B(n_246),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_289),
.A2(n_292),
.B(n_278),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_290),
.B(n_294),
.Y(n_297)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_272),
.B(n_246),
.CI(n_3),
.CON(n_291),
.SN(n_291)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_291),
.A2(n_8),
.B(n_9),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_2),
.B(n_4),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_280),
.C(n_266),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_4),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_277),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_295),
.A2(n_296),
.B1(n_292),
.B2(n_286),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_280),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_298),
.A2(n_308),
.B(n_289),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_301),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_285),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_271),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_303),
.B(n_288),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_282),
.B(n_274),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_306),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_5),
.C(n_6),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_294),
.C(n_293),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_7),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_8),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_308),
.Y(n_313)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_313),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_303),
.A2(n_296),
.B1(n_284),
.B2(n_290),
.Y(n_314)
);

OAI211xp5_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_316),
.B(n_317),
.C(n_291),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_295),
.Y(n_315)
);

AOI21xp33_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_300),
.B(n_298),
.Y(n_320)
);

OAI211xp5_ASAP7_75t_L g325 ( 
.A1(n_320),
.A2(n_323),
.B(n_319),
.C(n_321),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_297),
.C(n_305),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_310),
.C(n_315),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_316),
.A2(n_299),
.B(n_291),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_9),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_324),
.A2(n_325),
.B(n_326),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_318),
.B(n_9),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_10),
.C(n_313),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_10),
.Y(n_331)
);


endmodule