module real_jpeg_18000_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_622, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_622;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_195;
wire n_110;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_594;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_608;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_1),
.A2(n_83),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_1),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_1),
.A2(n_152),
.B1(n_266),
.B2(n_269),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_1),
.A2(n_152),
.B1(n_460),
.B2(n_463),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_SL g470 ( 
.A1(n_1),
.A2(n_152),
.B1(n_471),
.B2(n_473),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_2),
.A2(n_119),
.B1(n_123),
.B2(n_125),
.Y(n_118)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_2),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_2),
.A2(n_125),
.B1(n_195),
.B2(n_200),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_2),
.A2(n_125),
.B1(n_325),
.B2(n_334),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g558 ( 
.A1(n_2),
.A2(n_125),
.B1(n_318),
.B2(n_559),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_3),
.A2(n_128),
.B1(n_129),
.B2(n_131),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_3),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_3),
.A2(n_128),
.B1(n_292),
.B2(n_296),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_3),
.A2(n_128),
.B1(n_437),
.B2(n_442),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_3),
.A2(n_124),
.B1(n_128),
.B2(n_493),
.Y(n_492)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_4),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_4),
.Y(n_354)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_5),
.Y(n_89)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_5),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_5),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_5),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_6),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_6),
.A2(n_39),
.B1(n_247),
.B2(n_249),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_6),
.A2(n_39),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_6),
.A2(n_39),
.B1(n_447),
.B2(n_449),
.Y(n_446)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_7),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_7),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_7),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_7),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_8),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_8),
.A2(n_71),
.B1(n_275),
.B2(n_278),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_8),
.A2(n_71),
.B1(n_317),
.B2(n_320),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_8),
.A2(n_71),
.B1(n_407),
.B2(n_412),
.Y(n_406)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_9),
.B(n_155),
.Y(n_306)
);

OAI32xp33_ASAP7_75t_L g398 ( 
.A1(n_9),
.A2(n_47),
.A3(n_275),
.B1(n_399),
.B2(n_402),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_9),
.B(n_77),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_9),
.A2(n_101),
.B1(n_238),
.B2(n_492),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_SL g510 ( 
.A1(n_9),
.A2(n_81),
.B1(n_511),
.B2(n_512),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_10),
.A2(n_174),
.B1(n_176),
.B2(n_178),
.Y(n_173)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_10),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_10),
.A2(n_178),
.B1(n_346),
.B2(n_348),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_10),
.A2(n_178),
.B1(n_334),
.B2(n_566),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_SL g607 ( 
.A1(n_10),
.A2(n_178),
.B1(n_596),
.B2(n_608),
.Y(n_607)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_11),
.Y(n_106)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_11),
.Y(n_115)
);

BUFx4f_ASAP7_75t_L g122 ( 
.A(n_11),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_11),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_12),
.A2(n_162),
.B1(n_165),
.B2(n_166),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_12),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_12),
.A2(n_165),
.B1(n_340),
.B2(n_343),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_12),
.A2(n_165),
.B1(n_550),
.B2(n_552),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_SL g595 ( 
.A1(n_12),
.A2(n_82),
.B1(n_165),
.B2(n_596),
.Y(n_595)
);

OAI22xp33_ASAP7_75t_L g108 ( 
.A1(n_13),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_13),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_13),
.A2(n_110),
.B1(n_220),
.B2(n_222),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_13),
.A2(n_110),
.B1(n_323),
.B2(n_326),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g542 ( 
.A1(n_13),
.A2(n_110),
.B1(n_543),
.B2(n_546),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_21),
.B(n_23),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_16),
.A2(n_231),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_16),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_16),
.A2(n_233),
.B1(n_253),
.B2(n_255),
.Y(n_252)
);

OAI22x1_ASAP7_75t_SL g298 ( 
.A1(n_16),
.A2(n_233),
.B1(n_299),
.B2(n_301),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_16),
.A2(n_233),
.B1(n_318),
.B2(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_17),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_17),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_17),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_17),
.Y(n_236)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_17),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

BUFx8_ASAP7_75t_L g130 ( 
.A(n_19),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_19),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g319 ( 
.A(n_19),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_616),
.B(n_619),
.Y(n_24)
);

AO21x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_533),
.B(n_609),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_379),
.B(n_528),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_310),
.C(n_374),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_258),
.B(n_283),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_29),
.B(n_258),
.C(n_530),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_156),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_30),
.B(n_157),
.C(n_226),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_78),
.C(n_126),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_32),
.B(n_126),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_46),
.B1(n_68),
.B2(n_76),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_34),
.A2(n_77),
.B1(n_265),
.B2(n_270),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_43),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_45),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_45),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_45),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_45),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_46),
.A2(n_68),
.B1(n_76),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_46),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_46),
.A2(n_76),
.B1(n_252),
.B2(n_322),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_46),
.A2(n_76),
.B1(n_291),
.B2(n_510),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_46),
.A2(n_76),
.B1(n_333),
.B2(n_549),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_46),
.A2(n_76),
.B1(n_549),
.B2(n_565),
.Y(n_564)
);

AO21x2_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_53),
.B(n_61),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_58),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_60),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_62),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_62),
.Y(n_232)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_62),
.Y(n_342)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_66),
.Y(n_344)
);

INVx6_ASAP7_75t_L g420 ( 
.A(n_66),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_67),
.Y(n_277)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_77),
.A2(n_265),
.B1(n_270),
.B2(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_77),
.A2(n_270),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g591 ( 
.A1(n_77),
.A2(n_270),
.B(n_592),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_78),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_100),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_79),
.B(n_100),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_86),
.B1(n_94),
.B2(n_95),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_SL g272 ( 
.A1(n_80),
.A2(n_81),
.B(n_129),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_81),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_81),
.B(n_424),
.Y(n_423)
);

OAI21xp33_ASAP7_75t_SL g434 ( 
.A1(n_81),
.A2(n_423),
.B(n_435),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_81),
.B(n_305),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_81),
.B(n_182),
.Y(n_498)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g248 ( 
.A(n_85),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_85),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_93),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_96),
.A2(n_135),
.B(n_139),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_99),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_107),
.B1(n_116),
.B2(n_118),
.Y(n_100)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_101),
.A2(n_118),
.B1(n_161),
.B2(n_238),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_101),
.A2(n_173),
.B(n_353),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_101),
.A2(n_171),
.B1(n_446),
.B2(n_454),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_101),
.A2(n_470),
.B1(n_492),
.B2(n_496),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_105),
.Y(n_421)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_106),
.Y(n_300)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_106),
.Y(n_411)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22x1_ASAP7_75t_SL g297 ( 
.A1(n_108),
.A2(n_159),
.B1(n_298),
.B2(n_304),
.Y(n_297)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_113),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_114),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_115),
.Y(n_169)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_121),
.Y(n_412)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_122),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_122),
.Y(n_448)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_134),
.B1(n_150),
.B2(n_155),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_127),
.A2(n_134),
.B1(n_155),
.B2(n_272),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_134),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_134),
.A2(n_155),
.B1(n_557),
.B2(n_558),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_134),
.A2(n_155),
.B(n_618),
.Y(n_617)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_L g315 ( 
.A1(n_139),
.A2(n_244),
.B1(n_246),
.B2(n_316),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_139),
.A2(n_244),
.B1(n_316),
.B2(n_361),
.Y(n_360)
);

AOI22x1_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_143),
.B1(n_145),
.B2(n_148),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_146),
.Y(n_327)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_147),
.Y(n_569)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22x1_ASAP7_75t_SL g243 ( 
.A1(n_151),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_243)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_155),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_226),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_179),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_158),
.A2(n_180),
.B(n_205),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_170),
.B2(n_172),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_159),
.A2(n_239),
.B1(n_298),
.B2(n_406),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_159),
.A2(n_469),
.B1(n_476),
.B2(n_477),
.Y(n_468)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_205),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_193),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_181),
.A2(n_206),
.B1(n_274),
.B2(n_282),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_181),
.A2(n_206),
.B1(n_338),
.B2(n_345),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_181),
.A2(n_206),
.B1(n_434),
.B2(n_436),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_181),
.A2(n_206),
.B1(n_436),
.B2(n_459),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_181),
.A2(n_206),
.B1(n_389),
.B2(n_459),
.Y(n_518)
);

OA21x2_ASAP7_75t_L g539 ( 
.A1(n_181),
.A2(n_206),
.B(n_345),
.Y(n_539)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_182),
.A2(n_219),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_182),
.A2(n_194),
.B1(n_229),
.B2(n_339),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_182),
.A2(n_229),
.B1(n_388),
.B2(n_395),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_183),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_187),
.B1(n_188),
.B2(n_191),
.Y(n_183)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_190),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_190),
.Y(n_472)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_190),
.Y(n_489)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_192),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_199),
.Y(n_204)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_199),
.Y(n_281)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_218),
.Y(n_205)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_212),
.B1(n_215),
.B2(n_217),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_211),
.Y(n_347)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_211),
.Y(n_394)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_215),
.Y(n_422)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_221),
.Y(n_348)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_242),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_227),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_237),
.Y(n_227)
);

XOR2x2_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_237),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_230),
.Y(n_282)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_235),
.Y(n_464)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_238),
.Y(n_476)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_240),
.Y(n_305)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_251),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_243),
.B(n_251),
.C(n_373),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_244),
.A2(n_245),
.B1(n_361),
.B2(n_542),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_244),
.A2(n_245),
.B1(n_594),
.B2(n_595),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_244),
.A2(n_245),
.B1(n_595),
.B2(n_607),
.Y(n_606)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_256),
.Y(n_269)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_256),
.Y(n_553)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_257),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.C(n_263),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_259),
.A2(n_260),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_262),
.B(n_263),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_271),
.C(n_273),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_273),
.Y(n_286)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_286),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_274),
.Y(n_395)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_280),
.Y(n_403)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_307),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_284),
.B(n_307),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.C(n_288),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_285),
.B(n_382),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_287),
.B(n_288),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_297),
.C(n_306),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_289),
.B(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx2_ASAP7_75t_SL g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_295),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_295),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_297),
.B(n_306),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_299),
.Y(n_493)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

A2O1A1O1Ixp25_ASAP7_75t_L g528 ( 
.A1(n_310),
.A2(n_374),
.B(n_529),
.C(n_531),
.D(n_532),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_365),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_311),
.B(n_365),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_328),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_312),
.B(n_583),
.C(n_584),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.C(n_321),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_313),
.B(n_368),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_315),
.B(n_321),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_317),
.Y(n_320)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx8_ASAP7_75t_L g547 ( 
.A(n_319),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_322),
.Y(n_331)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_325),
.Y(n_511)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_325),
.Y(n_551)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_350),
.Y(n_328)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_329),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_330),
.A2(n_337),
.B(n_349),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_330),
.B(n_337),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_340),
.Y(n_435)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_342),
.Y(n_390)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_349),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_349),
.A2(n_575),
.B1(n_577),
.B2(n_587),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_350),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_351),
.A2(n_356),
.B1(n_357),
.B2(n_364),
.Y(n_350)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_351),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_355),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_352),
.A2(n_358),
.B1(n_359),
.B2(n_360),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_352),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_352),
.A2(n_355),
.B1(n_358),
.B2(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx12f_ASAP7_75t_L g497 ( 
.A(n_354),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_355),
.Y(n_370)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_358),
.A2(n_364),
.B1(n_579),
.B2(n_622),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_359),
.Y(n_580)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx5_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_369),
.C(n_371),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_366),
.A2(n_367),
.B1(n_369),
.B2(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_369),
.Y(n_377)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_372),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_378),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_375),
.B(n_378),
.Y(n_531)
);

AOI21x1_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_413),
.B(n_527),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_383),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_381),
.B(n_383),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_387),
.C(n_396),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_384),
.A2(n_385),
.B1(n_522),
.B2(n_523),
.Y(n_521)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_387),
.A2(n_396),
.B1(n_397),
.B2(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_387),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_404),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_398),
.A2(n_404),
.B1(n_405),
.B2(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_398),
.Y(n_506)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_403),
.Y(n_424)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_406),
.Y(n_454)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

OAI21x1_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_520),
.B(n_526),
.Y(n_413)
);

AOI21x1_ASAP7_75t_SL g414 ( 
.A1(n_415),
.A2(n_502),
.B(n_519),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g415 ( 
.A1(n_416),
.A2(n_466),
.B(n_501),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_444),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_417),
.B(n_444),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_432),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_418),
.A2(n_432),
.B1(n_433),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_418),
.Y(n_479)
);

OAI32xp33_ASAP7_75t_L g418 ( 
.A1(n_419),
.A2(n_421),
.A3(n_422),
.B1(n_423),
.B2(n_425),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_429),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_441),
.Y(n_443)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_441),
.Y(n_462)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_455),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_445),
.B(n_457),
.C(n_465),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_446),
.Y(n_477)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_456),
.A2(n_457),
.B1(n_458),
.B2(n_465),
.Y(n_455)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_456),
.Y(n_465)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_467),
.A2(n_480),
.B(n_500),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_478),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_468),
.B(n_478),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_475),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_481),
.A2(n_494),
.B(n_499),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_491),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_490),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_498),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_495),
.B(n_498),
.Y(n_499)
);

INVx6_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_504),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_504),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_507),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_505),
.B(n_508),
.C(n_518),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_508),
.A2(n_509),
.B1(n_517),
.B2(n_518),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_SL g520 ( 
.A(n_521),
.B(n_525),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_521),
.B(n_525),
.Y(n_526)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

NOR3xp33_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_588),
.C(n_604),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_581),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g611 ( 
.A1(n_536),
.A2(n_612),
.B(n_613),
.Y(n_611)
);

NOR2x1_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_574),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_537),
.B(n_574),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_554),
.Y(n_537)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_538),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_540),
.C(n_548),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_539),
.A2(n_564),
.B1(n_570),
.B2(n_571),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_539),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_539),
.B(n_548),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_539),
.B(n_556),
.C(n_571),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_540),
.A2(n_555),
.B1(n_572),
.B2(n_573),
.Y(n_554)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_540),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_540),
.B(n_576),
.Y(n_575)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_542),
.Y(n_557)
);

INVx6_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx5_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx8_ASAP7_75t_L g562 ( 
.A(n_545),
.Y(n_562)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_545),
.Y(n_600)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_547),
.Y(n_546)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_555),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_555),
.B(n_572),
.C(n_603),
.Y(n_602)
);

XNOR2x1_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_563),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_558),
.Y(n_594)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx6_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_564),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_565),
.Y(n_592)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_575),
.B(n_577),
.C(n_578),
.Y(n_574)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_575),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_578),
.B(n_586),
.Y(n_585)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_582),
.B(n_585),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_582),
.B(n_585),
.Y(n_612)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

A2O1A1O1Ixp25_ASAP7_75t_L g610 ( 
.A1(n_589),
.A2(n_605),
.B(n_611),
.C(n_614),
.D(n_615),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_590),
.B(n_602),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_590),
.B(n_606),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_590),
.B(n_602),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_590),
.B(n_606),
.Y(n_615)
);

FAx1_ASAP7_75t_SL g590 ( 
.A(n_591),
.B(n_593),
.CI(n_601),
.CON(n_590),
.SN(n_590)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_597),
.Y(n_608)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_606),
.B(n_617),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_606),
.B(n_617),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_607),
.Y(n_618)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

CKINVDCx16_ASAP7_75t_R g619 ( 
.A(n_620),
.Y(n_619)
);


endmodule