module fake_netlist_6_4259_n_503 (n_52, n_16, n_1, n_46, n_18, n_21, n_3, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_5, n_77, n_42, n_8, n_24, n_54, n_0, n_32, n_66, n_78, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_27, n_38, n_61, n_59, n_76, n_36, n_26, n_55, n_58, n_64, n_48, n_65, n_25, n_40, n_41, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_60, n_35, n_12, n_69, n_30, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_503);

input n_52;
input n_16;
input n_1;
input n_46;
input n_18;
input n_21;
input n_3;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_5;
input n_77;
input n_42;
input n_8;
input n_24;
input n_54;
input n_0;
input n_32;
input n_66;
input n_78;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_27;
input n_38;
input n_61;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_41;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_503;

wire n_435;
wire n_91;
wire n_326;
wire n_256;
wire n_440;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_106;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_495;
wire n_350;
wire n_84;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_114;
wire n_198;
wire n_86;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_468;
wire n_111;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_79;
wire n_375;
wire n_338;
wire n_466;
wire n_360;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_96;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_493;
wire n_397;
wire n_155;
wire n_109;
wire n_445;
wire n_425;
wire n_122;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_82;
wire n_236;
wire n_112;
wire n_172;
wire n_472;
wire n_270;
wire n_239;
wire n_126;
wire n_414;
wire n_97;
wire n_490;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_93;
wire n_80;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_460;
wire n_107;
wire n_417;
wire n_446;
wire n_498;
wire n_89;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_103;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_154;
wire n_456;
wire n_98;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_455;
wire n_83;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_152;
wire n_92;
wire n_321;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_406;
wire n_483;
wire n_102;
wire n_204;
wire n_482;
wire n_474;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_130;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_477;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_124;
wire n_94;
wire n_282;
wire n_436;
wire n_116;
wire n_211;
wire n_175;
wire n_117;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_95;
wire n_311;
wire n_403;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_487;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_88;
wire n_416;
wire n_277;
wire n_418;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_90;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_488;
wire n_429;
wire n_373;
wire n_87;
wire n_195;
wire n_285;
wire n_497;
wire n_85;
wire n_99;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_489;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_110;
wire n_412;
wire n_81;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVx1_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVxp67_ASAP7_75t_SL g80 ( 
.A(n_47),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_61),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_7),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_12),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_52),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_8),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_15),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVxp67_ASAP7_75t_SL g93 ( 
.A(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_7),
.Y(n_94)
);

INVxp33_ASAP7_75t_SL g95 ( 
.A(n_31),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_14),
.Y(n_96)
);

BUFx2_ASAP7_75t_SL g97 ( 
.A(n_13),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_45),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVxp33_ASAP7_75t_SL g101 ( 
.A(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_12),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_29),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_49),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_58),
.Y(n_107)
);

INVxp33_ASAP7_75t_SL g108 ( 
.A(n_38),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_35),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_8),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

NOR2xp67_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_56),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_32),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_1),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_11),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_1),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_11),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_48),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_41),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_30),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_20),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_44),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_17),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_14),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_72),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_16),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_5),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_22),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g140 ( 
.A(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_9),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_9),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_15),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_18),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_6),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_21),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_19),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_10),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_33),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_26),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_97),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_90),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_90),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_122),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_122),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_135),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_81),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_81),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_89),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_89),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_107),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_107),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_99),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_91),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

NOR2xp67_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_0),
.Y(n_174)
);

INVx3_ASAP7_75t_SL g175 ( 
.A(n_104),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_2),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_124),
.B(n_2),
.Y(n_177)
);

AND3x2_ASAP7_75t_L g178 ( 
.A(n_103),
.B(n_3),
.C(n_4),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_104),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_105),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_R g184 ( 
.A(n_146),
.B(n_28),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_125),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_129),
.B(n_3),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_95),
.B(n_4),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_R g190 ( 
.A(n_150),
.B(n_36),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_150),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_82),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_82),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_101),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_101),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_108),
.B(n_5),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_R g197 ( 
.A(n_96),
.B(n_37),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_147),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_108),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_96),
.Y(n_202)
);

AO21x2_ASAP7_75t_L g203 ( 
.A1(n_109),
.A2(n_148),
.B(n_113),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_136),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_79),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_136),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_142),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_142),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_143),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_121),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_83),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_143),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_R g213 ( 
.A(n_129),
.B(n_39),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_121),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_84),
.Y(n_215)
);

NAND2x1_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_121),
.Y(n_216)
);

AO22x2_ASAP7_75t_L g217 ( 
.A1(n_177),
.A2(n_120),
.B1(n_144),
.B2(n_133),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_111),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_171),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

AND2x6_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_148),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_153),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_157),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_185),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_176),
.A2(n_137),
.B1(n_113),
.B2(n_132),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_189),
.A2(n_196),
.B1(n_163),
.B2(n_200),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

AO22x2_ASAP7_75t_L g235 ( 
.A1(n_188),
.A2(n_154),
.B1(n_109),
.B2(n_199),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_180),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_174),
.B(n_114),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_201),
.Y(n_239)
);

OAI221xp5_ASAP7_75t_L g240 ( 
.A1(n_201),
.A2(n_126),
.B1(n_139),
.B2(n_138),
.C(n_131),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_175),
.B(n_85),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_173),
.Y(n_242)
);

NAND3xp33_ASAP7_75t_L g243 ( 
.A(n_199),
.B(n_172),
.C(n_169),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_203),
.A2(n_86),
.B1(n_130),
.B2(n_128),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

OR2x2_ASAP7_75t_SL g246 ( 
.A(n_152),
.B(n_123),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_186),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_186),
.Y(n_248)
);

NAND2x1p5_ASAP7_75t_L g249 ( 
.A(n_154),
.B(n_110),
.Y(n_249)
);

NOR2x1p5_ASAP7_75t_L g250 ( 
.A(n_191),
.B(n_140),
.Y(n_250)
);

AND2x6_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_117),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_185),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_179),
.B(n_116),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_93),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_194),
.A2(n_80),
.B1(n_100),
.B2(n_98),
.Y(n_255)
);

AND2x6_ASAP7_75t_L g256 ( 
.A(n_184),
.B(n_115),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_185),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_181),
.Y(n_258)
);

AND2x6_ASAP7_75t_SL g259 ( 
.A(n_192),
.B(n_92),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_194),
.A2(n_10),
.B1(n_13),
.B2(n_16),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_200),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_261)
);

NAND2xp33_ASAP7_75t_L g262 ( 
.A(n_191),
.B(n_25),
.Y(n_262)
);

AO22x2_ASAP7_75t_L g263 ( 
.A1(n_193),
.A2(n_40),
.B1(n_46),
.B2(n_67),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_156),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_233),
.A2(n_195),
.B1(n_187),
.B2(n_155),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_239),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_226),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_223),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_155),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_159),
.B1(n_162),
.B2(n_158),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_227),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_159),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_216),
.A2(n_162),
.B(n_158),
.Y(n_274)
);

BUFx4f_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_228),
.Y(n_276)
);

NAND3xp33_ASAP7_75t_SL g277 ( 
.A(n_255),
.B(n_197),
.C(n_170),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_221),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_238),
.B(n_190),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_230),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_SL g282 ( 
.A1(n_245),
.A2(n_178),
.B(n_161),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_231),
.A2(n_156),
.B1(n_168),
.B2(n_166),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_254),
.A2(n_167),
.B(n_165),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_242),
.B(n_161),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_224),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_254),
.A2(n_164),
.B(n_212),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_161),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_258),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_235),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_247),
.B(n_209),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_225),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_250),
.A2(n_204),
.B1(n_207),
.B2(n_206),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_246),
.A2(n_208),
.B1(n_202),
.B2(n_77),
.Y(n_295)
);

AOI221xp5_ASAP7_75t_L g296 ( 
.A1(n_217),
.A2(n_71),
.B1(n_75),
.B2(n_261),
.C(n_260),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_248),
.Y(n_297)
);

NAND2x1p5_ASAP7_75t_L g298 ( 
.A(n_253),
.B(n_218),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_220),
.Y(n_299)
);

O2A1O1Ixp33_ASAP7_75t_L g300 ( 
.A1(n_240),
.A2(n_222),
.B(n_262),
.C(n_234),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_219),
.B(n_249),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_236),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_241),
.A2(n_235),
.B(n_237),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_229),
.Y(n_304)
);

CKINVDCx6p67_ASAP7_75t_R g305 ( 
.A(n_256),
.Y(n_305)
);

O2A1O1Ixp33_ASAP7_75t_SL g306 ( 
.A1(n_243),
.A2(n_263),
.B(n_252),
.C(n_257),
.Y(n_306)
);

BUFx8_ASAP7_75t_L g307 ( 
.A(n_251),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_223),
.Y(n_308)
);

INVx3_ASAP7_75t_SL g309 ( 
.A(n_217),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_243),
.A2(n_263),
.B(n_251),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_251),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

INVx3_ASAP7_75t_SL g313 ( 
.A(n_278),
.Y(n_313)
);

O2A1O1Ixp33_ASAP7_75t_L g314 ( 
.A1(n_266),
.A2(n_291),
.B(n_300),
.C(n_301),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_269),
.B(n_301),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_267),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_282),
.Y(n_317)
);

AOI21xp33_ASAP7_75t_SL g318 ( 
.A1(n_283),
.A2(n_273),
.B(n_285),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_269),
.B(n_304),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_309),
.Y(n_320)
);

AND2x4_ASAP7_75t_L g321 ( 
.A(n_272),
.B(n_287),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_276),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_299),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_275),
.A2(n_311),
.B1(n_305),
.B2(n_270),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_297),
.Y(n_325)
);

OA21x2_ASAP7_75t_L g326 ( 
.A1(n_293),
.A2(n_286),
.B(n_302),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_271),
.B(n_309),
.Y(n_327)
);

OAI21x1_ASAP7_75t_L g328 ( 
.A1(n_274),
.A2(n_298),
.B(n_310),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_268),
.A2(n_265),
.B1(n_289),
.B2(n_298),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_290),
.Y(n_330)
);

OAI21x1_ASAP7_75t_L g331 ( 
.A1(n_295),
.A2(n_279),
.B(n_284),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_297),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_279),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_288),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_296),
.A2(n_277),
.B(n_292),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_307),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_307),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_306),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_294),
.A2(n_266),
.B1(n_244),
.B2(n_275),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_306),
.Y(n_341)
);

OAI21x1_ASAP7_75t_SL g342 ( 
.A1(n_310),
.A2(n_244),
.B(n_303),
.Y(n_342)
);

OAI21x1_ASAP7_75t_L g343 ( 
.A1(n_308),
.A2(n_245),
.B(n_239),
.Y(n_343)
);

OA21x2_ASAP7_75t_L g344 ( 
.A1(n_303),
.A2(n_245),
.B(n_239),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_266),
.B(n_245),
.Y(n_346)
);

OA21x2_ASAP7_75t_L g347 ( 
.A1(n_303),
.A2(n_245),
.B(n_239),
.Y(n_347)
);

O2A1O1Ixp33_ASAP7_75t_L g348 ( 
.A1(n_266),
.A2(n_239),
.B(n_245),
.C(n_291),
.Y(n_348)
);

NAND2x1p5_ASAP7_75t_L g349 ( 
.A(n_275),
.B(n_268),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_266),
.B(n_245),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_266),
.B(n_245),
.Y(n_351)
);

AO21x1_ASAP7_75t_L g352 ( 
.A1(n_266),
.A2(n_188),
.B(n_310),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_267),
.Y(n_353)
);

OR3x4_ASAP7_75t_SL g354 ( 
.A(n_296),
.B(n_120),
.C(n_93),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_267),
.Y(n_355)
);

OA21x2_ASAP7_75t_L g356 ( 
.A1(n_303),
.A2(n_245),
.B(n_239),
.Y(n_356)
);

OAI21x1_ASAP7_75t_L g357 ( 
.A1(n_308),
.A2(n_245),
.B(n_239),
.Y(n_357)
);

AO21x2_ASAP7_75t_L g358 ( 
.A1(n_266),
.A2(n_303),
.B(n_239),
.Y(n_358)
);

A2O1A1Ixp33_ASAP7_75t_L g359 ( 
.A1(n_266),
.A2(n_245),
.B(n_310),
.C(n_189),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_297),
.Y(n_360)
);

OAI21x1_ASAP7_75t_L g361 ( 
.A1(n_308),
.A2(n_245),
.B(n_239),
.Y(n_361)
);

OAI21x1_ASAP7_75t_L g362 ( 
.A1(n_308),
.A2(n_245),
.B(n_239),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_266),
.A2(n_245),
.B(n_244),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_291),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_316),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_320),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_313),
.Y(n_367)
);

O2A1O1Ixp33_ASAP7_75t_SL g368 ( 
.A1(n_359),
.A2(n_338),
.B(n_363),
.C(n_314),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_322),
.Y(n_369)
);

AND2x4_ASAP7_75t_SL g370 ( 
.A(n_337),
.B(n_332),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_319),
.B(n_360),
.Y(n_371)
);

AO31x2_ASAP7_75t_L g372 ( 
.A1(n_352),
.A2(n_359),
.A3(n_340),
.B(n_350),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_353),
.Y(n_373)
);

OR2x6_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_337),
.Y(n_374)
);

INVx8_ASAP7_75t_L g375 ( 
.A(n_332),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_325),
.B(n_315),
.Y(n_376)
);

AO31x2_ASAP7_75t_L g377 ( 
.A1(n_352),
.A2(n_351),
.A3(n_329),
.B(n_317),
.Y(n_377)
);

AO32x2_ASAP7_75t_L g378 ( 
.A1(n_324),
.A2(n_354),
.A3(n_358),
.B1(n_342),
.B2(n_348),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_315),
.B(n_313),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_335),
.A2(n_333),
.B1(n_334),
.B2(n_317),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_355),
.Y(n_381)
);

NAND2xp33_ASAP7_75t_R g382 ( 
.A(n_327),
.B(n_345),
.Y(n_382)
);

OR2x6_ASAP7_75t_L g383 ( 
.A(n_332),
.B(n_328),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_326),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_330),
.B(n_332),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_326),
.Y(n_386)
);

OR2x6_ASAP7_75t_L g387 ( 
.A(n_332),
.B(n_328),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_330),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_312),
.B(n_364),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_318),
.B(n_345),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_R g391 ( 
.A(n_337),
.B(n_320),
.Y(n_391)
);

NOR3xp33_ASAP7_75t_SL g392 ( 
.A(n_323),
.B(n_354),
.C(n_327),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_321),
.B(n_346),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_346),
.A2(n_335),
.B1(n_341),
.B2(n_321),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_341),
.A2(n_331),
.B1(n_321),
.B2(n_336),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_331),
.B(n_341),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_358),
.B(n_347),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_344),
.B(n_356),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_339),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_339),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_341),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_343),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_344),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_339),
.Y(n_406)
);

INVx6_ASAP7_75t_L g407 ( 
.A(n_375),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_384),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_401),
.A2(n_395),
.B1(n_393),
.B2(n_403),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_389),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_390),
.A2(n_371),
.B1(n_376),
.B2(n_380),
.Y(n_411)
);

OAI21xp33_ASAP7_75t_L g412 ( 
.A1(n_392),
.A2(n_357),
.B(n_362),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_386),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_382),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_394),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_379),
.B(n_385),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_401),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_404),
.Y(n_419)
);

AOI221xp5_ASAP7_75t_L g420 ( 
.A1(n_365),
.A2(n_339),
.B1(n_349),
.B2(n_357),
.C(n_361),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_405),
.Y(n_421)
);

AOI221xp5_ASAP7_75t_L g422 ( 
.A1(n_369),
.A2(n_361),
.B1(n_362),
.B2(n_373),
.C(n_381),
.Y(n_422)
);

A2O1A1Ixp33_ASAP7_75t_L g423 ( 
.A1(n_397),
.A2(n_396),
.B(n_370),
.C(n_398),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_368),
.Y(n_424)
);

OR2x2_ASAP7_75t_SL g425 ( 
.A(n_366),
.B(n_391),
.Y(n_425)
);

NOR3xp33_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_367),
.C(n_388),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_399),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_397),
.Y(n_428)
);

NOR3xp33_ASAP7_75t_L g429 ( 
.A(n_367),
.B(n_388),
.C(n_400),
.Y(n_429)
);

INVxp33_ASAP7_75t_L g430 ( 
.A(n_410),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_417),
.B(n_378),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_408),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_408),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_417),
.B(n_372),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_413),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_428),
.B(n_370),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_414),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_413),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_418),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_415),
.B(n_372),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_378),
.Y(n_441)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_407),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_409),
.A2(n_374),
.B1(n_383),
.B2(n_387),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_427),
.B(n_378),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_416),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_416),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_372),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_372),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_425),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_432),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_448),
.A2(n_426),
.B1(n_429),
.B2(n_409),
.Y(n_451)
);

NAND3xp33_ASAP7_75t_L g452 ( 
.A(n_437),
.B(n_420),
.C(n_400),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_432),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_418),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_433),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_436),
.B(n_423),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_433),
.Y(n_457)
);

AO21x2_ASAP7_75t_L g458 ( 
.A1(n_443),
.A2(n_412),
.B(n_419),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_421),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_434),
.B(n_377),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_435),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_430),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_448),
.Y(n_464)
);

AOI33xp33_ASAP7_75t_L g465 ( 
.A1(n_438),
.A2(n_446),
.A3(n_445),
.B1(n_441),
.B2(n_431),
.B3(n_422),
.Y(n_465)
);

NOR2x1_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_374),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_464),
.B(n_431),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_460),
.B(n_441),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_453),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_459),
.B(n_440),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_438),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_447),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_451),
.B(n_446),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_453),
.B(n_444),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_462),
.Y(n_475)
);

AOI221xp5_ASAP7_75t_L g476 ( 
.A1(n_452),
.A2(n_412),
.B1(n_391),
.B2(n_402),
.C(n_424),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_462),
.B(n_444),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_475),
.B(n_456),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_471),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_476),
.B(n_456),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_465),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_475),
.Y(n_482)
);

NAND3xp33_ASAP7_75t_L g483 ( 
.A(n_473),
.B(n_465),
.C(n_443),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_472),
.Y(n_484)
);

OAI31xp33_ASAP7_75t_SL g485 ( 
.A1(n_467),
.A2(n_456),
.A3(n_466),
.B(n_454),
.Y(n_485)
);

AOI221xp5_ASAP7_75t_L g486 ( 
.A1(n_483),
.A2(n_469),
.B1(n_467),
.B2(n_468),
.C(n_450),
.Y(n_486)
);

AOI221xp5_ASAP7_75t_L g487 ( 
.A1(n_481),
.A2(n_479),
.B1(n_484),
.B2(n_480),
.C(n_478),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_R g488 ( 
.A(n_478),
.B(n_402),
.Y(n_488)
);

OAI21xp33_ASAP7_75t_L g489 ( 
.A1(n_485),
.A2(n_468),
.B(n_374),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_480),
.A2(n_439),
.B(n_461),
.Y(n_490)
);

AOI32xp33_ASAP7_75t_L g491 ( 
.A1(n_482),
.A2(n_474),
.A3(n_454),
.B1(n_457),
.B2(n_455),
.Y(n_491)
);

OAI211xp5_ASAP7_75t_L g492 ( 
.A1(n_482),
.A2(n_366),
.B(n_439),
.C(n_477),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_486),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_490),
.A2(n_383),
.B(n_387),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_489),
.A2(n_383),
.B(n_387),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_493),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_494),
.Y(n_497)
);

AOI222xp33_ASAP7_75t_L g498 ( 
.A1(n_495),
.A2(n_487),
.B1(n_492),
.B2(n_474),
.C1(n_454),
.C2(n_424),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_496),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_499),
.Y(n_500)
);

OAI221xp5_ASAP7_75t_L g501 ( 
.A1(n_500),
.A2(n_497),
.B1(n_498),
.B2(n_491),
.C(n_488),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_501),
.A2(n_498),
.B1(n_458),
.B2(n_442),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_502),
.A2(n_458),
.B1(n_445),
.B2(n_442),
.Y(n_503)
);


endmodule