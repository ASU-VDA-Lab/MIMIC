module fake_jpeg_19158_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_22),
.Y(n_45)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_25),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_41),
.B(n_36),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_33),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_32),
.A2(n_28),
.B1(n_27),
.B2(n_15),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_32),
.B1(n_37),
.B2(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_34),
.B1(n_32),
.B2(n_37),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_59),
.B1(n_55),
.B2(n_47),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_34),
.B1(n_27),
.B2(n_28),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_60),
.A2(n_34),
.B1(n_47),
.B2(n_55),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_61),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_39),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_64),
.B(n_70),
.Y(n_85)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_43),
.B(n_21),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_32),
.B1(n_37),
.B2(n_33),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_43),
.B(n_21),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_81),
.Y(n_100)
);

NAND2x1_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_33),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_40),
.Y(n_106)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_82),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_84),
.A2(n_89),
.B(n_106),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_25),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_37),
.C(n_35),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_106),
.C(n_86),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_54),
.B1(n_72),
.B2(n_80),
.Y(n_121)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_108),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_105),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_40),
.Y(n_105)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_58),
.A2(n_17),
.B1(n_44),
.B2(n_54),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_109),
.A2(n_72),
.B1(n_76),
.B2(n_53),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_61),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_111),
.Y(n_115)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_75),
.B(n_82),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_114),
.A2(n_119),
.B(n_51),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_56),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_123),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_83),
.A2(n_76),
.B1(n_80),
.B2(n_44),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_108),
.B1(n_99),
.B2(n_53),
.Y(n_151)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_94),
.Y(n_123)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_127),
.A2(n_91),
.B1(n_51),
.B2(n_38),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_131),
.Y(n_168)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_92),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_100),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_19),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_132),
.B(n_135),
.Y(n_139)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_85),
.B(n_65),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_136),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_103),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_105),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_138),
.B(n_98),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_133),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_140),
.B(n_154),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_117),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_84),
.B(n_96),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_145),
.A2(n_149),
.B(n_159),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_166),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_113),
.A2(n_31),
.B(n_23),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_90),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_150),
.B(n_163),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_118),
.B1(n_128),
.B2(n_130),
.Y(n_176)
);

BUFx12_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_134),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_111),
.B1(n_90),
.B2(n_91),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_153),
.A2(n_165),
.B1(n_127),
.B2(n_123),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_125),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_155),
.A2(n_51),
.B1(n_38),
.B2(n_23),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_115),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_157),
.B(n_162),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g190 ( 
.A1(n_158),
.A2(n_149),
.B(n_145),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_26),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_115),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_31),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_17),
.B1(n_38),
.B2(n_56),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_112),
.B(n_30),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_112),
.B(n_40),
.C(n_56),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_51),
.C(n_22),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_40),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_23),
.B(n_26),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_178),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_172),
.A2(n_199),
.B1(n_202),
.B2(n_151),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_173),
.B(n_185),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_122),
.B1(n_120),
.B2(n_136),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_176),
.B1(n_170),
.B2(n_165),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_168),
.A2(n_135),
.B1(n_120),
.B2(n_132),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_182),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_142),
.B(n_116),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_181),
.B(n_191),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_129),
.Y(n_185)
);

AND2x6_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_120),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_166),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_156),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_188),
.B(n_189),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_30),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_190),
.A2(n_1),
.B(n_2),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_139),
.B(n_1),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_169),
.A2(n_30),
.B1(n_26),
.B2(n_20),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_193),
.A2(n_195),
.B(n_199),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_200),
.C(n_155),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_29),
.B1(n_24),
.B2(n_30),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_198),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_22),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_148),
.B(n_29),
.C(n_24),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_224),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_163),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_194),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_186),
.A2(n_161),
.B(n_143),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_206),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_183),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_220),
.B1(n_178),
.B2(n_200),
.Y(n_234)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_175),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_214),
.Y(n_231)
);

NOR3xp33_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_164),
.C(n_146),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_174),
.B(n_20),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_177),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_223),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_26),
.Y(n_225)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

XOR2x2_ASAP7_75t_SL g229 ( 
.A(n_224),
.B(n_190),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_229),
.B(n_246),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_243),
.Y(n_262)
);

XOR2x2_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_192),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_232),
.A2(n_218),
.B(n_205),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_180),
.B1(n_172),
.B2(n_171),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_238),
.A2(n_210),
.B1(n_218),
.B2(n_219),
.Y(n_250)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_187),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_198),
.B1(n_202),
.B2(n_196),
.Y(n_244)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_244),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_187),
.C(n_193),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_215),
.C(n_223),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_23),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_213),
.C(n_207),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_250),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_206),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_248),
.Y(n_271)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_253),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_254),
.B(n_256),
.Y(n_266)
);

OA21x2_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_216),
.B(n_219),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_246),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_215),
.C(n_212),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_259),
.C(n_260),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_217),
.C(n_209),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_2),
.C(n_3),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_2),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_261),
.A2(n_239),
.B(n_227),
.Y(n_265)
);

BUFx12_ASAP7_75t_L g263 ( 
.A(n_255),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_9),
.Y(n_288)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_265),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_243),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_270),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_251),
.A2(n_237),
.B1(n_236),
.B2(n_235),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_268),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_230),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_252),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_262),
.B(n_238),
.Y(n_270)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_272),
.Y(n_281)
);

BUFx12f_ASAP7_75t_SL g274 ( 
.A(n_258),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_274),
.A2(n_252),
.B(n_249),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_229),
.C(n_4),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_258),
.C(n_261),
.Y(n_277)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_270),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_3),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_284),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_4),
.B(n_5),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_4),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_10),
.B(n_11),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_276),
.B1(n_263),
.B2(n_13),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_6),
.C(n_9),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_288),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_296),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_271),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_286),
.B(n_277),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_279),
.B(n_264),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_297),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

AOI322xp5_ASAP7_75t_L g304 ( 
.A1(n_300),
.A2(n_302),
.A3(n_303),
.B1(n_292),
.B2(n_282),
.C1(n_268),
.C2(n_290),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_291),
.A2(n_285),
.B(n_263),
.Y(n_301)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_301),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_287),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_304),
.Y(n_307)
);

AOI321xp33_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_267),
.A3(n_282),
.B1(n_13),
.B2(n_14),
.C(n_11),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_307),
.A2(n_305),
.B(n_299),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_298),
.C(n_306),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_12),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_12),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_13),
.Y(n_313)
);


endmodule