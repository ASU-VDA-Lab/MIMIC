module real_jpeg_27925_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_333, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_332, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_333;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_332;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_0),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_92),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_0),
.A2(n_50),
.B1(n_52),
.B2(n_92),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_0),
.A2(n_55),
.B1(n_56),
.B2(n_92),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_1),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_1),
.A2(n_27),
.B1(n_50),
.B2(n_52),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_1),
.A2(n_27),
.B1(n_55),
.B2(n_56),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_2),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_107),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_107),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_2),
.A2(n_50),
.B1(n_52),
.B2(n_107),
.Y(n_200)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_3),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_4),
.B(n_50),
.Y(n_112)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_4),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_5),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_5),
.A2(n_45),
.B1(n_55),
.B2(n_56),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_45),
.Y(n_273)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_90),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_7),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_90),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_7),
.A2(n_55),
.B1(n_56),
.B2(n_90),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_7),
.A2(n_50),
.B1(n_52),
.B2(n_90),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_8),
.A2(n_55),
.B1(n_56),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_8),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_8),
.A2(n_50),
.B1(n_52),
.B2(n_100),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_100),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_100),
.Y(n_281)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_10),
.A2(n_36),
.B1(n_55),
.B2(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_10),
.A2(n_36),
.B1(n_50),
.B2(n_52),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_11),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_97),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_11),
.A2(n_50),
.B1(n_52),
.B2(n_97),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_97),
.Y(n_254)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_13),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_13),
.A2(n_29),
.B(n_33),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_13),
.B(n_31),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_13),
.A2(n_55),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_13),
.B(n_55),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_13),
.B(n_68),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_13),
.A2(n_115),
.B1(n_134),
.B2(n_200),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_13),
.A2(n_32),
.B(n_215),
.Y(n_214)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_16),
.A2(n_55),
.B1(n_56),
.B2(n_66),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_17),
.A2(n_43),
.B1(n_50),
.B2(n_52),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_17),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_43),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_78),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_76),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_21),
.B(n_37),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_23),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_29),
.Y(n_30)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_25),
.A2(n_34),
.B(n_104),
.C(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_31),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_28),
.A2(n_31),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_28),
.A2(n_31),
.B1(n_142),
.B2(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_28),
.A2(n_31),
.B1(n_161),
.B2(n_254),
.Y(n_253)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_31),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_32),
.A2(n_62),
.B(n_64),
.C(n_65),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_62),
.Y(n_64)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_32),
.A2(n_56),
.A3(n_62),
.B1(n_216),
.B2(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_33),
.B(n_104),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_69),
.C(n_71),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_38),
.A2(n_39),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_58),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_40),
.B(n_313),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_42),
.A2(n_73),
.B1(n_75),
.B2(n_281),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_46),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_46),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_46),
.A2(n_58),
.B1(n_307),
.B2(n_314),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_53),
.B(n_57),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_54),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_47),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_47),
.A2(n_53),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_47),
.A2(n_53),
.B1(n_132),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_47),
.A2(n_53),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_47),
.A2(n_53),
.B1(n_175),
.B2(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_47),
.B(n_104),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_47),
.A2(n_53),
.B1(n_96),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_47),
.A2(n_53),
.B1(n_57),
.B2(n_263),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

OAI32xp33_ASAP7_75t_L g177 ( 
.A1(n_48),
.A2(n_52),
.A3(n_55),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_49),
.B(n_50),
.Y(n_179)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_50),
.B(n_205),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_55),
.B(n_66),
.Y(n_224)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_58),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_59),
.A2(n_60),
.B1(n_68),
.B2(n_305),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_60),
.A2(n_68),
.B1(n_89),
.B2(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_60),
.A2(n_68),
.B1(n_145),
.B2(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_60),
.A2(n_68),
.B1(n_163),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_65),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_65),
.B1(n_88),
.B2(n_91),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_61),
.A2(n_65),
.B1(n_91),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_61),
.A2(n_65),
.B1(n_123),
.B2(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_61),
.A2(n_65),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_327),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_69),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_73),
.A2(n_75),
.B1(n_106),
.B2(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_73),
.A2(n_75),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_322),
.B(n_328),
.Y(n_78)
);

OAI321xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_298),
.A3(n_317),
.B1(n_320),
.B2(n_321),
.C(n_332),
.Y(n_79)
);

AOI321xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_250),
.A3(n_287),
.B1(n_292),
.B2(n_297),
.C(n_333),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_147),
.C(n_165),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_127),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_83),
.B(n_127),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_108),
.C(n_119),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_84),
.B(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_102),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_93),
.B2(n_94),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_86),
.B(n_94),
.C(n_102),
.Y(n_137)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_98),
.A2(n_101),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_98),
.A2(n_101),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_104),
.B(n_115),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_108),
.A2(n_119),
.B1(n_120),
.B2(n_248),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_108),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_111),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_118),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_112),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_112),
.A2(n_114),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_115),
.A2(n_134),
.B1(n_136),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_115),
.A2(n_134),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_115),
.A2(n_134),
.B1(n_194),
.B2(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_115),
.A2(n_134),
.B1(n_189),
.B2(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_115),
.A2(n_134),
.B(n_154),
.Y(n_265)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_126),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_121),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_124),
.B(n_126),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_125),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_138),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_137),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_137),
.C(n_138),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_133),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_146),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_143),
.C(n_146),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_148),
.A2(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_149),
.B(n_150),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_164),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_157),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_152),
.B(n_157),
.C(n_164),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_153),
.B(n_155),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_156),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_244),
.B(n_249),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_230),
.B(n_243),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_209),
.B(n_229),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_190),
.B(n_208),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_180),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_170),
.B(n_180),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_171),
.A2(n_172),
.B1(n_176),
.B2(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_174),
.Y(n_178)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_187),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_185),
.C(n_187),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_188),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_197),
.B(n_207),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_192),
.B(n_196),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_202),
.B(n_206),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_199),
.B(n_201),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_210),
.B(n_211),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_222),
.B1(n_227),
.B2(n_228),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_213),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_217),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_221),
.C(n_228),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_225),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_231),
.B(n_232),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_239),
.C(n_241),
.Y(n_245)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_238),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_246),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_267),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_267),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_258),
.C(n_266),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_252),
.B(n_258),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_252),
.Y(n_329)
);

FAx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.CI(n_257),
.CON(n_252),
.SN(n_252)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_255),
.C(n_257),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_254),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_256),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_264),
.B2(n_265),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_259),
.B(n_265),
.Y(n_283)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_265),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_264),
.A2(n_279),
.B(n_282),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_285),
.B2(n_286),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_276),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_270),
.B(n_276),
.C(n_286),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_274),
.B(n_275),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_274),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_273),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_300),
.C(n_309),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g319 ( 
.A(n_275),
.B(n_300),
.CI(n_309),
.CON(n_319),
.SN(n_319)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_276)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_277),
.Y(n_284)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_285),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_288),
.A2(n_293),
.B(n_296),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_289),
.B(n_290),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_310),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_310),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_308),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_301),
.A2(n_302),
.B1(n_312),
.B2(n_315),
.Y(n_311)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_304),
.C(n_307),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_315),
.C(n_316),
.Y(n_323)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_303),
.Y(n_308)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_304),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_316),
.Y(n_310)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_312),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_318),
.B(n_319),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_319),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);


endmodule