module fake_netlist_6_3655_n_4354 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_442, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_443, n_246, n_38, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_466, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_433, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_464, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_328, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4354);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_466;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_433;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_464;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_328;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4354;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_801;
wire n_3766;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_3783;
wire n_700;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_3844;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4168;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_509;
wire n_1342;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_677;
wire n_805;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1009;
wire n_1930;
wire n_1743;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_471;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4087;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_1371;
wire n_1285;
wire n_873;
wire n_2974;
wire n_2886;
wire n_3946;
wire n_1985;
wire n_4213;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_852;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_836;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_3979;
wire n_616;
wire n_658;
wire n_4308;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2739;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2510;
wire n_3023;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_4325;
wire n_2212;
wire n_3929;
wire n_758;
wire n_516;
wire n_3494;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_491;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_4187;
wire n_940;
wire n_770;
wire n_567;
wire n_1971;
wire n_1781;
wire n_2090;
wire n_2058;
wire n_2603;
wire n_2660;
wire n_538;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_494;
wire n_539;
wire n_493;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_1404;
wire n_638;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2551;
wire n_2364;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_4262;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_1815;
wire n_659;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_913;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4071;
wire n_4255;
wire n_3506;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_473;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_551;
wire n_699;
wire n_1986;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_564;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4349;
wire n_824;
wire n_686;
wire n_4102;
wire n_4297;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_577;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_619;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_572;
wire n_4314;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_1441;
wire n_606;
wire n_818;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_3910;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4296;
wire n_4009;
wire n_2633;
wire n_483;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_630;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_792;
wire n_2522;
wire n_476;
wire n_3949;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_982;
wire n_4257;
wire n_2674;
wire n_2832;
wire n_4226;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_932;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_3446;
wire n_4158;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_905;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_993;
wire n_2692;
wire n_3842;
wire n_689;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_966;
wire n_3888;
wire n_2908;
wire n_3168;
wire n_764;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4161;
wire n_4337;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3055;
wire n_3092;
wire n_3492;
wire n_3966;
wire n_3895;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_1014;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_882;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_586;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1950;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_702;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_835;
wire n_928;
wire n_1801;
wire n_850;
wire n_690;
wire n_1886;
wire n_1214;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_4043;
wire n_825;
wire n_4313;
wire n_728;
wire n_4353;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_515;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_696;
wire n_1515;
wire n_961;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_2824;
wire n_593;
wire n_4169;
wire n_514;
wire n_4055;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_3271;
wire n_950;
wire n_4248;
wire n_2812;
wire n_484;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_590;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_1052;
wire n_2794;
wire n_1033;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_3073;
wire n_2431;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_1634;
wire n_2078;
wire n_3252;
wire n_2932;
wire n_595;
wire n_1767;
wire n_627;
wire n_1779;
wire n_524;
wire n_1465;
wire n_3253;
wire n_3450;
wire n_3431;
wire n_3209;
wire n_4002;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_4289;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4288;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_495;
wire n_815;
wire n_3953;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_4191;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_639;
wire n_963;
wire n_2767;
wire n_794;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1139;
wire n_1714;
wire n_872;
wire n_3922;
wire n_3179;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_542;
wire n_847;
wire n_851;
wire n_644;
wire n_682;
wire n_2537;
wire n_2897;
wire n_3970;
wire n_4345;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_3171;
wire n_791;
wire n_1913;
wire n_4216;
wire n_3608;
wire n_510;
wire n_837;
wire n_4315;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_3353;
wire n_3150;
wire n_3018;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_765;
wire n_987;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2933;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_738;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_705;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_2134;
wire n_1176;
wire n_1004;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_3887;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_4123;
wire n_1431;
wire n_4096;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_4286;
wire n_1809;
wire n_3119;
wire n_4280;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_3731;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_4218;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_3557;
wire n_927;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_478;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4264;
wire n_2857;
wire n_3693;
wire n_3788;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_777;
wire n_1299;
wire n_2896;
wire n_526;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_4175;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_1507;
wire n_2482;
wire n_552;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_745;
wire n_1604;
wire n_2424;
wire n_2296;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_623;
wire n_716;
wire n_1201;
wire n_1398;
wire n_884;
wire n_2354;
wire n_2682;
wire n_1048;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_3393;
wire n_474;
wire n_811;
wire n_527;
wire n_1207;
wire n_683;
wire n_2442;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3451;
wire n_3480;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_2545;
wire n_3577;
wire n_3540;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_589;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_3641;
wire n_767;
wire n_3591;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_477;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1736;
wire n_1564;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_505;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_3944;
wire n_3909;
wire n_546;
wire n_1141;
wire n_562;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_3265;
wire n_2464;
wire n_2846;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_2329;
wire n_1092;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_511;
wire n_2990;
wire n_3847;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3323;
wire n_3226;
wire n_3364;
wire n_4020;
wire n_4176;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_4261;
wire n_1745;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_497;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1892;
wire n_1459;
wire n_1614;
wire n_3188;
wire n_3742;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4034;
wire n_1617;
wire n_4056;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_4206;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_4132;
wire n_2995;
wire n_2955;
wire n_1731;
wire n_2158;
wire n_3360;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_3917;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_3016;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2993;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_1129;
wire n_3870;
wire n_4030;
wire n_4126;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_664;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_607;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3276;
wire n_3194;
wire n_1934;
wire n_3250;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_617;
wire n_3886;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_4234;
wire n_4304;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_517;
wire n_4211;
wire n_4182;
wire n_3337;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_1037;
wire n_621;
wire n_1397;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_923;
wire n_504;
wire n_1409;
wire n_4230;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_4274;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4270;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_4155;
wire n_2740;
wire n_746;
wire n_4238;
wire n_1601;
wire n_609;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4109;
wire n_4192;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4159;
wire n_4195;
wire n_3784;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_1870;
wire n_2964;
wire n_4174;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_662;
wire n_3475;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_711;
wire n_1352;
wire n_579;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_4258;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_972;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3988;
wire n_1974;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_482;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3439;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_4135;
wire n_2871;
wire n_4209;
wire n_4279;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_3858;
wire n_4183;
wire n_1489;
wire n_4321;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_543;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_4040;
wire n_804;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_799;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_3007;
wire n_2809;
wire n_787;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_4343;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_652;
wire n_2154;
wire n_2727;
wire n_3377;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1914;
wire n_1318;
wire n_737;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_3762;
wire n_3469;
wire n_3958;
wire n_2266;
wire n_2960;
wire n_3932;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_502;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_655;
wire n_1045;
wire n_1650;
wire n_1794;
wire n_786;
wire n_1962;
wire n_1236;
wire n_706;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_4317;
wire n_834;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_743;
wire n_766;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2923;
wire n_2793;
wire n_2715;
wire n_2888;
wire n_1804;
wire n_2885;
wire n_3711;
wire n_3776;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4170;
wire n_4143;
wire n_729;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_841;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3458;
wire n_3216;
wire n_3515;
wire n_1150;
wire n_4203;
wire n_3808;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1929;
wire n_1007;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_853;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_680;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2163;
wire n_2186;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_2969;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_4295;
wire n_1120;
wire n_832;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_691;
wire n_535;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_1147;
wire n_1785;
wire n_763;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_4352;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_1303;
wire n_761;
wire n_2769;
wire n_4342;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_3062;
wire n_2858;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_4106;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4027;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_647;
wire n_4160;
wire n_4231;
wire n_844;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_1028;
wire n_576;
wire n_3836;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_2744;
wire n_4309;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_2743;
wire n_3962;
wire n_708;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_4166;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_498;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4142;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3697;
wire n_3643;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_492;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_719;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4105;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_4244;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_829;
wire n_1156;
wire n_1362;
wire n_4259;
wire n_3123;
wire n_984;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_859;
wire n_570;
wire n_2033;
wire n_3086;
wire n_735;
wire n_4104;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_3285;
wire n_519;
wire n_4208;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_4346;
wire n_4351;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_4316;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_3101;
wire n_2844;
wire n_3989;
wire n_756;
wire n_2478;
wire n_1619;
wire n_2303;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_1606;
wire n_4332;
wire n_810;
wire n_4108;
wire n_1133;
wire n_635;
wire n_1194;
wire n_3374;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_4051;
wire n_1051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_4293;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_3709;
wire n_753;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_4148;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_679;
wire n_4057;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_633;
wire n_1629;
wire n_1170;
wire n_665;
wire n_2221;
wire n_588;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1890;
wire n_1632;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_3903;
wire n_730;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_640;
wire n_4129;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3584;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_629;
wire n_4275;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_900;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_531;
wire n_827;
wire n_2912;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g469 ( 
.A(n_213),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_119),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_403),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_365),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_462),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_166),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_0),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_260),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_283),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_167),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_133),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_236),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_69),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_321),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_439),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_366),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_218),
.Y(n_485)
);

BUFx8_ASAP7_75t_SL g486 ( 
.A(n_220),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_348),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_177),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_50),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_413),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_294),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_404),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_69),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_10),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_323),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_437),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_447),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_425),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_1),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_123),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_285),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_47),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_397),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_197),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_182),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_146),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_50),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_220),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_364),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_434),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_385),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_428),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_0),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_151),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_386),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_158),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_261),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_159),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_175),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_29),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_57),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_370),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_110),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_130),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_157),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_49),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_61),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_153),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_267),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_287),
.Y(n_530)
);

BUFx5_ASAP7_75t_L g531 ( 
.A(n_320),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_81),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_2),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_85),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_102),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_8),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_357),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_143),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_8),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_358),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_114),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_368),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_126),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_117),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_254),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_316),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_5),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_332),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_241),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_30),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_66),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_174),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_416),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_334),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_420),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_66),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_419),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_34),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_188),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_251),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_165),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_400),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_174),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_231),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_401),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_461),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_294),
.Y(n_567)
);

BUFx8_ASAP7_75t_SL g568 ( 
.A(n_367),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_168),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_103),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_291),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_143),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_433),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_375),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_291),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_73),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_232),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_339),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_282),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_331),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_109),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_173),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_429),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_31),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_426),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_446),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_309),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_173),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_105),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_167),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_326),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_47),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_19),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_25),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_305),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_318),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_298),
.Y(n_597)
);

BUFx10_ASAP7_75t_L g598 ( 
.A(n_86),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_39),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_261),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_242),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_249),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_276),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_40),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_252),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_309),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_307),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_215),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_20),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_93),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_353),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_417),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_181),
.Y(n_613)
);

BUFx5_ASAP7_75t_L g614 ( 
.A(n_226),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_211),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_82),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_249),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_239),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_381),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_184),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_228),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_436),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_467),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_86),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_74),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_112),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_122),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_456),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_17),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_77),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_125),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_346),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_377),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_77),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_243),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_231),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_359),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_49),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_117),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_103),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_390),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_247),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_376),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_124),
.Y(n_644)
);

CKINVDCx16_ASAP7_75t_R g645 ( 
.A(n_79),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_27),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_138),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_13),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_411),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_338),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_5),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_300),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_179),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_120),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_412),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_222),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_186),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_168),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_171),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_121),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_123),
.Y(n_661)
);

CKINVDCx14_ASAP7_75t_R g662 ( 
.A(n_93),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_341),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_324),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_155),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_209),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_297),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_197),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_333),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_28),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_289),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_24),
.Y(n_672)
);

BUFx5_ASAP7_75t_L g673 ( 
.A(n_256),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_137),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_265),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_153),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_144),
.Y(n_677)
);

BUFx10_ASAP7_75t_L g678 ( 
.A(n_306),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_180),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_243),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_290),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_169),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_105),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_62),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_115),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_219),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_48),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_345),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_107),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_405),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_126),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_10),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_92),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_11),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_111),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_435),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_95),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_101),
.Y(n_698)
);

CKINVDCx16_ASAP7_75t_R g699 ( 
.A(n_239),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_170),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_340),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_424),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_328),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_391),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_11),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_111),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_432),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_374),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_459),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_454),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_45),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_292),
.Y(n_712)
);

BUFx10_ASAP7_75t_L g713 ( 
.A(n_254),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_360),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_194),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_236),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_260),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_115),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_179),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_205),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_444),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_15),
.Y(n_722)
);

BUFx10_ASAP7_75t_L g723 ( 
.A(n_292),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_7),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_43),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_245),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_139),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_269),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_61),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_9),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_113),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_65),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_312),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_269),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_233),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_90),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_181),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_2),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_166),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_369),
.Y(n_740)
);

INVxp67_ASAP7_75t_SL g741 ( 
.A(n_282),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_125),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_70),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_297),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_20),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_90),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_35),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_289),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_351),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_319),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_183),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_361),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_352),
.Y(n_753)
);

CKINVDCx16_ASAP7_75t_R g754 ( 
.A(n_194),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_350),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_449),
.Y(n_756)
);

INVx4_ASAP7_75t_R g757 ( 
.A(n_296),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_177),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_427),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_164),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_267),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_414),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_238),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_204),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_187),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_290),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_300),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_531),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_495),
.Y(n_769)
);

INVxp67_ASAP7_75t_SL g770 ( 
.A(n_495),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_531),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_497),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_510),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_531),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_531),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_531),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_531),
.Y(n_777)
);

CKINVDCx16_ASAP7_75t_R g778 ( 
.A(n_618),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_531),
.Y(n_779)
);

CKINVDCx16_ASAP7_75t_R g780 ( 
.A(n_618),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_531),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_531),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_486),
.Y(n_783)
);

INVxp67_ASAP7_75t_SL g784 ( 
.A(n_497),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_614),
.Y(n_785)
);

CKINVDCx14_ASAP7_75t_R g786 ( 
.A(n_662),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_598),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_614),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_614),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_614),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_614),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_614),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_614),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_568),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_614),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_614),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_673),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_673),
.B(n_1),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_673),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_673),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_673),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_673),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_645),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_673),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_673),
.Y(n_805)
);

INVxp33_ASAP7_75t_SL g806 ( 
.A(n_685),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_739),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_573),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_673),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_481),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_573),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_481),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_481),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_481),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_481),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_594),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_594),
.Y(n_817)
);

CKINVDCx16_ASAP7_75t_R g818 ( 
.A(n_645),
.Y(n_818)
);

INVxp67_ASAP7_75t_SL g819 ( 
.A(n_574),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_594),
.Y(n_820)
);

INVxp33_ASAP7_75t_L g821 ( 
.A(n_739),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_594),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_594),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_599),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_599),
.Y(n_825)
);

BUFx2_ASAP7_75t_SL g826 ( 
.A(n_619),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_699),
.Y(n_827)
);

CKINVDCx16_ASAP7_75t_R g828 ( 
.A(n_699),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_599),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_599),
.Y(n_830)
);

CKINVDCx16_ASAP7_75t_R g831 ( 
.A(n_754),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_599),
.Y(n_832)
);

INVxp33_ASAP7_75t_SL g833 ( 
.A(n_475),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_676),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_676),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_676),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_676),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_471),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_471),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_509),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_469),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_509),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_522),
.Y(n_843)
);

CKINVDCx16_ASAP7_75t_R g844 ( 
.A(n_754),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_522),
.Y(n_845)
);

NOR2xp67_ASAP7_75t_L g846 ( 
.A(n_557),
.B(n_3),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_622),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_622),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_676),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_628),
.Y(n_850)
);

INVxp67_ASAP7_75t_SL g851 ( 
.A(n_574),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_628),
.Y(n_852)
);

INVxp33_ASAP7_75t_L g853 ( 
.A(n_469),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_632),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_632),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_472),
.Y(n_856)
);

CKINVDCx16_ASAP7_75t_R g857 ( 
.A(n_598),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_720),
.Y(n_858)
);

INVxp33_ASAP7_75t_L g859 ( 
.A(n_478),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_485),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_664),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_477),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_664),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_669),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_669),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_688),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_688),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_701),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_507),
.Y(n_869)
);

INVxp67_ASAP7_75t_SL g870 ( 
.A(n_637),
.Y(n_870)
);

INVxp67_ASAP7_75t_SL g871 ( 
.A(n_637),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_701),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_703),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_703),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_720),
.Y(n_875)
);

INVxp33_ASAP7_75t_SL g876 ( 
.A(n_479),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_710),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_473),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_720),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_720),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_548),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_480),
.Y(n_882)
);

INVxp33_ASAP7_75t_SL g883 ( 
.A(n_482),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_720),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_474),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_474),
.Y(n_886)
);

INVxp67_ASAP7_75t_SL g887 ( 
.A(n_710),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_476),
.Y(n_888)
);

INVxp67_ASAP7_75t_SL g889 ( 
.A(n_557),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_494),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_476),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_518),
.Y(n_892)
);

CKINVDCx16_ASAP7_75t_R g893 ( 
.A(n_598),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_483),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_518),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_478),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_484),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_672),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_672),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_707),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_489),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_489),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_499),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_487),
.Y(n_904)
);

INVxp33_ASAP7_75t_L g905 ( 
.A(n_491),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_491),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_530),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_508),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_508),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_513),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_501),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_513),
.Y(n_912)
);

INVxp67_ASAP7_75t_L g913 ( 
.A(n_516),
.Y(n_913)
);

INVxp33_ASAP7_75t_SL g914 ( 
.A(n_502),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_516),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_504),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_521),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_521),
.Y(n_918)
);

INVx4_ASAP7_75t_R g919 ( 
.A(n_619),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_771),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_881),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_770),
.B(n_520),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_771),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_889),
.B(n_557),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_784),
.B(n_752),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_846),
.B(n_752),
.Y(n_926)
);

INVx5_ASAP7_75t_L g927 ( 
.A(n_881),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_849),
.B(n_623),
.Y(n_928)
);

BUFx12f_ASAP7_75t_L g929 ( 
.A(n_783),
.Y(n_929)
);

INVx5_ASAP7_75t_L g930 ( 
.A(n_881),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_796),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_881),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_806),
.A2(n_546),
.B1(n_600),
.B2(n_547),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_810),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_810),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_812),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_812),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_803),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_803),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_857),
.B(n_583),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_769),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_796),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_881),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_801),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_801),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_890),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_808),
.B(n_520),
.Y(n_947)
);

BUFx8_ASAP7_75t_SL g948 ( 
.A(n_794),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_849),
.B(n_623),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_827),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_858),
.Y(n_951)
);

OAI21x1_ASAP7_75t_L g952 ( 
.A1(n_809),
.A2(n_696),
.B(n_655),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_809),
.Y(n_953)
);

OA21x2_ASAP7_75t_L g954 ( 
.A1(n_798),
.A2(n_709),
.B(n_707),
.Y(n_954)
);

INVx5_ASAP7_75t_L g955 ( 
.A(n_858),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_827),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_768),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_774),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_774),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_813),
.Y(n_960)
);

BUFx8_ASAP7_75t_SL g961 ( 
.A(n_783),
.Y(n_961)
);

OA21x2_ASAP7_75t_L g962 ( 
.A1(n_775),
.A2(n_721),
.B(n_709),
.Y(n_962)
);

INVx5_ASAP7_75t_L g963 ( 
.A(n_900),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_862),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_862),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_819),
.B(n_490),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_813),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_833),
.B(n_914),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_851),
.B(n_870),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_814),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_786),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_814),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_871),
.B(n_655),
.Y(n_973)
);

BUFx12f_ASAP7_75t_L g974 ( 
.A(n_882),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_856),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_815),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_775),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_876),
.B(n_762),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_815),
.Y(n_979)
);

CKINVDCx14_ASAP7_75t_R g980 ( 
.A(n_773),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_877),
.B(n_696),
.Y(n_981)
);

INVxp67_ASAP7_75t_L g982 ( 
.A(n_807),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_816),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_776),
.Y(n_984)
);

INVxp33_ASAP7_75t_SL g985 ( 
.A(n_882),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_769),
.Y(n_986)
);

AOI22x1_ASAP7_75t_SL g987 ( 
.A1(n_860),
.A2(n_626),
.B1(n_635),
.B2(n_630),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_776),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_777),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_787),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_777),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_772),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_779),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_816),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_817),
.B(n_820),
.Y(n_995)
);

INVx5_ASAP7_75t_L g996 ( 
.A(n_900),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_817),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_903),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_820),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_779),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_887),
.B(n_532),
.Y(n_1001)
);

OAI22x1_ASAP7_75t_R g1002 ( 
.A1(n_778),
.A2(n_666),
.B1(n_691),
.B2(n_653),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_878),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_822),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_822),
.Y(n_1005)
);

INVx5_ASAP7_75t_L g1006 ( 
.A(n_772),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_823),
.Y(n_1007)
);

AND2x6_ASAP7_75t_L g1008 ( 
.A(n_781),
.B(n_548),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_811),
.B(n_826),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_823),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_824),
.Y(n_1011)
);

BUFx8_ASAP7_75t_SL g1012 ( 
.A(n_903),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_824),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_825),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_781),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_825),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_782),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_826),
.B(n_492),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_782),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_883),
.B(n_721),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_785),
.Y(n_1021)
);

INVx6_ASAP7_75t_L g1022 ( 
.A(n_811),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_785),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_829),
.B(n_496),
.Y(n_1024)
);

NAND2xp33_ASAP7_75t_L g1025 ( 
.A(n_911),
.B(n_505),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_829),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_780),
.A2(n_728),
.B1(n_717),
.B2(n_731),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_818),
.A2(n_828),
.B1(n_844),
.B2(n_831),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_830),
.B(n_753),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_853),
.B(n_532),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_788),
.Y(n_1031)
);

AND2x2_ASAP7_75t_SL g1032 ( 
.A(n_838),
.B(n_548),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_830),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_788),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_789),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_832),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_832),
.B(n_755),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_834),
.B(n_498),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_SL g1039 ( 
.A1(n_869),
.A2(n_603),
.B1(n_533),
.B2(n_536),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_834),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_835),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_835),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_836),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_836),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_837),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_911),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_837),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_875),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_789),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_1012),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1009),
.B(n_875),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_920),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_969),
.B(n_894),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1036),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1009),
.B(n_879),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1036),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1036),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1041),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_1030),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1041),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_924),
.B(n_879),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1041),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_920),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_957),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_975),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_920),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_1003),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_924),
.B(n_880),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_974),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_957),
.Y(n_1070)
);

AND2x6_ASAP7_75t_L g1071 ( 
.A(n_924),
.B(n_926),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_1028),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_923),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_974),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_1030),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_923),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_974),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_921),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_1028),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_923),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_924),
.B(n_880),
.Y(n_1081)
);

CKINVDCx8_ASAP7_75t_R g1082 ( 
.A(n_939),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_R g1083 ( 
.A(n_980),
.B(n_897),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_957),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_941),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_931),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_989),
.Y(n_1087)
);

NOR2xp67_ASAP7_75t_L g1088 ( 
.A(n_964),
.B(n_916),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_933),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_R g1090 ( 
.A(n_1025),
.B(n_904),
.Y(n_1090)
);

OA21x2_ASAP7_75t_L g1091 ( 
.A1(n_952),
.A2(n_791),
.B(n_790),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_990),
.B(n_787),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_921),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_941),
.B(n_986),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_961),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_971),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_986),
.B(n_821),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_921),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_989),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_971),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_948),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_985),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_989),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_939),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_966),
.B(n_884),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_929),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_929),
.Y(n_1107)
);

AND2x6_ASAP7_75t_L g1108 ( 
.A(n_926),
.B(n_753),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_921),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_989),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_SL g1111 ( 
.A(n_968),
.B(n_893),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1031),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_921),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_931),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_966),
.B(n_884),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_933),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1032),
.B(n_790),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_929),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1031),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_931),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_950),
.Y(n_1121)
);

XNOR2xp5_ASAP7_75t_L g1122 ( 
.A(n_1027),
.B(n_907),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_1002),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1031),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_978),
.B(n_916),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_992),
.B(n_859),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_992),
.B(n_905),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_921),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_932),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1031),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_928),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_950),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_1002),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_928),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_932),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1032),
.B(n_791),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_932),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_928),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_1046),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1046),
.Y(n_1140)
);

NAND2xp33_ASAP7_75t_R g1141 ( 
.A(n_922),
.B(n_506),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_928),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_942),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_949),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_949),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_987),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_1027),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1032),
.B(n_792),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_941),
.B(n_1029),
.Y(n_1149)
);

BUFx10_ASAP7_75t_L g1150 ( 
.A(n_1020),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_949),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_938),
.Y(n_1152)
);

INVxp67_ASAP7_75t_SL g1153 ( 
.A(n_1038),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_956),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_987),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_965),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_942),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_932),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_932),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_949),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_926),
.B(n_792),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_995),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_998),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_995),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_946),
.A2(n_741),
.B1(n_493),
.B2(n_517),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_995),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_982),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1029),
.B(n_839),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_942),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_932),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_995),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_958),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_944),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1029),
.B(n_840),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1039),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_1039),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_940),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_943),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_944),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_922),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_943),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_958),
.Y(n_1182)
);

CKINVDCx20_ASAP7_75t_R g1183 ( 
.A(n_947),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_947),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1018),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_958),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_1001),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1001),
.B(n_925),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_1022),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_944),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_959),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1022),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1022),
.Y(n_1193)
);

AND2x2_ASAP7_75t_SL g1194 ( 
.A(n_926),
.B(n_548),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1022),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_959),
.Y(n_1196)
);

BUFx8_ASAP7_75t_L g1197 ( 
.A(n_1029),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_959),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_945),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1022),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_973),
.B(n_841),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_943),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_981),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_945),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1038),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1006),
.B(n_583),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1006),
.B(n_583),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_945),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1006),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_977),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_953),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1006),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1006),
.B(n_896),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_943),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1006),
.B(n_583),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_953),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_977),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_977),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_984),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_943),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1024),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1037),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_953),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_952),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_934),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_984),
.Y(n_1226)
);

NAND2xp33_ASAP7_75t_R g1227 ( 
.A(n_954),
.B(n_514),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_954),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_984),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_988),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_943),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_988),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_951),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_954),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_951),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_934),
.B(n_842),
.Y(n_1236)
);

INVxp67_ASAP7_75t_SL g1237 ( 
.A(n_951),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_988),
.B(n_793),
.Y(n_1238)
);

OA21x2_ASAP7_75t_L g1239 ( 
.A1(n_935),
.A2(n_795),
.B(n_793),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_954),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_935),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_936),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_991),
.Y(n_1243)
);

AND2x6_ASAP7_75t_L g1244 ( 
.A(n_991),
.B(n_548),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_951),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_951),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_951),
.Y(n_1247)
);

BUFx10_ASAP7_75t_L g1248 ( 
.A(n_1008),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_962),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_936),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_991),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_962),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_937),
.Y(n_1253)
);

CKINVDCx8_ASAP7_75t_R g1254 ( 
.A(n_962),
.Y(n_1254)
);

BUFx10_ASAP7_75t_L g1255 ( 
.A(n_1008),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_993),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_962),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_993),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_993),
.Y(n_1259)
);

BUFx8_ASAP7_75t_L g1260 ( 
.A(n_937),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1000),
.B(n_708),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1000),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1000),
.Y(n_1263)
);

INVxp67_ASAP7_75t_L g1264 ( 
.A(n_960),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1015),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1015),
.B(n_795),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_960),
.B(n_901),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_970),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1015),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1017),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_970),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_983),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1017),
.Y(n_1273)
);

AND2x6_ASAP7_75t_L g1274 ( 
.A(n_1017),
.B(n_663),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_967),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_983),
.B(n_843),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1019),
.A2(n_799),
.B(n_797),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_1147),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1149),
.B(n_902),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1131),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1224),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1188),
.B(n_913),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1224),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1134),
.Y(n_1284)
);

NAND2xp33_ASAP7_75t_L g1285 ( 
.A(n_1071),
.B(n_663),
.Y(n_1285)
);

NAND2xp33_ASAP7_75t_SL g1286 ( 
.A(n_1177),
.B(n_470),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1050),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1205),
.B(n_503),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1277),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1059),
.B(n_1184),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1205),
.B(n_511),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1138),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1277),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1071),
.A2(n_1019),
.B1(n_1023),
.B2(n_1021),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1126),
.B(n_845),
.Y(n_1295)
);

NAND3xp33_ASAP7_75t_L g1296 ( 
.A(n_1187),
.B(n_523),
.C(n_519),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1149),
.B(n_902),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1239),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1239),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1053),
.B(n_524),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1239),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1221),
.B(n_512),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1094),
.Y(n_1303)
);

INVx4_ASAP7_75t_L g1304 ( 
.A(n_1071),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1142),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1185),
.B(n_1221),
.Y(n_1306)
);

NAND3xp33_ASAP7_75t_L g1307 ( 
.A(n_1141),
.B(n_526),
.C(n_525),
.Y(n_1307)
);

NAND2xp33_ASAP7_75t_SL g1308 ( 
.A(n_1177),
.B(n_470),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_1127),
.Y(n_1309)
);

BUFx4f_ASAP7_75t_L g1310 ( 
.A(n_1071),
.Y(n_1310)
);

INVx4_ASAP7_75t_L g1311 ( 
.A(n_1071),
.Y(n_1311)
);

AND3x2_ASAP7_75t_L g1312 ( 
.A(n_1111),
.B(n_533),
.C(n_529),
.Y(n_1312)
);

AND3x2_ASAP7_75t_L g1313 ( 
.A(n_1104),
.B(n_536),
.C(n_529),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1075),
.B(n_906),
.Y(n_1314)
);

INVxp33_ASAP7_75t_L g1315 ( 
.A(n_1122),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1144),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1052),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1052),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1063),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1063),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1097),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1066),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1145),
.Y(n_1323)
);

OR2x2_ASAP7_75t_SL g1324 ( 
.A(n_1167),
.B(n_561),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1151),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1249),
.A2(n_537),
.B1(n_540),
.B2(n_515),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1222),
.B(n_1125),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1066),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1222),
.B(n_1150),
.Y(n_1329)
);

INVx4_ASAP7_75t_L g1330 ( 
.A(n_1071),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1073),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1153),
.B(n_1019),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1073),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1150),
.B(n_527),
.Y(n_1334)
);

OAI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1249),
.A2(n_500),
.B1(n_604),
.B2(n_488),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1076),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1160),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1257),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1162),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1076),
.Y(n_1340)
);

INVxp67_ASAP7_75t_SL g1341 ( 
.A(n_1275),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1105),
.B(n_1021),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1201),
.B(n_847),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1115),
.B(n_1021),
.Y(n_1344)
);

INVx4_ASAP7_75t_L g1345 ( 
.A(n_1189),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1164),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1166),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1180),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1149),
.B(n_906),
.Y(n_1349)
);

OR2x6_ASAP7_75t_L g1350 ( 
.A(n_1094),
.B(n_488),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1092),
.B(n_1094),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1150),
.B(n_528),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1088),
.B(n_542),
.Y(n_1353)
);

OAI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1252),
.A2(n_604),
.B1(n_621),
.B2(n_500),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1194),
.B(n_1023),
.Y(n_1355)
);

NAND2xp33_ASAP7_75t_L g1356 ( 
.A(n_1252),
.B(n_663),
.Y(n_1356)
);

INVx5_ASAP7_75t_L g1357 ( 
.A(n_1248),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1171),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1225),
.B(n_848),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1080),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1194),
.B(n_1023),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1080),
.Y(n_1362)
);

BUFx4f_ASAP7_75t_L g1363 ( 
.A(n_1108),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1225),
.B(n_850),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1117),
.A2(n_1034),
.B1(n_1049),
.B2(n_1035),
.Y(n_1365)
);

NAND3xp33_ASAP7_75t_L g1366 ( 
.A(n_1242),
.B(n_535),
.C(n_534),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1091),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1061),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1068),
.Y(n_1369)
);

NAND3xp33_ASAP7_75t_L g1370 ( 
.A(n_1242),
.B(n_539),
.C(n_538),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1085),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1180),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1086),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1267),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1091),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1051),
.B(n_1034),
.Y(n_1376)
);

XOR2x2_ASAP7_75t_L g1377 ( 
.A(n_1165),
.B(n_3),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1086),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1114),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1091),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1081),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1087),
.Y(n_1382)
);

NAND3xp33_ASAP7_75t_L g1383 ( 
.A(n_1250),
.B(n_543),
.C(n_541),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1250),
.B(n_852),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1114),
.Y(n_1385)
);

BUFx10_ASAP7_75t_L g1386 ( 
.A(n_1101),
.Y(n_1386)
);

BUFx4f_ASAP7_75t_L g1387 ( 
.A(n_1108),
.Y(n_1387)
);

CKINVDCx11_ASAP7_75t_R g1388 ( 
.A(n_1123),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1253),
.B(n_854),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1136),
.A2(n_1034),
.B1(n_1049),
.B2(n_1035),
.Y(n_1390)
);

INVx5_ASAP7_75t_L g1391 ( 
.A(n_1248),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1120),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1257),
.Y(n_1393)
);

NAND2xp33_ASAP7_75t_L g1394 ( 
.A(n_1148),
.B(n_663),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1099),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1120),
.Y(n_1396)
);

INVx4_ASAP7_75t_L g1397 ( 
.A(n_1189),
.Y(n_1397)
);

NAND2xp33_ASAP7_75t_R g1398 ( 
.A(n_1139),
.B(n_553),
.Y(n_1398)
);

AND3x1_ASAP7_75t_L g1399 ( 
.A(n_1241),
.B(n_567),
.C(n_561),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1253),
.B(n_855),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1183),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1203),
.B(n_544),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1192),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1143),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1143),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_SL g1406 ( 
.A(n_1268),
.B(n_554),
.Y(n_1406)
);

INVx4_ASAP7_75t_L g1407 ( 
.A(n_1192),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1234),
.A2(n_1035),
.B1(n_1049),
.B2(n_1008),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1157),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1157),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1103),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1169),
.Y(n_1412)
);

INVxp33_ASAP7_75t_L g1413 ( 
.A(n_1083),
.Y(n_1413)
);

OR2x6_ASAP7_75t_L g1414 ( 
.A(n_1055),
.B(n_621),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1110),
.Y(n_1415)
);

NAND3xp33_ASAP7_75t_L g1416 ( 
.A(n_1268),
.B(n_549),
.C(n_545),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1254),
.Y(n_1417)
);

INVxp33_ASAP7_75t_L g1418 ( 
.A(n_1090),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1271),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1169),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1161),
.B(n_994),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1054),
.B(n_994),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1112),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1197),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1119),
.Y(n_1425)
);

AND3x2_ASAP7_75t_L g1426 ( 
.A(n_1272),
.B(n_575),
.C(n_567),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_SL g1427 ( 
.A(n_1271),
.B(n_555),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1124),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1254),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1168),
.B(n_861),
.Y(n_1430)
);

AND2x6_ASAP7_75t_L g1431 ( 
.A(n_1130),
.B(n_663),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1056),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1248),
.Y(n_1433)
);

NAND3xp33_ASAP7_75t_L g1434 ( 
.A(n_1227),
.B(n_551),
.C(n_550),
.Y(n_1434)
);

NAND3xp33_ASAP7_75t_L g1435 ( 
.A(n_1264),
.B(n_556),
.C(n_552),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_1168),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1183),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1173),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1057),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1197),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1058),
.B(n_997),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1168),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1203),
.B(n_558),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1060),
.B(n_997),
.Y(n_1444)
);

NOR3xp33_ASAP7_75t_L g1445 ( 
.A(n_1139),
.B(n_758),
.C(n_750),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1062),
.B(n_1174),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1226),
.Y(n_1447)
);

INVx6_ASAP7_75t_L g1448 ( 
.A(n_1197),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1226),
.Y(n_1449)
);

INVx5_ASAP7_75t_L g1450 ( 
.A(n_1255),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1251),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_SL g1452 ( 
.A(n_1174),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1251),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1174),
.B(n_863),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1173),
.Y(n_1455)
);

BUFx10_ASAP7_75t_L g1456 ( 
.A(n_1101),
.Y(n_1456)
);

NOR2x1p5_ASAP7_75t_L g1457 ( 
.A(n_1069),
.B(n_576),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1179),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1179),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1259),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1228),
.A2(n_565),
.B1(n_566),
.B2(n_562),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1193),
.B(n_578),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1102),
.B(n_559),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1193),
.B(n_1195),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1240),
.A2(n_1008),
.B1(n_799),
.B2(n_800),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1050),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1228),
.A2(n_585),
.B1(n_586),
.B2(n_580),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1195),
.B(n_591),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1259),
.Y(n_1469)
);

INVx1_ASAP7_75t_SL g1470 ( 
.A(n_1140),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1190),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1121),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1269),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1200),
.B(n_999),
.Y(n_1474)
);

INVx4_ASAP7_75t_L g1475 ( 
.A(n_1200),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_1147),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1102),
.B(n_1156),
.Y(n_1477)
);

INVx2_ASAP7_75t_SL g1478 ( 
.A(n_1213),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1255),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1269),
.Y(n_1480)
);

NAND3xp33_ASAP7_75t_L g1481 ( 
.A(n_1175),
.B(n_563),
.C(n_560),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1273),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1245),
.B(n_999),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1140),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1273),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1108),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1108),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1190),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1199),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1199),
.Y(n_1490)
);

INVx1_ASAP7_75t_SL g1491 ( 
.A(n_1121),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1108),
.A2(n_1008),
.B1(n_800),
.B2(n_802),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1204),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1108),
.A2(n_612),
.B1(n_633),
.B2(n_611),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1156),
.B(n_564),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1246),
.A2(n_643),
.B1(n_649),
.B2(n_641),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1163),
.B(n_650),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1204),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1208),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1163),
.B(n_569),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1261),
.B(n_908),
.Y(n_1501)
);

AND3x2_ASAP7_75t_L g1502 ( 
.A(n_1236),
.B(n_581),
.C(n_575),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1206),
.A2(n_1215),
.B1(n_1207),
.B2(n_1276),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1208),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1064),
.A2(n_1008),
.B1(n_802),
.B2(n_804),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1211),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1211),
.Y(n_1507)
);

BUFx8_ASAP7_75t_SL g1508 ( 
.A(n_1095),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1216),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1216),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1223),
.B(n_864),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1223),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1132),
.B(n_570),
.Y(n_1513)
);

NAND2xp33_ASAP7_75t_L g1514 ( 
.A(n_1244),
.B(n_1008),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1070),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1235),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1132),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1082),
.B(n_690),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1082),
.B(n_865),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1084),
.A2(n_1008),
.B1(n_804),
.B2(n_805),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1172),
.A2(n_805),
.B1(n_797),
.B2(n_758),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1289),
.Y(n_1522)
);

INVx4_ASAP7_75t_SL g1523 ( 
.A(n_1338),
.Y(n_1523)
);

AND2x6_ASAP7_75t_L g1524 ( 
.A(n_1338),
.B(n_1393),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1303),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_SL g1526 ( 
.A1(n_1327),
.A2(n_1116),
.B1(n_1089),
.B2(n_1176),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1290),
.B(n_1175),
.Y(n_1527)
);

AO22x2_ASAP7_75t_L g1528 ( 
.A1(n_1419),
.A2(n_750),
.B1(n_581),
.B2(n_587),
.Y(n_1528)
);

NAND2x1p5_ASAP7_75t_L g1529 ( 
.A(n_1338),
.B(n_1235),
.Y(n_1529)
);

OR2x2_ASAP7_75t_SL g1530 ( 
.A(n_1401),
.B(n_1176),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1338),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1339),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1303),
.B(n_1235),
.Y(n_1533)
);

OAI22x1_ASAP7_75t_L g1534 ( 
.A1(n_1419),
.A2(n_1067),
.B1(n_1065),
.B2(n_1146),
.Y(n_1534)
);

INVx8_ASAP7_75t_L g1535 ( 
.A(n_1452),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1289),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1339),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1346),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1282),
.B(n_1065),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1371),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1300),
.B(n_1182),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1346),
.Y(n_1542)
);

NAND3xp33_ASAP7_75t_L g1543 ( 
.A(n_1306),
.B(n_1067),
.C(n_1096),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1338),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1393),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1371),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1282),
.B(n_1096),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1293),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1293),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1436),
.B(n_1247),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1359),
.B(n_1100),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1347),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1393),
.Y(n_1553)
);

NAND2xp33_ASAP7_75t_SL g1554 ( 
.A(n_1393),
.B(n_1100),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1436),
.B(n_1247),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1442),
.B(n_1247),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1359),
.B(n_1069),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1347),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1368),
.B(n_1186),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1508),
.Y(n_1560)
);

NAND2x1_ASAP7_75t_L g1561 ( 
.A(n_1393),
.B(n_1093),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1364),
.B(n_1074),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1368),
.B(n_1191),
.Y(n_1563)
);

OAI21xp33_ASAP7_75t_L g1564 ( 
.A1(n_1364),
.A2(n_572),
.B(n_571),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1310),
.B(n_1255),
.Y(n_1565)
);

INVx8_ASAP7_75t_L g1566 ( 
.A(n_1452),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1442),
.B(n_1237),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1290),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1321),
.B(n_1329),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1309),
.B(n_1089),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1486),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1279),
.B(n_1196),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1310),
.B(n_1198),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1437),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1358),
.Y(n_1575)
);

OR2x2_ASAP7_75t_SL g1576 ( 
.A(n_1481),
.B(n_1116),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1358),
.Y(n_1577)
);

INVx8_ASAP7_75t_L g1578 ( 
.A(n_1452),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1310),
.B(n_1304),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1280),
.Y(n_1580)
);

INVxp67_ASAP7_75t_L g1581 ( 
.A(n_1519),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1309),
.B(n_1374),
.Y(n_1582)
);

INVx4_ASAP7_75t_L g1583 ( 
.A(n_1304),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1374),
.B(n_1074),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1279),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1280),
.Y(n_1586)
);

AND2x4_ASAP7_75t_L g1587 ( 
.A(n_1279),
.B(n_1210),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1369),
.B(n_1217),
.Y(n_1588)
);

INVx1_ASAP7_75t_SL g1589 ( 
.A(n_1470),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_1448),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1486),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1284),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1284),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1292),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1516),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1317),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1292),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1317),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1318),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1318),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1305),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1516),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1319),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1305),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1384),
.B(n_1077),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1448),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1516),
.Y(n_1607)
);

NAND2x1p5_ASAP7_75t_L g1608 ( 
.A(n_1304),
.B(n_1275),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1311),
.B(n_1218),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1417),
.A2(n_1229),
.B1(n_1230),
.B2(n_1219),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1348),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1418),
.B(n_1077),
.Y(n_1612)
);

INVx4_ASAP7_75t_L g1613 ( 
.A(n_1311),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1297),
.B(n_1232),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1319),
.Y(n_1615)
);

NAND2x1p5_ASAP7_75t_L g1616 ( 
.A(n_1311),
.B(n_1275),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1316),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1320),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1316),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1519),
.B(n_1152),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1323),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1369),
.B(n_1243),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1323),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1325),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1384),
.B(n_1106),
.Y(n_1625)
);

AO22x2_ASAP7_75t_L g1626 ( 
.A1(n_1417),
.A2(n_1429),
.B1(n_1434),
.B2(n_1356),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1320),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1325),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1337),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1484),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1381),
.B(n_1256),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1322),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1491),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_1487),
.Y(n_1634)
);

AO22x2_ASAP7_75t_L g1635 ( 
.A1(n_1417),
.A2(n_584),
.B1(n_588),
.B2(n_587),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1337),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1348),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1297),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_1487),
.Y(n_1639)
);

INVx4_ASAP7_75t_L g1640 ( 
.A(n_1330),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1389),
.B(n_1106),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1297),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1349),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1389),
.B(n_1400),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1381),
.B(n_1258),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1343),
.B(n_1262),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1349),
.Y(n_1647)
);

NAND2xp33_ASAP7_75t_L g1648 ( 
.A(n_1433),
.B(n_1479),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1372),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1448),
.Y(n_1650)
);

AO22x2_ASAP7_75t_L g1651 ( 
.A1(n_1429),
.A2(n_584),
.B1(n_593),
.B2(n_588),
.Y(n_1651)
);

INVx3_ASAP7_75t_L g1652 ( 
.A(n_1281),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1322),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1343),
.B(n_1295),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1349),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1382),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1382),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1395),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1395),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1314),
.Y(n_1660)
);

INVx5_ASAP7_75t_L g1661 ( 
.A(n_1433),
.Y(n_1661)
);

AO22x2_ASAP7_75t_L g1662 ( 
.A1(n_1429),
.A2(n_1356),
.B1(n_1461),
.B2(n_1400),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1411),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1411),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1415),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1328),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1415),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1295),
.B(n_1118),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1351),
.A2(n_1079),
.B1(n_1072),
.B2(n_1263),
.Y(n_1669)
);

AO22x2_ASAP7_75t_L g1670 ( 
.A1(n_1326),
.A2(n_1445),
.B1(n_1377),
.B2(n_1307),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1430),
.B(n_1265),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1423),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1332),
.B(n_1270),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1287),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1448),
.Y(n_1675)
);

BUFx6f_ASAP7_75t_L g1676 ( 
.A(n_1363),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1423),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1334),
.B(n_1118),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1314),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1425),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1425),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1428),
.Y(n_1682)
);

AO22x2_ASAP7_75t_L g1683 ( 
.A1(n_1377),
.A2(n_593),
.B1(n_605),
.B2(n_595),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1430),
.B(n_1093),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1454),
.B(n_1093),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1428),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1515),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1454),
.B(n_1128),
.Y(n_1688)
);

AO22x2_ASAP7_75t_L g1689 ( 
.A1(n_1281),
.A2(n_595),
.B1(n_615),
.B2(n_605),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1352),
.B(n_1107),
.Y(n_1690)
);

INVx3_ASAP7_75t_L g1691 ( 
.A(n_1281),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1495),
.B(n_1152),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1515),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1517),
.B(n_1095),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1287),
.Y(n_1695)
);

INVx4_ASAP7_75t_L g1696 ( 
.A(n_1330),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1363),
.Y(n_1697)
);

BUFx6f_ASAP7_75t_L g1698 ( 
.A(n_1363),
.Y(n_1698)
);

AO22x2_ASAP7_75t_L g1699 ( 
.A1(n_1283),
.A2(n_615),
.B1(n_617),
.B2(n_616),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1330),
.B(n_1128),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1432),
.B(n_1128),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1432),
.B(n_1129),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1500),
.B(n_1154),
.Y(n_1703)
);

BUFx3_ASAP7_75t_L g1704 ( 
.A(n_1424),
.Y(n_1704)
);

INVx3_ASAP7_75t_L g1705 ( 
.A(n_1283),
.Y(n_1705)
);

INVx5_ASAP7_75t_L g1706 ( 
.A(n_1433),
.Y(n_1706)
);

BUFx4f_ASAP7_75t_L g1707 ( 
.A(n_1372),
.Y(n_1707)
);

A2O1A1Ixp33_ASAP7_75t_L g1708 ( 
.A1(n_1439),
.A2(n_616),
.B(n_625),
.C(n_617),
.Y(n_1708)
);

CKINVDCx20_ASAP7_75t_R g1709 ( 
.A(n_1278),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1439),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1464),
.B(n_1238),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1513),
.B(n_1154),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1447),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1478),
.B(n_1446),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1447),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1472),
.Y(n_1716)
);

CKINVDCx16_ASAP7_75t_R g1717 ( 
.A(n_1386),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1478),
.B(n_1129),
.Y(n_1718)
);

BUFx3_ASAP7_75t_L g1719 ( 
.A(n_1424),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1449),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1328),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1449),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1345),
.B(n_1129),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1483),
.B(n_1266),
.Y(n_1724)
);

INVxp67_ASAP7_75t_L g1725 ( 
.A(n_1472),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1331),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1451),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1331),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1463),
.B(n_1072),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1451),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1333),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1402),
.B(n_1079),
.Y(n_1732)
);

AO22x2_ASAP7_75t_L g1733 ( 
.A1(n_1283),
.A2(n_625),
.B1(n_646),
.B2(n_644),
.Y(n_1733)
);

INVx3_ASAP7_75t_L g1734 ( 
.A(n_1458),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1433),
.B(n_1275),
.Y(n_1735)
);

INVxp67_ASAP7_75t_L g1736 ( 
.A(n_1443),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1477),
.B(n_1288),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_1387),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1453),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1345),
.B(n_1135),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1333),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1453),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1460),
.Y(n_1743)
);

INVx2_ASAP7_75t_SL g1744 ( 
.A(n_1350),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1460),
.Y(n_1745)
);

INVx4_ASAP7_75t_L g1746 ( 
.A(n_1433),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1469),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1474),
.B(n_1135),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1345),
.B(n_1135),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1469),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1342),
.B(n_1137),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1473),
.Y(n_1752)
);

BUFx6f_ASAP7_75t_L g1753 ( 
.A(n_1387),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1291),
.B(n_598),
.Y(n_1754)
);

AO22x2_ASAP7_75t_L g1755 ( 
.A1(n_1335),
.A2(n_1354),
.B1(n_1299),
.B2(n_1301),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1285),
.A2(n_1158),
.B1(n_1159),
.B2(n_1137),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1278),
.Y(n_1757)
);

INVx2_ASAP7_75t_SL g1758 ( 
.A(n_1350),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1336),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_1466),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_1466),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1473),
.Y(n_1762)
);

NAND2x1p5_ASAP7_75t_L g1763 ( 
.A(n_1387),
.B(n_1137),
.Y(n_1763)
);

INVx3_ASAP7_75t_L g1764 ( 
.A(n_1458),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1302),
.B(n_1260),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1336),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1480),
.Y(n_1767)
);

NAND2xp33_ASAP7_75t_L g1768 ( 
.A(n_1524),
.B(n_1479),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1644),
.B(n_1397),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1654),
.B(n_1397),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1644),
.B(n_1397),
.Y(n_1771)
);

NOR2xp67_ASAP7_75t_L g1772 ( 
.A(n_1543),
.B(n_1296),
.Y(n_1772)
);

NOR2xp67_ASAP7_75t_SL g1773 ( 
.A(n_1661),
.B(n_1403),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1532),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1539),
.B(n_1737),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1724),
.B(n_1403),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1590),
.B(n_1440),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_1560),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1581),
.B(n_1315),
.Y(n_1779)
);

INVxp67_ASAP7_75t_L g1780 ( 
.A(n_1527),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1661),
.B(n_1403),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1547),
.B(n_1399),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_1560),
.Y(n_1783)
);

NAND2x1p5_ASAP7_75t_L g1784 ( 
.A(n_1661),
.B(n_1407),
.Y(n_1784)
);

NAND2x1p5_ASAP7_75t_L g1785 ( 
.A(n_1661),
.B(n_1407),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1736),
.B(n_1413),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1711),
.B(n_1660),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1570),
.A2(n_1670),
.B1(n_1527),
.B2(n_1569),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1660),
.B(n_1407),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1596),
.Y(n_1790)
);

NOR2x1p5_ASAP7_75t_L g1791 ( 
.A(n_1704),
.B(n_1440),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1679),
.B(n_1475),
.Y(n_1792)
);

O2A1O1Ixp5_ASAP7_75t_L g1793 ( 
.A1(n_1541),
.A2(n_1353),
.B(n_1468),
.C(n_1462),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_SL g1794 ( 
.A(n_1706),
.B(n_1475),
.Y(n_1794)
);

INVx5_ASAP7_75t_L g1795 ( 
.A(n_1524),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1706),
.B(n_1475),
.Y(n_1796)
);

O2A1O1Ixp5_ASAP7_75t_L g1797 ( 
.A1(n_1573),
.A2(n_1735),
.B(n_1610),
.C(n_1609),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1679),
.B(n_1501),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1646),
.B(n_1501),
.Y(n_1799)
);

AOI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1570),
.A2(n_1467),
.B1(n_1427),
.B2(n_1406),
.Y(n_1800)
);

NAND2x1_ASAP7_75t_L g1801 ( 
.A(n_1524),
.B(n_1479),
.Y(n_1801)
);

INVx2_ASAP7_75t_SL g1802 ( 
.A(n_1568),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1569),
.B(n_1366),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1537),
.B(n_1501),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1596),
.Y(n_1805)
);

INVx8_ASAP7_75t_L g1806 ( 
.A(n_1535),
.Y(n_1806)
);

AND2x6_ASAP7_75t_SL g1807 ( 
.A(n_1620),
.B(n_1388),
.Y(n_1807)
);

INVx1_ASAP7_75t_SL g1808 ( 
.A(n_1716),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1538),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_SL g1810 ( 
.A(n_1706),
.B(n_1479),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1568),
.B(n_1370),
.Y(n_1811)
);

OAI21xp33_ASAP7_75t_L g1812 ( 
.A1(n_1526),
.A2(n_1416),
.B(n_1383),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1542),
.B(n_1344),
.Y(n_1813)
);

OR2x6_ASAP7_75t_L g1814 ( 
.A(n_1535),
.B(n_1350),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1706),
.B(n_1479),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1670),
.A2(n_1503),
.B1(n_1398),
.B2(n_1435),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1552),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1598),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1714),
.B(n_1357),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1598),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1558),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1575),
.B(n_1577),
.Y(n_1822)
);

NAND3xp33_ASAP7_75t_SL g1823 ( 
.A(n_1678),
.B(n_1476),
.C(n_1133),
.Y(n_1823)
);

INVx2_ASAP7_75t_SL g1824 ( 
.A(n_1540),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_SL g1825 ( 
.A1(n_1670),
.A2(n_1123),
.B1(n_1133),
.B2(n_1260),
.Y(n_1825)
);

OAI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1573),
.A2(n_1361),
.B(n_1355),
.Y(n_1826)
);

BUFx3_ASAP7_75t_L g1827 ( 
.A(n_1540),
.Y(n_1827)
);

NOR2x2_ASAP7_75t_L g1828 ( 
.A(n_1683),
.B(n_1350),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1662),
.A2(n_1408),
.B1(n_1294),
.B2(n_1465),
.Y(n_1829)
);

INVxp67_ASAP7_75t_L g1830 ( 
.A(n_1637),
.Y(n_1830)
);

NOR2x2_ASAP7_75t_L g1831 ( 
.A(n_1683),
.B(n_1414),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1580),
.B(n_1511),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1586),
.B(n_1511),
.Y(n_1833)
);

AOI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1551),
.A2(n_1286),
.B1(n_1308),
.B2(n_1414),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1714),
.B(n_1583),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1700),
.Y(n_1836)
);

AND2x4_ASAP7_75t_L g1837 ( 
.A(n_1590),
.B(n_1457),
.Y(n_1837)
);

INVx2_ASAP7_75t_SL g1838 ( 
.A(n_1546),
.Y(n_1838)
);

INVx2_ASAP7_75t_SL g1839 ( 
.A(n_1546),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1592),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1593),
.B(n_1376),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1714),
.B(n_1357),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1583),
.B(n_1357),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1594),
.B(n_1421),
.Y(n_1844)
);

HB1xp67_ASAP7_75t_L g1845 ( 
.A(n_1637),
.Y(n_1845)
);

A2O1A1Ixp33_ASAP7_75t_L g1846 ( 
.A1(n_1597),
.A2(n_1285),
.B(n_1394),
.C(n_1422),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1683),
.A2(n_1414),
.B1(n_1394),
.B2(n_697),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1601),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_SL g1849 ( 
.A(n_1583),
.B(n_1357),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1604),
.B(n_1414),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1668),
.B(n_1357),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1617),
.B(n_1312),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1648),
.A2(n_1391),
.B(n_1357),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1751),
.A2(n_1390),
.B(n_1365),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1619),
.B(n_1441),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1620),
.B(n_1497),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1621),
.B(n_1444),
.Y(n_1857)
);

OAI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1559),
.A2(n_1299),
.B(n_1298),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1623),
.B(n_1367),
.Y(n_1859)
);

NAND2xp33_ASAP7_75t_L g1860 ( 
.A(n_1524),
.B(n_1391),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1599),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1624),
.B(n_1367),
.Y(n_1862)
);

NOR2x1p5_ASAP7_75t_L g1863 ( 
.A(n_1704),
.B(n_1146),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1599),
.Y(n_1864)
);

NOR2xp67_ASAP7_75t_L g1865 ( 
.A(n_1612),
.B(n_1518),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1628),
.B(n_1367),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1662),
.A2(n_697),
.B1(n_712),
.B2(n_576),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1600),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1629),
.B(n_1375),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1636),
.B(n_1375),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1600),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1710),
.B(n_1656),
.Y(n_1872)
);

BUFx8_ASAP7_75t_L g1873 ( 
.A(n_1757),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1557),
.B(n_1457),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1657),
.B(n_1375),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1658),
.B(n_1380),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1659),
.B(n_1380),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1663),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1664),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_1613),
.B(n_1640),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1665),
.B(n_1380),
.Y(n_1881)
);

INVx3_ASAP7_75t_L g1882 ( 
.A(n_1700),
.Y(n_1882)
);

BUFx6f_ASAP7_75t_L g1883 ( 
.A(n_1531),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1667),
.B(n_1480),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1662),
.A2(n_712),
.B1(n_646),
.B2(n_647),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1603),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1672),
.B(n_1482),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1613),
.B(n_1391),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1677),
.B(n_1482),
.Y(n_1889)
);

INVx2_ASAP7_75t_SL g1890 ( 
.A(n_1649),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1626),
.A2(n_1450),
.B1(n_1391),
.B2(n_1341),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1680),
.B(n_1485),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1681),
.B(n_1485),
.Y(n_1893)
);

OAI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1563),
.A2(n_1301),
.B(n_1298),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1603),
.Y(n_1895)
);

NAND2x1p5_ASAP7_75t_L g1896 ( 
.A(n_1531),
.B(n_1613),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1682),
.B(n_1490),
.Y(n_1897)
);

BUFx3_ASAP7_75t_L g1898 ( 
.A(n_1535),
.Y(n_1898)
);

AOI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1562),
.A2(n_1496),
.B1(n_1494),
.B2(n_1476),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1686),
.B(n_1490),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_SL g1901 ( 
.A(n_1640),
.B(n_1391),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_L g1902 ( 
.A1(n_1635),
.A2(n_1651),
.B1(n_1699),
.B2(n_1689),
.Y(n_1902)
);

INVxp67_ASAP7_75t_L g1903 ( 
.A(n_1649),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1574),
.B(n_1324),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1713),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1715),
.Y(n_1906)
);

BUFx3_ASAP7_75t_L g1907 ( 
.A(n_1566),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1687),
.B(n_1498),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1693),
.B(n_1498),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1640),
.B(n_1391),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1648),
.A2(n_1450),
.B(n_1492),
.Y(n_1911)
);

INVx2_ASAP7_75t_SL g1912 ( 
.A(n_1611),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1671),
.B(n_1499),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1671),
.B(n_1582),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1615),
.Y(n_1915)
);

INVx4_ASAP7_75t_L g1916 ( 
.A(n_1524),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1605),
.A2(n_1155),
.B1(n_704),
.B2(n_714),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1729),
.B(n_1589),
.Y(n_1918)
);

A2O1A1Ixp33_ASAP7_75t_L g1919 ( 
.A1(n_1582),
.A2(n_1504),
.B(n_1510),
.C(n_1499),
.Y(n_1919)
);

AOI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1625),
.A2(n_1155),
.B1(n_740),
.B2(n_749),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1630),
.B(n_1324),
.Y(n_1921)
);

BUFx3_ASAP7_75t_L g1922 ( 
.A(n_1566),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1671),
.B(n_1510),
.Y(n_1923)
);

NOR2xp67_ASAP7_75t_L g1924 ( 
.A(n_1612),
.B(n_1504),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1588),
.B(n_1512),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1622),
.B(n_1512),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1633),
.B(n_1386),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1635),
.A2(n_647),
.B1(n_651),
.B2(n_644),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1735),
.A2(n_1450),
.B(n_1505),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1631),
.B(n_1340),
.Y(n_1930)
);

AO22x1_ASAP7_75t_L g1931 ( 
.A1(n_1732),
.A2(n_1260),
.B1(n_579),
.B2(n_582),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1645),
.B(n_1340),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1725),
.B(n_1386),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1585),
.B(n_1360),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1585),
.B(n_1360),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1638),
.B(n_1362),
.Y(n_1936)
);

AOI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1641),
.A2(n_756),
.B1(n_759),
.B2(n_702),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1615),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1720),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1722),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1618),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1642),
.B(n_1362),
.Y(n_1942)
);

INVx2_ASAP7_75t_SL g1943 ( 
.A(n_1707),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1669),
.B(n_1456),
.Y(n_1944)
);

A2O1A1Ixp33_ASAP7_75t_SL g1945 ( 
.A1(n_1652),
.A2(n_1459),
.B(n_1489),
.C(n_1458),
.Y(n_1945)
);

OAI22xp5_ASAP7_75t_SL g1946 ( 
.A1(n_1709),
.A2(n_609),
.B1(n_634),
.B2(n_592),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1727),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1765),
.A2(n_1521),
.B1(n_1378),
.B2(n_1379),
.Y(n_1948)
);

INVx2_ASAP7_75t_SL g1949 ( 
.A(n_1707),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1643),
.B(n_1373),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1531),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1647),
.B(n_1373),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1655),
.B(n_1378),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1692),
.B(n_1703),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1684),
.B(n_1379),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1684),
.B(n_1385),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1684),
.B(n_1385),
.Y(n_1957)
);

NAND2xp33_ASAP7_75t_L g1958 ( 
.A(n_1676),
.B(n_1450),
.Y(n_1958)
);

O2A1O1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1708),
.A2(n_652),
.B(n_656),
.C(n_651),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1685),
.B(n_1392),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1730),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1739),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1685),
.B(n_1392),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1696),
.B(n_1450),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1712),
.B(n_1456),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1606),
.B(n_1426),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1685),
.B(n_1396),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1618),
.Y(n_1968)
);

INVxp67_ASAP7_75t_L g1969 ( 
.A(n_1584),
.Y(n_1969)
);

AOI22xp33_ASAP7_75t_L g1970 ( 
.A1(n_1635),
.A2(n_656),
.B1(n_657),
.B2(n_652),
.Y(n_1970)
);

AOI22xp33_ASAP7_75t_L g1971 ( 
.A1(n_1651),
.A2(n_1689),
.B1(n_1733),
.B2(n_1699),
.Y(n_1971)
);

NAND2xp33_ASAP7_75t_L g1972 ( 
.A(n_1676),
.B(n_1450),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1690),
.B(n_1456),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1742),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1688),
.B(n_1396),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1688),
.B(n_1404),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1564),
.B(n_1459),
.Y(n_1977)
);

AOI22xp33_ASAP7_75t_L g1978 ( 
.A1(n_1651),
.A2(n_658),
.B1(n_660),
.B2(n_657),
.Y(n_1978)
);

AND2x6_ASAP7_75t_L g1979 ( 
.A(n_1836),
.B(n_1676),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_R g1980 ( 
.A(n_1778),
.B(n_1674),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1787),
.B(n_1754),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1774),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1809),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1954),
.B(n_1584),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1803),
.B(n_1688),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1817),
.Y(n_1986)
);

BUFx2_ASAP7_75t_L g1987 ( 
.A(n_1912),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1790),
.Y(n_1988)
);

HB1xp67_ASAP7_75t_L g1989 ( 
.A(n_1845),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1803),
.B(n_1626),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1805),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1818),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1776),
.B(n_1626),
.Y(n_1993)
);

NOR2xp33_ASAP7_75t_L g1994 ( 
.A(n_1780),
.B(n_1674),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1914),
.B(n_1673),
.Y(n_1995)
);

NAND2xp33_ASAP7_75t_SL g1996 ( 
.A(n_1916),
.B(n_1676),
.Y(n_1996)
);

INVx5_ASAP7_75t_L g1997 ( 
.A(n_1795),
.Y(n_1997)
);

AND2x4_ASAP7_75t_L g1998 ( 
.A(n_1898),
.B(n_1606),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1844),
.B(n_1567),
.Y(n_1999)
);

AOI22xp33_ASAP7_75t_L g2000 ( 
.A1(n_1788),
.A2(n_1528),
.B1(n_1765),
.B2(n_1699),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1820),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1799),
.B(n_1567),
.Y(n_2002)
);

BUFx6f_ASAP7_75t_L g2003 ( 
.A(n_1883),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1861),
.Y(n_2004)
);

NAND3xp33_ASAP7_75t_SL g2005 ( 
.A(n_1816),
.B(n_1800),
.C(n_1856),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_1898),
.B(n_1650),
.Y(n_2006)
);

AND2x6_ASAP7_75t_L g2007 ( 
.A(n_1836),
.B(n_1697),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_1783),
.Y(n_2008)
);

INVx2_ASAP7_75t_SL g2009 ( 
.A(n_1827),
.Y(n_2009)
);

BUFx2_ASAP7_75t_L g2010 ( 
.A(n_1845),
.Y(n_2010)
);

AOI22xp33_ASAP7_75t_SL g2011 ( 
.A1(n_1944),
.A2(n_1528),
.B1(n_1755),
.B2(n_1695),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1782),
.B(n_1760),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1864),
.Y(n_2013)
);

BUFx5_ASAP7_75t_L g2014 ( 
.A(n_1905),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1821),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1868),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1840),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_1873),
.Y(n_2018)
);

BUFx3_ASAP7_75t_L g2019 ( 
.A(n_1806),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1871),
.Y(n_2020)
);

AND2x4_ASAP7_75t_L g2021 ( 
.A(n_1907),
.B(n_1650),
.Y(n_2021)
);

INVx2_ASAP7_75t_SL g2022 ( 
.A(n_1827),
.Y(n_2022)
);

BUFx6f_ASAP7_75t_L g2023 ( 
.A(n_1883),
.Y(n_2023)
);

INVxp67_ASAP7_75t_L g2024 ( 
.A(n_1890),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1848),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1770),
.B(n_1769),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1878),
.Y(n_2027)
);

AND2x4_ASAP7_75t_L g2028 ( 
.A(n_1907),
.B(n_1675),
.Y(n_2028)
);

AND2x6_ASAP7_75t_L g2029 ( 
.A(n_1882),
.B(n_1697),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1879),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1906),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1918),
.B(n_1760),
.Y(n_2032)
);

BUFx3_ASAP7_75t_L g2033 ( 
.A(n_1806),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1939),
.Y(n_2034)
);

AND2x6_ASAP7_75t_L g2035 ( 
.A(n_1882),
.B(n_1697),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1918),
.B(n_1761),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1813),
.B(n_1567),
.Y(n_2037)
);

BUFx12f_ASAP7_75t_L g2038 ( 
.A(n_1873),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1940),
.Y(n_2039)
);

NOR2xp33_ASAP7_75t_L g2040 ( 
.A(n_1775),
.B(n_1695),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1947),
.Y(n_2041)
);

OR2x2_ASAP7_75t_SL g2042 ( 
.A(n_1823),
.B(n_1717),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1922),
.B(n_1675),
.Y(n_2043)
);

BUFx6f_ASAP7_75t_L g2044 ( 
.A(n_1883),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1886),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1961),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1962),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1895),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_R g2049 ( 
.A(n_1943),
.B(n_1761),
.Y(n_2049)
);

AND2x4_ASAP7_75t_L g2050 ( 
.A(n_1922),
.B(n_1744),
.Y(n_2050)
);

INVxp67_ASAP7_75t_L g2051 ( 
.A(n_1808),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1874),
.B(n_1744),
.Y(n_2052)
);

CKINVDCx9p33_ASAP7_75t_R g2053 ( 
.A(n_1927),
.Y(n_2053)
);

NAND2x1p5_ASAP7_75t_L g2054 ( 
.A(n_1795),
.B(n_1531),
.Y(n_2054)
);

BUFx3_ASAP7_75t_L g2055 ( 
.A(n_1806),
.Y(n_2055)
);

BUFx4f_ASAP7_75t_L g2056 ( 
.A(n_1837),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1974),
.Y(n_2057)
);

INVx1_ASAP7_75t_SL g2058 ( 
.A(n_1802),
.Y(n_2058)
);

AOI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_1856),
.A2(n_1554),
.B1(n_1534),
.B2(n_1694),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1841),
.B(n_1748),
.Y(n_2060)
);

HB1xp67_ASAP7_75t_L g2061 ( 
.A(n_1830),
.Y(n_2061)
);

INVx3_ASAP7_75t_L g2062 ( 
.A(n_1916),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_1769),
.B(n_1697),
.Y(n_2063)
);

BUFx10_ASAP7_75t_L g2064 ( 
.A(n_1927),
.Y(n_2064)
);

INVx3_ASAP7_75t_L g2065 ( 
.A(n_1896),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1822),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1872),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1855),
.B(n_1525),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1915),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1938),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1965),
.B(n_1758),
.Y(n_2071)
);

BUFx2_ASAP7_75t_L g2072 ( 
.A(n_1903),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1941),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1857),
.B(n_1525),
.Y(n_2074)
);

NOR2x1_ASAP7_75t_R g2075 ( 
.A(n_1777),
.B(n_1719),
.Y(n_2075)
);

AND2x4_ASAP7_75t_L g2076 ( 
.A(n_1837),
.B(n_1758),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1968),
.Y(n_2077)
);

BUFx10_ASAP7_75t_L g2078 ( 
.A(n_1786),
.Y(n_2078)
);

BUFx6f_ASAP7_75t_L g2079 ( 
.A(n_1883),
.Y(n_2079)
);

CKINVDCx5p33_ASAP7_75t_R g2080 ( 
.A(n_1807),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1969),
.B(n_1572),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1921),
.B(n_1528),
.Y(n_2082)
);

BUFx6f_ASAP7_75t_L g2083 ( 
.A(n_1951),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1884),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1887),
.Y(n_2085)
);

AO21x1_ASAP7_75t_L g2086 ( 
.A1(n_1771),
.A2(n_1554),
.B(n_1609),
.Y(n_2086)
);

INVxp33_ASAP7_75t_L g2087 ( 
.A(n_1779),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_SL g2088 ( 
.A(n_1771),
.B(n_1698),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_R g2089 ( 
.A(n_1949),
.B(n_1709),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1936),
.Y(n_2090)
);

AND2x6_ASAP7_75t_L g2091 ( 
.A(n_1951),
.B(n_1698),
.Y(n_2091)
);

BUFx3_ASAP7_75t_L g2092 ( 
.A(n_1777),
.Y(n_2092)
);

AND2x2_ASAP7_75t_SL g2093 ( 
.A(n_1885),
.B(n_1698),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1942),
.Y(n_2094)
);

INVx3_ASAP7_75t_L g2095 ( 
.A(n_1896),
.Y(n_2095)
);

INVx3_ASAP7_75t_L g2096 ( 
.A(n_1795),
.Y(n_2096)
);

AND2x4_ASAP7_75t_L g2097 ( 
.A(n_1791),
.B(n_1814),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1859),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1832),
.B(n_1572),
.Y(n_2099)
);

INVx2_ASAP7_75t_SL g2100 ( 
.A(n_1824),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_1814),
.B(n_1719),
.Y(n_2101)
);

BUFx3_ASAP7_75t_L g2102 ( 
.A(n_1838),
.Y(n_2102)
);

INVx4_ASAP7_75t_L g2103 ( 
.A(n_1795),
.Y(n_2103)
);

NOR3xp33_ASAP7_75t_SL g2104 ( 
.A(n_1812),
.B(n_1786),
.C(n_1944),
.Y(n_2104)
);

INVx3_ASAP7_75t_L g2105 ( 
.A(n_1951),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1889),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_1921),
.B(n_1572),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_R g2108 ( 
.A(n_1973),
.B(n_1566),
.Y(n_2108)
);

INVx2_ASAP7_75t_SL g2109 ( 
.A(n_1839),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1862),
.Y(n_2110)
);

INVxp67_ASAP7_75t_SL g2111 ( 
.A(n_1768),
.Y(n_2111)
);

NOR3xp33_ASAP7_75t_SL g2112 ( 
.A(n_1779),
.B(n_1708),
.C(n_589),
.Y(n_2112)
);

NOR3xp33_ASAP7_75t_SL g2113 ( 
.A(n_1946),
.B(n_590),
.C(n_577),
.Y(n_2113)
);

NOR2xp33_ASAP7_75t_L g2114 ( 
.A(n_1798),
.B(n_1576),
.Y(n_2114)
);

OR2x2_ASAP7_75t_L g2115 ( 
.A(n_1850),
.B(n_1530),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_1814),
.B(n_1587),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1892),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1833),
.B(n_1804),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_1966),
.B(n_1587),
.Y(n_2119)
);

BUFx3_ASAP7_75t_L g2120 ( 
.A(n_1966),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1865),
.B(n_1587),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1811),
.B(n_1614),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1893),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1811),
.B(n_1614),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1897),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1925),
.B(n_1614),
.Y(n_2126)
);

NOR3xp33_ASAP7_75t_SL g2127 ( 
.A(n_1904),
.B(n_597),
.C(n_596),
.Y(n_2127)
);

AND2x4_ASAP7_75t_L g2128 ( 
.A(n_1863),
.B(n_1772),
.Y(n_2128)
);

NOR3xp33_ASAP7_75t_SL g2129 ( 
.A(n_1904),
.B(n_602),
.C(n_601),
.Y(n_2129)
);

BUFx4f_ASAP7_75t_L g2130 ( 
.A(n_1951),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1926),
.B(n_1755),
.Y(n_2131)
);

NAND2x1p5_ASAP7_75t_L g2132 ( 
.A(n_1773),
.B(n_1746),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1924),
.B(n_1755),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1950),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_R g2135 ( 
.A(n_1933),
.B(n_1578),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1930),
.B(n_1743),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1900),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1932),
.B(n_1745),
.Y(n_2138)
);

INVx2_ASAP7_75t_SL g2139 ( 
.A(n_1933),
.Y(n_2139)
);

NOR2xp33_ASAP7_75t_L g2140 ( 
.A(n_1852),
.B(n_1571),
.Y(n_2140)
);

NOR2xp33_ASAP7_75t_L g2141 ( 
.A(n_1899),
.B(n_1571),
.Y(n_2141)
);

BUFx2_ASAP7_75t_L g2142 ( 
.A(n_1828),
.Y(n_2142)
);

NOR2xp33_ASAP7_75t_L g2143 ( 
.A(n_1789),
.B(n_1792),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1908),
.Y(n_2144)
);

AND2x4_ASAP7_75t_L g2145 ( 
.A(n_1835),
.B(n_1523),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1866),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1909),
.Y(n_2147)
);

CKINVDCx11_ASAP7_75t_R g2148 ( 
.A(n_1931),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1913),
.B(n_1747),
.Y(n_2149)
);

BUFx3_ASAP7_75t_L g2150 ( 
.A(n_1784),
.Y(n_2150)
);

BUFx2_ASAP7_75t_L g2151 ( 
.A(n_1831),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1923),
.B(n_1750),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1952),
.Y(n_2153)
);

INVx3_ASAP7_75t_L g2154 ( 
.A(n_1801),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1834),
.B(n_1752),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1847),
.B(n_1928),
.Y(n_2156)
);

BUFx3_ASAP7_75t_L g2157 ( 
.A(n_1784),
.Y(n_2157)
);

AND2x4_ASAP7_75t_L g2158 ( 
.A(n_1835),
.B(n_1523),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1847),
.B(n_1762),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1953),
.Y(n_2160)
);

BUFx4f_ASAP7_75t_SL g2161 ( 
.A(n_1851),
.Y(n_2161)
);

NAND2xp33_ASAP7_75t_R g2162 ( 
.A(n_1911),
.B(n_1652),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_1917),
.Y(n_2163)
);

NAND2x1_ASAP7_75t_L g2164 ( 
.A(n_1934),
.B(n_1746),
.Y(n_2164)
);

INVx1_ASAP7_75t_SL g2165 ( 
.A(n_1955),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1869),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1870),
.Y(n_2167)
);

INVx3_ASAP7_75t_L g2168 ( 
.A(n_1785),
.Y(n_2168)
);

AND2x4_ASAP7_75t_L g2169 ( 
.A(n_1956),
.B(n_1523),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1978),
.B(n_1767),
.Y(n_2170)
);

NOR3xp33_ASAP7_75t_SL g2171 ( 
.A(n_1959),
.B(n_607),
.C(n_606),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1957),
.Y(n_2172)
);

BUFx6f_ASAP7_75t_L g2173 ( 
.A(n_1785),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1960),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1875),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_1928),
.B(n_1970),
.Y(n_2176)
);

AOI22xp5_ASAP7_75t_SL g2177 ( 
.A1(n_1825),
.A2(n_610),
.B1(n_613),
.B2(n_608),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1876),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1978),
.B(n_1970),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1826),
.B(n_1718),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1877),
.Y(n_2181)
);

AND2x4_ASAP7_75t_L g2182 ( 
.A(n_1963),
.B(n_1571),
.Y(n_2182)
);

INVx4_ASAP7_75t_L g2183 ( 
.A(n_1958),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1881),
.Y(n_2184)
);

NOR2xp33_ASAP7_75t_R g2185 ( 
.A(n_1972),
.B(n_1578),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1935),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_1967),
.Y(n_2187)
);

AND2x4_ASAP7_75t_L g2188 ( 
.A(n_1975),
.B(n_1571),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1976),
.Y(n_2189)
);

HB1xp67_ASAP7_75t_L g2190 ( 
.A(n_1819),
.Y(n_2190)
);

AND2x4_ASAP7_75t_L g2191 ( 
.A(n_1819),
.B(n_1591),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1885),
.B(n_1718),
.Y(n_2192)
);

CKINVDCx5p33_ASAP7_75t_R g2193 ( 
.A(n_1920),
.Y(n_2193)
);

OAI21xp5_ASAP7_75t_L g2194 ( 
.A1(n_1797),
.A2(n_1579),
.B(n_1718),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1948),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1919),
.Y(n_2196)
);

NOR2xp33_ASAP7_75t_R g2197 ( 
.A(n_1860),
.B(n_1578),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_L g2198 ( 
.A(n_1937),
.B(n_1591),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1867),
.B(n_1533),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1977),
.Y(n_2200)
);

INVx3_ASAP7_75t_L g2201 ( 
.A(n_1880),
.Y(n_2201)
);

O2A1O1Ixp33_ASAP7_75t_L g2202 ( 
.A1(n_1846),
.A2(n_867),
.B(n_868),
.C(n_866),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1977),
.Y(n_2203)
);

BUFx6f_ASAP7_75t_L g2204 ( 
.A(n_1810),
.Y(n_2204)
);

NOR2xp33_ASAP7_75t_SL g2205 ( 
.A(n_1829),
.B(n_1591),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_1867),
.B(n_1502),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1858),
.Y(n_2207)
);

NAND2xp33_ASAP7_75t_R g2208 ( 
.A(n_1854),
.B(n_1652),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1902),
.B(n_1533),
.Y(n_2209)
);

AND2x4_ASAP7_75t_L g2210 ( 
.A(n_1842),
.B(n_1591),
.Y(n_2210)
);

AOI21xp5_ASAP7_75t_L g2211 ( 
.A1(n_2111),
.A2(n_1853),
.B(n_1880),
.Y(n_2211)
);

BUFx6f_ASAP7_75t_L g2212 ( 
.A(n_2130),
.Y(n_2212)
);

OAI21x1_ASAP7_75t_L g2213 ( 
.A1(n_2194),
.A2(n_1891),
.B(n_1894),
.Y(n_2213)
);

A2O1A1Ixp33_ASAP7_75t_L g2214 ( 
.A1(n_2005),
.A2(n_1793),
.B(n_1902),
.C(n_1971),
.Y(n_2214)
);

OAI22xp5_ASAP7_75t_L g2215 ( 
.A1(n_2093),
.A2(n_2179),
.B1(n_2176),
.B2(n_2156),
.Y(n_2215)
);

OAI21x1_ASAP7_75t_L g2216 ( 
.A1(n_2202),
.A2(n_1842),
.B(n_1843),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2084),
.B(n_1971),
.Y(n_2217)
);

OAI21x1_ASAP7_75t_L g2218 ( 
.A1(n_2202),
.A2(n_1964),
.B(n_1849),
.Y(n_2218)
);

AOI21xp5_ASAP7_75t_L g2219 ( 
.A1(n_2111),
.A2(n_1849),
.B(n_1843),
.Y(n_2219)
);

AO31x2_ASAP7_75t_L g2220 ( 
.A1(n_2086),
.A2(n_1929),
.A3(n_1536),
.B(n_1548),
.Y(n_2220)
);

NOR2xp67_ASAP7_75t_R g2221 ( 
.A(n_1997),
.B(n_1698),
.Y(n_2221)
);

INVx4_ASAP7_75t_L g2222 ( 
.A(n_1997),
.Y(n_2222)
);

BUFx6f_ASAP7_75t_L g2223 ( 
.A(n_2130),
.Y(n_2223)
);

OAI21x1_ASAP7_75t_L g2224 ( 
.A1(n_2201),
.A2(n_1888),
.B(n_1901),
.Y(n_2224)
);

OAI21xp5_ASAP7_75t_L g2225 ( 
.A1(n_2005),
.A2(n_1794),
.B(n_1781),
.Y(n_2225)
);

AOI21xp5_ASAP7_75t_SL g2226 ( 
.A1(n_2183),
.A2(n_1753),
.B(n_1738),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2085),
.B(n_1689),
.Y(n_2227)
);

AOI21xp5_ASAP7_75t_L g2228 ( 
.A1(n_2060),
.A2(n_1901),
.B(n_1888),
.Y(n_2228)
);

OAI21x1_ASAP7_75t_L g2229 ( 
.A1(n_2201),
.A2(n_2164),
.B(n_2088),
.Y(n_2229)
);

OAI21x1_ASAP7_75t_L g2230 ( 
.A1(n_2063),
.A2(n_2088),
.B(n_2196),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2106),
.B(n_1733),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1982),
.Y(n_2232)
);

OAI21xp5_ASAP7_75t_L g2233 ( 
.A1(n_2026),
.A2(n_1794),
.B(n_1781),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2117),
.B(n_1733),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2123),
.B(n_1796),
.Y(n_2235)
);

AO31x2_ASAP7_75t_L g2236 ( 
.A1(n_2207),
.A2(n_1536),
.A3(n_1548),
.B(n_1522),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2125),
.B(n_1796),
.Y(n_2237)
);

AO21x2_ASAP7_75t_L g2238 ( 
.A1(n_2026),
.A2(n_1945),
.B(n_1810),
.Y(n_2238)
);

OAI21x1_ASAP7_75t_L g2239 ( 
.A1(n_2063),
.A2(n_1910),
.B(n_1964),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2137),
.B(n_1544),
.Y(n_2240)
);

AOI21x1_ASAP7_75t_SL g2241 ( 
.A1(n_1990),
.A2(n_1740),
.B(n_1723),
.Y(n_2241)
);

OAI21x1_ASAP7_75t_L g2242 ( 
.A1(n_2180),
.A2(n_1910),
.B(n_1549),
.Y(n_2242)
);

AOI21xp5_ASAP7_75t_L g2243 ( 
.A1(n_1995),
.A2(n_1579),
.B(n_1815),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1983),
.Y(n_2244)
);

AOI21x1_ASAP7_75t_L g2245 ( 
.A1(n_1993),
.A2(n_1815),
.B(n_1549),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2144),
.B(n_1544),
.Y(n_2246)
);

BUFx6f_ASAP7_75t_L g2247 ( 
.A(n_2092),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_1980),
.Y(n_2248)
);

OAI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_2093),
.A2(n_2066),
.B1(n_2067),
.B2(n_2000),
.Y(n_2249)
);

AOI21xp5_ASAP7_75t_L g2250 ( 
.A1(n_2037),
.A2(n_1746),
.B(n_1565),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2147),
.B(n_1544),
.Y(n_2251)
);

BUFx3_ASAP7_75t_L g2252 ( 
.A(n_1987),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2118),
.B(n_1545),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_1984),
.B(n_1701),
.Y(n_2254)
);

OAI21xp5_ASAP7_75t_L g2255 ( 
.A1(n_2195),
.A2(n_1945),
.B(n_1756),
.Y(n_2255)
);

OAI21x1_ASAP7_75t_L g2256 ( 
.A1(n_2154),
.A2(n_1522),
.B(n_1691),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2143),
.B(n_1545),
.Y(n_2257)
);

AOI21xp5_ASAP7_75t_L g2258 ( 
.A1(n_2205),
.A2(n_1565),
.B(n_1696),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2143),
.B(n_1545),
.Y(n_2259)
);

OAI21xp5_ASAP7_75t_L g2260 ( 
.A1(n_2104),
.A2(n_1705),
.B(n_1691),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_L g2261 ( 
.A(n_2087),
.B(n_1313),
.Y(n_2261)
);

AOI21xp5_ASAP7_75t_L g2262 ( 
.A1(n_1999),
.A2(n_1696),
.B(n_1753),
.Y(n_2262)
);

AOI21xp5_ASAP7_75t_L g2263 ( 
.A1(n_2002),
.A2(n_1753),
.B(n_1738),
.Y(n_2263)
);

AOI21x1_ASAP7_75t_L g2264 ( 
.A1(n_2200),
.A2(n_1561),
.B(n_1723),
.Y(n_2264)
);

AO31x2_ASAP7_75t_L g2265 ( 
.A1(n_2203),
.A2(n_1632),
.A3(n_1653),
.B(n_1627),
.Y(n_2265)
);

AOI21xp5_ASAP7_75t_L g2266 ( 
.A1(n_1996),
.A2(n_1753),
.B(n_1738),
.Y(n_2266)
);

OAI21x1_ASAP7_75t_L g2267 ( 
.A1(n_2154),
.A2(n_2110),
.B(n_2098),
.Y(n_2267)
);

OAI21x1_ASAP7_75t_L g2268 ( 
.A1(n_2098),
.A2(n_1705),
.B(n_1691),
.Y(n_2268)
);

AOI21xp5_ASAP7_75t_L g2269 ( 
.A1(n_1996),
.A2(n_1738),
.B(n_1616),
.Y(n_2269)
);

OAI21x1_ASAP7_75t_L g2270 ( 
.A1(n_2110),
.A2(n_1705),
.B(n_1763),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2107),
.B(n_1701),
.Y(n_2271)
);

A2O1A1Ixp33_ASAP7_75t_L g2272 ( 
.A1(n_2104),
.A2(n_2114),
.B(n_2141),
.C(n_2112),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1986),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_1981),
.B(n_1701),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_1985),
.B(n_2122),
.Y(n_2275)
);

BUFx6f_ASAP7_75t_L g2276 ( 
.A(n_2092),
.Y(n_2276)
);

OAI21x1_ASAP7_75t_L g2277 ( 
.A1(n_2146),
.A2(n_1763),
.B(n_1602),
.Y(n_2277)
);

AOI21x1_ASAP7_75t_SL g2278 ( 
.A1(n_2128),
.A2(n_1740),
.B(n_1723),
.Y(n_2278)
);

OAI21xp5_ASAP7_75t_L g2279 ( 
.A1(n_2131),
.A2(n_1632),
.B(n_1627),
.Y(n_2279)
);

NAND2x1_ASAP7_75t_L g2280 ( 
.A(n_2183),
.B(n_1553),
.Y(n_2280)
);

AOI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_2136),
.A2(n_1616),
.B(n_1608),
.Y(n_2281)
);

AND2x4_ASAP7_75t_L g2282 ( 
.A(n_2097),
.B(n_1634),
.Y(n_2282)
);

OAI22x1_ASAP7_75t_L g2283 ( 
.A1(n_2059),
.A2(n_660),
.B1(n_670),
.B2(n_658),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2124),
.B(n_1702),
.Y(n_2284)
);

NAND2x1p5_ASAP7_75t_L g2285 ( 
.A(n_1997),
.B(n_1553),
.Y(n_2285)
);

OAI21x1_ASAP7_75t_L g2286 ( 
.A1(n_2146),
.A2(n_2132),
.B(n_2168),
.Y(n_2286)
);

INVx3_ASAP7_75t_L g2287 ( 
.A(n_2103),
.Y(n_2287)
);

AO21x1_ASAP7_75t_L g2288 ( 
.A1(n_2155),
.A2(n_2133),
.B(n_2114),
.Y(n_2288)
);

INVx4_ASAP7_75t_L g2289 ( 
.A(n_1997),
.Y(n_2289)
);

OR2x6_ASAP7_75t_L g2290 ( 
.A(n_2132),
.B(n_1740),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2165),
.B(n_1702),
.Y(n_2291)
);

AOI21xp5_ASAP7_75t_L g2292 ( 
.A1(n_2138),
.A2(n_1608),
.B(n_1529),
.Y(n_2292)
);

AOI21xp5_ASAP7_75t_L g2293 ( 
.A1(n_2126),
.A2(n_1529),
.B(n_1749),
.Y(n_2293)
);

NOR2x1_ASAP7_75t_L g2294 ( 
.A(n_1994),
.B(n_1749),
.Y(n_2294)
);

INVx3_ASAP7_75t_L g2295 ( 
.A(n_2103),
.Y(n_2295)
);

OA21x2_ASAP7_75t_L g2296 ( 
.A1(n_2190),
.A2(n_873),
.B(n_872),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_SL g2297 ( 
.A(n_2163),
.B(n_1634),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_1980),
.Y(n_2298)
);

NAND2x1p5_ASAP7_75t_L g2299 ( 
.A(n_2062),
.B(n_2150),
.Y(n_2299)
);

OAI22x1_ASAP7_75t_L g2300 ( 
.A1(n_2151),
.A2(n_674),
.B1(n_675),
.B2(n_670),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_L g2301 ( 
.A(n_2087),
.B(n_1702),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2153),
.B(n_1653),
.Y(n_2302)
);

A2O1A1Ixp33_ASAP7_75t_L g2303 ( 
.A1(n_2141),
.A2(n_1749),
.B(n_1639),
.C(n_1634),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2015),
.Y(n_2304)
);

BUFx6f_ASAP7_75t_L g2305 ( 
.A(n_2056),
.Y(n_2305)
);

A2O1A1Ixp33_ASAP7_75t_L g2306 ( 
.A1(n_2112),
.A2(n_1639),
.B(n_1634),
.C(n_1533),
.Y(n_2306)
);

BUFx2_ASAP7_75t_L g2307 ( 
.A(n_2051),
.Y(n_2307)
);

NAND2x1p5_ASAP7_75t_L g2308 ( 
.A(n_2062),
.B(n_1639),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_2008),
.Y(n_2309)
);

AO31x2_ASAP7_75t_L g2310 ( 
.A1(n_2159),
.A2(n_1721),
.A3(n_1726),
.B(n_1666),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2160),
.B(n_1666),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_2032),
.B(n_708),
.Y(n_2312)
);

BUFx3_ASAP7_75t_L g2313 ( 
.A(n_2010),
.Y(n_2313)
);

BUFx6f_ASAP7_75t_L g2314 ( 
.A(n_2056),
.Y(n_2314)
);

AOI21xp5_ASAP7_75t_L g2315 ( 
.A1(n_2068),
.A2(n_1700),
.B(n_1639),
.Y(n_2315)
);

A2O1A1Ixp33_ASAP7_75t_L g2316 ( 
.A1(n_2177),
.A2(n_874),
.B(n_1555),
.C(n_1550),
.Y(n_2316)
);

BUFx3_ASAP7_75t_L g2317 ( 
.A(n_2072),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2166),
.B(n_1721),
.Y(n_2318)
);

OA22x2_ASAP7_75t_L g2319 ( 
.A1(n_2193),
.A2(n_675),
.B1(n_679),
.B2(n_674),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2013),
.Y(n_2320)
);

AOI21xp5_ASAP7_75t_L g2321 ( 
.A1(n_2074),
.A2(n_1602),
.B(n_1595),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2090),
.B(n_1726),
.Y(n_2322)
);

INVx1_ASAP7_75t_SL g2323 ( 
.A(n_1989),
.Y(n_2323)
);

AO31x2_ASAP7_75t_L g2324 ( 
.A1(n_2192),
.A2(n_1731),
.A3(n_1741),
.B(n_1728),
.Y(n_2324)
);

AOI21xp5_ASAP7_75t_L g2325 ( 
.A1(n_2198),
.A2(n_1602),
.B(n_1595),
.Y(n_2325)
);

OAI21xp5_ASAP7_75t_L g2326 ( 
.A1(n_2199),
.A2(n_1731),
.B(n_1728),
.Y(n_2326)
);

OAI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_2000),
.A2(n_1759),
.B1(n_1766),
.B2(n_1741),
.Y(n_2327)
);

OAI21x1_ASAP7_75t_L g2328 ( 
.A1(n_2168),
.A2(n_1607),
.B(n_1595),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2094),
.B(n_1759),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2134),
.B(n_2036),
.Y(n_2330)
);

AOI21xp5_ASAP7_75t_L g2331 ( 
.A1(n_2198),
.A2(n_1607),
.B(n_1766),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2172),
.B(n_1550),
.Y(n_2332)
);

NOR2x1_ASAP7_75t_SL g2333 ( 
.A(n_2173),
.B(n_2150),
.Y(n_2333)
);

AND2x4_ASAP7_75t_L g2334 ( 
.A(n_2097),
.B(n_1550),
.Y(n_2334)
);

OAI21xp5_ASAP7_75t_L g2335 ( 
.A1(n_2011),
.A2(n_1405),
.B(n_1404),
.Y(n_2335)
);

AOI21xp5_ASAP7_75t_L g2336 ( 
.A1(n_2149),
.A2(n_1607),
.B(n_1734),
.Y(n_2336)
);

AOI21x1_ASAP7_75t_L g2337 ( 
.A1(n_2190),
.A2(n_1409),
.B(n_1405),
.Y(n_2337)
);

AOI21x1_ASAP7_75t_L g2338 ( 
.A1(n_2170),
.A2(n_2121),
.B(n_2209),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2013),
.Y(n_2339)
);

NAND2xp33_ASAP7_75t_L g2340 ( 
.A(n_2185),
.B(n_1734),
.Y(n_2340)
);

AOI21xp33_ASAP7_75t_L g2341 ( 
.A1(n_2208),
.A2(n_1556),
.B(n_1555),
.Y(n_2341)
);

OAI21x1_ASAP7_75t_L g2342 ( 
.A1(n_2096),
.A2(n_1764),
.B(n_1410),
.Y(n_2342)
);

OAI22x1_ASAP7_75t_L g2343 ( 
.A1(n_2142),
.A2(n_681),
.B1(n_682),
.B2(n_679),
.Y(n_2343)
);

AND2x4_ASAP7_75t_L g2344 ( 
.A(n_1998),
.B(n_1555),
.Y(n_2344)
);

OAI21x1_ASAP7_75t_L g2345 ( 
.A1(n_2096),
.A2(n_2054),
.B(n_2065),
.Y(n_2345)
);

A2O1A1Ixp33_ASAP7_75t_L g2346 ( 
.A1(n_2171),
.A2(n_2040),
.B(n_2140),
.C(n_2129),
.Y(n_2346)
);

AND3x4_ASAP7_75t_L g2347 ( 
.A(n_2128),
.B(n_1556),
.C(n_713),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2167),
.B(n_1764),
.Y(n_2348)
);

AOI21xp5_ASAP7_75t_L g2349 ( 
.A1(n_2152),
.A2(n_2178),
.B(n_2175),
.Y(n_2349)
);

BUFx6f_ASAP7_75t_L g2350 ( 
.A(n_2019),
.Y(n_2350)
);

BUFx3_ASAP7_75t_L g2351 ( 
.A(n_2102),
.Y(n_2351)
);

OAI21x1_ASAP7_75t_L g2352 ( 
.A1(n_2054),
.A2(n_1410),
.B(n_1409),
.Y(n_2352)
);

AOI21xp5_ASAP7_75t_L g2353 ( 
.A1(n_2181),
.A2(n_1556),
.B(n_1489),
.Y(n_2353)
);

AO31x2_ASAP7_75t_L g2354 ( 
.A1(n_2184),
.A2(n_1420),
.A3(n_1438),
.B(n_1412),
.Y(n_2354)
);

OAI21xp5_ASAP7_75t_L g2355 ( 
.A1(n_2011),
.A2(n_1420),
.B(n_1412),
.Y(n_2355)
);

HB1xp67_ASAP7_75t_L g2356 ( 
.A(n_2051),
.Y(n_2356)
);

OAI21x1_ASAP7_75t_L g2357 ( 
.A1(n_2065),
.A2(n_1455),
.B(n_1438),
.Y(n_2357)
);

OAI21x1_ASAP7_75t_L g2358 ( 
.A1(n_2095),
.A2(n_1471),
.B(n_1455),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2082),
.B(n_708),
.Y(n_2359)
);

OAI22xp5_ASAP7_75t_L g2360 ( 
.A1(n_2115),
.A2(n_682),
.B1(n_683),
.B2(n_681),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2174),
.B(n_1471),
.Y(n_2361)
);

INVx4_ASAP7_75t_L g2362 ( 
.A(n_2091),
.Y(n_2362)
);

CKINVDCx8_ASAP7_75t_R g2363 ( 
.A(n_2018),
.Y(n_2363)
);

AOI21xp5_ASAP7_75t_L g2364 ( 
.A1(n_2099),
.A2(n_1489),
.B(n_1459),
.Y(n_2364)
);

AOI21xp5_ASAP7_75t_L g2365 ( 
.A1(n_2186),
.A2(n_2158),
.B(n_2145),
.Y(n_2365)
);

AOI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2145),
.A2(n_1493),
.B(n_1488),
.Y(n_2366)
);

OAI21xp5_ASAP7_75t_L g2367 ( 
.A1(n_2171),
.A2(n_1493),
.B(n_1488),
.Y(n_2367)
);

NOR2xp67_ASAP7_75t_L g2368 ( 
.A(n_2024),
.B(n_1506),
.Y(n_2368)
);

NAND2x1_ASAP7_75t_L g2369 ( 
.A(n_2091),
.B(n_1506),
.Y(n_2369)
);

AOI21xp5_ASAP7_75t_L g2370 ( 
.A1(n_2158),
.A2(n_1509),
.B(n_1507),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2187),
.B(n_1507),
.Y(n_2371)
);

AOI21x1_ASAP7_75t_L g2372 ( 
.A1(n_2191),
.A2(n_1509),
.B(n_1011),
.Y(n_2372)
);

OAI22xp5_ASAP7_75t_L g2373 ( 
.A1(n_2040),
.A2(n_692),
.B1(n_694),
.B2(n_683),
.Y(n_2373)
);

BUFx6f_ASAP7_75t_L g2374 ( 
.A(n_2019),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2077),
.Y(n_2375)
);

OAI21xp5_ASAP7_75t_L g2376 ( 
.A1(n_2140),
.A2(n_1011),
.B(n_1010),
.Y(n_2376)
);

AOI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_2189),
.A2(n_1514),
.B(n_1212),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_1994),
.B(n_620),
.Y(n_2378)
);

BUFx2_ASAP7_75t_L g2379 ( 
.A(n_2089),
.Y(n_2379)
);

BUFx12f_ASAP7_75t_L g2380 ( 
.A(n_2038),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2012),
.B(n_708),
.Y(n_2381)
);

HAxp5_ASAP7_75t_L g2382 ( 
.A(n_2078),
.B(n_678),
.CON(n_2382),
.SN(n_2382)
);

OAI21x1_ASAP7_75t_L g2383 ( 
.A1(n_2095),
.A2(n_1159),
.B(n_1158),
.Y(n_2383)
);

AND2x6_ASAP7_75t_L g2384 ( 
.A(n_2191),
.B(n_692),
.Y(n_2384)
);

AOI21xp5_ASAP7_75t_L g2385 ( 
.A1(n_2162),
.A2(n_1514),
.B(n_1212),
.Y(n_2385)
);

AO31x2_ASAP7_75t_L g2386 ( 
.A1(n_2077),
.A2(n_1013),
.A3(n_1014),
.B(n_1010),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2081),
.B(n_624),
.Y(n_2387)
);

AOI21x1_ASAP7_75t_L g2388 ( 
.A1(n_2210),
.A2(n_1014),
.B(n_1013),
.Y(n_2388)
);

BUFx2_ASAP7_75t_L g2389 ( 
.A(n_2089),
.Y(n_2389)
);

OAI21x1_ASAP7_75t_L g2390 ( 
.A1(n_2069),
.A2(n_1159),
.B(n_1158),
.Y(n_2390)
);

OAI21x1_ASAP7_75t_L g2391 ( 
.A1(n_2073),
.A2(n_1178),
.B(n_1170),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2071),
.B(n_627),
.Y(n_2392)
);

OAI21x1_ASAP7_75t_L g2393 ( 
.A1(n_1988),
.A2(n_1178),
.B(n_1170),
.Y(n_2393)
);

OAI21x1_ASAP7_75t_L g2394 ( 
.A1(n_1991),
.A2(n_1178),
.B(n_1170),
.Y(n_2394)
);

BUFx3_ASAP7_75t_L g2395 ( 
.A(n_2102),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2017),
.Y(n_2396)
);

BUFx6f_ASAP7_75t_L g2397 ( 
.A(n_2033),
.Y(n_2397)
);

INVx2_ASAP7_75t_SL g2398 ( 
.A(n_2009),
.Y(n_2398)
);

AOI21xp5_ASAP7_75t_L g2399 ( 
.A1(n_2162),
.A2(n_1209),
.B(n_1233),
.Y(n_2399)
);

HB1xp67_ASAP7_75t_L g2400 ( 
.A(n_1989),
.Y(n_2400)
);

A2O1A1Ixp33_ASAP7_75t_L g2401 ( 
.A1(n_2127),
.A2(n_698),
.B(n_711),
.C(n_694),
.Y(n_2401)
);

OAI21x1_ASAP7_75t_L g2402 ( 
.A1(n_1992),
.A2(n_1220),
.B(n_1042),
.Y(n_2402)
);

AOI21xp5_ASAP7_75t_L g2403 ( 
.A1(n_2182),
.A2(n_1209),
.B(n_1233),
.Y(n_2403)
);

AND2x2_ASAP7_75t_SL g2404 ( 
.A(n_2206),
.B(n_2101),
.Y(n_2404)
);

NOR3xp33_ASAP7_75t_L g2405 ( 
.A(n_2148),
.B(n_711),
.C(n_698),
.Y(n_2405)
);

AOI21xp5_ASAP7_75t_L g2406 ( 
.A1(n_2182),
.A2(n_1233),
.B(n_1520),
.Y(n_2406)
);

AO31x2_ASAP7_75t_L g2407 ( 
.A1(n_2025),
.A2(n_1042),
.A3(n_1043),
.B(n_1026),
.Y(n_2407)
);

AOI21xp5_ASAP7_75t_L g2408 ( 
.A1(n_2188),
.A2(n_2210),
.B(n_2208),
.Y(n_2408)
);

AO31x2_ASAP7_75t_L g2409 ( 
.A1(n_2027),
.A2(n_1043),
.A3(n_1045),
.B(n_1026),
.Y(n_2409)
);

INVx1_ASAP7_75t_SL g2410 ( 
.A(n_2061),
.Y(n_2410)
);

INVx3_ASAP7_75t_L g2411 ( 
.A(n_2003),
.Y(n_2411)
);

AOI21x1_ASAP7_75t_L g2412 ( 
.A1(n_2030),
.A2(n_1047),
.B(n_1045),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2031),
.Y(n_2413)
);

OAI21x1_ASAP7_75t_L g2414 ( 
.A1(n_2001),
.A2(n_1220),
.B(n_1047),
.Y(n_2414)
);

OAI21x1_ASAP7_75t_L g2415 ( 
.A1(n_2004),
.A2(n_2020),
.B(n_2016),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2034),
.Y(n_2416)
);

OAI21xp5_ASAP7_75t_L g2417 ( 
.A1(n_2188),
.A2(n_1431),
.B(n_1220),
.Y(n_2417)
);

AND2x4_ASAP7_75t_L g2418 ( 
.A(n_1998),
.B(n_908),
.Y(n_2418)
);

AOI21xp5_ASAP7_75t_L g2419 ( 
.A1(n_2173),
.A2(n_1233),
.B(n_1098),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2039),
.Y(n_2420)
);

AOI21xp5_ASAP7_75t_L g2421 ( 
.A1(n_2173),
.A2(n_1098),
.B(n_1078),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2139),
.B(n_629),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2052),
.B(n_631),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2061),
.B(n_636),
.Y(n_2424)
);

OAI21x1_ASAP7_75t_L g2425 ( 
.A1(n_2045),
.A2(n_910),
.B(n_909),
.Y(n_2425)
);

OAI21xp33_ASAP7_75t_L g2426 ( 
.A1(n_2113),
.A2(n_639),
.B(n_638),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2119),
.B(n_640),
.Y(n_2427)
);

OAI21xp5_ASAP7_75t_L g2428 ( 
.A1(n_2048),
.A2(n_1431),
.B(n_910),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2119),
.B(n_909),
.Y(n_2429)
);

AOI21xp5_ASAP7_75t_L g2430 ( 
.A1(n_2173),
.A2(n_1098),
.B(n_1078),
.Y(n_2430)
);

AOI21xp5_ASAP7_75t_L g2431 ( 
.A1(n_2116),
.A2(n_1098),
.B(n_1078),
.Y(n_2431)
);

AND2x4_ASAP7_75t_L g2432 ( 
.A(n_2006),
.B(n_912),
.Y(n_2432)
);

OAI21x1_ASAP7_75t_L g2433 ( 
.A1(n_2070),
.A2(n_2105),
.B(n_2046),
.Y(n_2433)
);

AOI21xp5_ASAP7_75t_L g2434 ( 
.A1(n_2116),
.A2(n_1109),
.B(n_1078),
.Y(n_2434)
);

OAI21x1_ASAP7_75t_L g2435 ( 
.A1(n_2105),
.A2(n_915),
.B(n_912),
.Y(n_2435)
);

AOI21xp5_ASAP7_75t_SL g2436 ( 
.A1(n_2157),
.A2(n_1113),
.B(n_1109),
.Y(n_2436)
);

AOI21xp5_ASAP7_75t_L g2437 ( 
.A1(n_2169),
.A2(n_1113),
.B(n_1109),
.Y(n_2437)
);

OAI21x1_ASAP7_75t_L g2438 ( 
.A1(n_2041),
.A2(n_917),
.B(n_915),
.Y(n_2438)
);

AOI21xp5_ASAP7_75t_L g2439 ( 
.A1(n_2169),
.A2(n_1113),
.B(n_1109),
.Y(n_2439)
);

OAI21xp5_ASAP7_75t_L g2440 ( 
.A1(n_2127),
.A2(n_1431),
.B(n_918),
.Y(n_2440)
);

OAI22xp5_ASAP7_75t_L g2441 ( 
.A1(n_2047),
.A2(n_722),
.B1(n_724),
.B2(n_718),
.Y(n_2441)
);

A2O1A1Ixp33_ASAP7_75t_L g2442 ( 
.A1(n_2129),
.A2(n_722),
.B(n_724),
.C(n_718),
.Y(n_2442)
);

AOI22xp5_ASAP7_75t_SL g2443 ( 
.A1(n_2080),
.A2(n_648),
.B1(n_654),
.B2(n_642),
.Y(n_2443)
);

HB1xp67_ASAP7_75t_L g2444 ( 
.A(n_2024),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2057),
.Y(n_2445)
);

AOI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2113),
.A2(n_661),
.B1(n_665),
.B2(n_659),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2014),
.Y(n_2447)
);

OAI21x1_ASAP7_75t_L g2448 ( 
.A1(n_2014),
.A2(n_918),
.B(n_917),
.Y(n_2448)
);

AND2x4_ASAP7_75t_L g2449 ( 
.A(n_2006),
.B(n_725),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_SL g2450 ( 
.A(n_2078),
.B(n_678),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2014),
.B(n_725),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2014),
.B(n_727),
.Y(n_2452)
);

AOI21xp5_ASAP7_75t_L g2453 ( 
.A1(n_2157),
.A2(n_1181),
.B(n_1113),
.Y(n_2453)
);

BUFx6f_ASAP7_75t_L g2454 ( 
.A(n_2033),
.Y(n_2454)
);

AOI21xp33_ASAP7_75t_L g2455 ( 
.A1(n_2204),
.A2(n_2053),
.B(n_2075),
.Y(n_2455)
);

AOI21xp5_ASAP7_75t_L g2456 ( 
.A1(n_2204),
.A2(n_1202),
.B(n_1181),
.Y(n_2456)
);

OAI21xp5_ASAP7_75t_L g2457 ( 
.A1(n_1979),
.A2(n_1431),
.B(n_729),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2014),
.B(n_727),
.Y(n_2458)
);

AOI21xp33_ASAP7_75t_L g2459 ( 
.A1(n_2204),
.A2(n_730),
.B(n_729),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2014),
.Y(n_2460)
);

BUFx4f_ASAP7_75t_L g2461 ( 
.A(n_2101),
.Y(n_2461)
);

AOI21x1_ASAP7_75t_L g2462 ( 
.A1(n_2050),
.A2(n_886),
.B(n_885),
.Y(n_2462)
);

OR2x6_ASAP7_75t_L g2463 ( 
.A(n_2204),
.B(n_730),
.Y(n_2463)
);

INVx3_ASAP7_75t_SL g2464 ( 
.A(n_2076),
.Y(n_2464)
);

AO31x2_ASAP7_75t_L g2465 ( 
.A1(n_2053),
.A2(n_734),
.A3(n_737),
.B(n_732),
.Y(n_2465)
);

AOI21xp5_ASAP7_75t_L g2466 ( 
.A1(n_2197),
.A2(n_1202),
.B(n_1181),
.Y(n_2466)
);

NOR2x1_ASAP7_75t_L g2467 ( 
.A(n_2055),
.B(n_732),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_1979),
.B(n_734),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2058),
.B(n_2076),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2003),
.Y(n_2470)
);

OAI21xp5_ASAP7_75t_L g2471 ( 
.A1(n_1979),
.A2(n_1431),
.B(n_738),
.Y(n_2471)
);

AOI21xp5_ASAP7_75t_L g2472 ( 
.A1(n_2197),
.A2(n_1202),
.B(n_1181),
.Y(n_2472)
);

OAI21x1_ASAP7_75t_L g2473 ( 
.A1(n_1979),
.A2(n_886),
.B(n_885),
.Y(n_2473)
);

INVx2_ASAP7_75t_SL g2474 ( 
.A(n_2022),
.Y(n_2474)
);

AOI22xp5_ASAP7_75t_L g2475 ( 
.A1(n_2161),
.A2(n_668),
.B1(n_671),
.B2(n_667),
.Y(n_2475)
);

OAI21x1_ASAP7_75t_L g2476 ( 
.A1(n_1979),
.A2(n_891),
.B(n_888),
.Y(n_2476)
);

AOI21xp5_ASAP7_75t_L g2477 ( 
.A1(n_2050),
.A2(n_1214),
.B(n_1202),
.Y(n_2477)
);

BUFx12f_ASAP7_75t_L g2478 ( 
.A(n_2148),
.Y(n_2478)
);

AND2x2_ASAP7_75t_L g2479 ( 
.A(n_2120),
.B(n_2064),
.Y(n_2479)
);

A2O1A1Ixp33_ASAP7_75t_L g2480 ( 
.A1(n_2120),
.A2(n_738),
.B(n_743),
.C(n_737),
.Y(n_2480)
);

INVx3_ASAP7_75t_L g2481 ( 
.A(n_2305),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2232),
.Y(n_2482)
);

BUFx3_ASAP7_75t_L g2483 ( 
.A(n_2351),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2420),
.Y(n_2484)
);

NOR2xp67_ASAP7_75t_SL g2485 ( 
.A(n_2478),
.B(n_2055),
.Y(n_2485)
);

BUFx8_ASAP7_75t_L g2486 ( 
.A(n_2380),
.Y(n_2486)
);

OAI22xp33_ASAP7_75t_L g2487 ( 
.A1(n_2297),
.A2(n_2319),
.B1(n_2330),
.B2(n_2283),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2275),
.B(n_2161),
.Y(n_2488)
);

BUFx6f_ASAP7_75t_L g2489 ( 
.A(n_2212),
.Y(n_2489)
);

AOI21xp5_ASAP7_75t_L g2490 ( 
.A1(n_2211),
.A2(n_2023),
.B(n_2003),
.Y(n_2490)
);

O2A1O1Ixp33_ASAP7_75t_L g2491 ( 
.A1(n_2272),
.A2(n_745),
.B(n_751),
.C(n_743),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2445),
.Y(n_2492)
);

AOI21xp5_ASAP7_75t_L g2493 ( 
.A1(n_2258),
.A2(n_2023),
.B(n_2003),
.Y(n_2493)
);

AOI22xp5_ASAP7_75t_L g2494 ( 
.A1(n_2347),
.A2(n_2064),
.B1(n_2021),
.B2(n_2043),
.Y(n_2494)
);

BUFx2_ASAP7_75t_L g2495 ( 
.A(n_2313),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2244),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_L g2497 ( 
.A(n_2378),
.B(n_2042),
.Y(n_2497)
);

HB1xp67_ASAP7_75t_L g2498 ( 
.A(n_2410),
.Y(n_2498)
);

AOI221xp5_ASAP7_75t_L g2499 ( 
.A1(n_2373),
.A2(n_680),
.B1(n_686),
.B2(n_684),
.C(n_677),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2273),
.Y(n_2500)
);

HB1xp67_ASAP7_75t_L g2501 ( 
.A(n_2410),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2215),
.B(n_2007),
.Y(n_2502)
);

INVx3_ASAP7_75t_L g2503 ( 
.A(n_2305),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_2317),
.B(n_2100),
.Y(n_2504)
);

NAND2x1p5_ASAP7_75t_L g2505 ( 
.A(n_2362),
.B(n_2021),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_SL g2506 ( 
.A(n_2294),
.B(n_2135),
.Y(n_2506)
);

AOI21x1_ASAP7_75t_L g2507 ( 
.A1(n_2412),
.A2(n_891),
.B(n_888),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2254),
.B(n_2028),
.Y(n_2508)
);

HB1xp67_ASAP7_75t_L g2509 ( 
.A(n_2400),
.Y(n_2509)
);

AND2x6_ASAP7_75t_L g2510 ( 
.A(n_2447),
.B(n_2023),
.Y(n_2510)
);

INVxp67_ASAP7_75t_L g2511 ( 
.A(n_2323),
.Y(n_2511)
);

HB1xp67_ASAP7_75t_L g2512 ( 
.A(n_2323),
.Y(n_2512)
);

BUFx6f_ASAP7_75t_L g2513 ( 
.A(n_2212),
.Y(n_2513)
);

INVx2_ASAP7_75t_SL g2514 ( 
.A(n_2395),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2215),
.B(n_2288),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2304),
.Y(n_2516)
);

INVx2_ASAP7_75t_SL g2517 ( 
.A(n_2252),
.Y(n_2517)
);

AND2x4_ASAP7_75t_L g2518 ( 
.A(n_2479),
.B(n_2028),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_2320),
.Y(n_2519)
);

NAND2x1_ASAP7_75t_L g2520 ( 
.A(n_2362),
.B(n_2091),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2396),
.Y(n_2521)
);

BUFx2_ASAP7_75t_L g2522 ( 
.A(n_2307),
.Y(n_2522)
);

OR2x6_ASAP7_75t_L g2523 ( 
.A(n_2408),
.B(n_2043),
.Y(n_2523)
);

CKINVDCx5p33_ASAP7_75t_R g2524 ( 
.A(n_2309),
.Y(n_2524)
);

AOI22xp5_ASAP7_75t_L g2525 ( 
.A1(n_2261),
.A2(n_2109),
.B1(n_2029),
.B2(n_2035),
.Y(n_2525)
);

OAI21x1_ASAP7_75t_L g2526 ( 
.A1(n_2390),
.A2(n_895),
.B(n_892),
.Y(n_2526)
);

INVxp67_ASAP7_75t_L g2527 ( 
.A(n_2356),
.Y(n_2527)
);

BUFx3_ASAP7_75t_L g2528 ( 
.A(n_2350),
.Y(n_2528)
);

AOI21xp33_ASAP7_75t_L g2529 ( 
.A1(n_2249),
.A2(n_751),
.B(n_745),
.Y(n_2529)
);

AOI22xp5_ASAP7_75t_L g2530 ( 
.A1(n_2450),
.A2(n_2029),
.B1(n_2035),
.B2(n_2007),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2413),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2339),
.Y(n_2532)
);

AOI22xp5_ASAP7_75t_L g2533 ( 
.A1(n_2346),
.A2(n_2381),
.B1(n_2312),
.B2(n_2297),
.Y(n_2533)
);

AOI221xp5_ASAP7_75t_L g2534 ( 
.A1(n_2373),
.A2(n_689),
.B1(n_695),
.B2(n_693),
.C(n_687),
.Y(n_2534)
);

AO21x2_ASAP7_75t_L g2535 ( 
.A1(n_2225),
.A2(n_2255),
.B(n_2326),
.Y(n_2535)
);

INVx1_ASAP7_75t_SL g2536 ( 
.A(n_2444),
.Y(n_2536)
);

INVx3_ASAP7_75t_L g2537 ( 
.A(n_2305),
.Y(n_2537)
);

BUFx3_ASAP7_75t_L g2538 ( 
.A(n_2350),
.Y(n_2538)
);

AOI22xp33_ASAP7_75t_SL g2539 ( 
.A1(n_2319),
.A2(n_2135),
.B1(n_2108),
.B2(n_2185),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_L g2540 ( 
.A(n_2469),
.B(n_700),
.Y(n_2540)
);

INVx1_ASAP7_75t_SL g2541 ( 
.A(n_2257),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2416),
.Y(n_2542)
);

OAI21xp5_ASAP7_75t_L g2543 ( 
.A1(n_2243),
.A2(n_2029),
.B(n_2007),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2249),
.B(n_2007),
.Y(n_2544)
);

INVx5_ASAP7_75t_L g2545 ( 
.A(n_2463),
.Y(n_2545)
);

INVx2_ASAP7_75t_SL g2546 ( 
.A(n_2398),
.Y(n_2546)
);

AND2x4_ASAP7_75t_L g2547 ( 
.A(n_2333),
.B(n_2023),
.Y(n_2547)
);

AOI21xp33_ASAP7_75t_SL g2548 ( 
.A1(n_2405),
.A2(n_761),
.B(n_760),
.Y(n_2548)
);

AOI21xp5_ASAP7_75t_L g2549 ( 
.A1(n_2281),
.A2(n_2079),
.B(n_2044),
.Y(n_2549)
);

BUFx3_ASAP7_75t_L g2550 ( 
.A(n_2350),
.Y(n_2550)
);

HB1xp67_ASAP7_75t_L g2551 ( 
.A(n_2470),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2217),
.B(n_2007),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2265),
.Y(n_2553)
);

AOI21xp5_ASAP7_75t_SL g2554 ( 
.A1(n_2303),
.A2(n_2316),
.B(n_2306),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2359),
.B(n_2108),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2217),
.B(n_2029),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2265),
.Y(n_2557)
);

HB1xp67_ASAP7_75t_L g2558 ( 
.A(n_2230),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2265),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2349),
.B(n_2029),
.Y(n_2560)
);

AOI21xp5_ASAP7_75t_L g2561 ( 
.A1(n_2228),
.A2(n_2079),
.B(n_2044),
.Y(n_2561)
);

AOI22xp33_ASAP7_75t_L g2562 ( 
.A1(n_2384),
.A2(n_713),
.B1(n_723),
.B2(n_678),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2375),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2429),
.B(n_2044),
.Y(n_2564)
);

NAND2xp33_ASAP7_75t_L g2565 ( 
.A(n_2248),
.B(n_2049),
.Y(n_2565)
);

INVx3_ASAP7_75t_L g2566 ( 
.A(n_2314),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2257),
.B(n_2035),
.Y(n_2567)
);

BUFx2_ASAP7_75t_L g2568 ( 
.A(n_2247),
.Y(n_2568)
);

BUFx6f_ASAP7_75t_L g2569 ( 
.A(n_2212),
.Y(n_2569)
);

INVx5_ASAP7_75t_L g2570 ( 
.A(n_2463),
.Y(n_2570)
);

AOI21xp5_ASAP7_75t_L g2571 ( 
.A1(n_2399),
.A2(n_2079),
.B(n_2044),
.Y(n_2571)
);

CKINVDCx5p33_ASAP7_75t_R g2572 ( 
.A(n_2298),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2407),
.Y(n_2573)
);

AOI21xp5_ASAP7_75t_L g2574 ( 
.A1(n_2292),
.A2(n_2083),
.B(n_2079),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2404),
.B(n_2083),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2271),
.B(n_2083),
.Y(n_2576)
);

BUFx2_ASAP7_75t_L g2577 ( 
.A(n_2247),
.Y(n_2577)
);

AOI22xp5_ASAP7_75t_L g2578 ( 
.A1(n_2426),
.A2(n_2035),
.B1(n_705),
.B2(n_715),
.Y(n_2578)
);

BUFx12f_ASAP7_75t_L g2579 ( 
.A(n_2374),
.Y(n_2579)
);

CKINVDCx5p33_ASAP7_75t_R g2580 ( 
.A(n_2363),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2407),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2415),
.Y(n_2582)
);

AOI22xp33_ASAP7_75t_L g2583 ( 
.A1(n_2384),
.A2(n_713),
.B1(n_723),
.B2(n_678),
.Y(n_2583)
);

BUFx2_ASAP7_75t_L g2584 ( 
.A(n_2247),
.Y(n_2584)
);

O2A1O1Ixp33_ASAP7_75t_L g2585 ( 
.A1(n_2401),
.A2(n_761),
.B(n_767),
.C(n_760),
.Y(n_2585)
);

BUFx3_ASAP7_75t_L g2586 ( 
.A(n_2374),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2433),
.Y(n_2587)
);

AND2x4_ASAP7_75t_L g2588 ( 
.A(n_2314),
.B(n_2083),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_SL g2589 ( 
.A(n_2455),
.B(n_2049),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2407),
.Y(n_2590)
);

BUFx6f_ASAP7_75t_L g2591 ( 
.A(n_2223),
.Y(n_2591)
);

AOI22xp33_ASAP7_75t_L g2592 ( 
.A1(n_2384),
.A2(n_713),
.B1(n_723),
.B2(n_767),
.Y(n_2592)
);

INVx2_ASAP7_75t_SL g2593 ( 
.A(n_2474),
.Y(n_2593)
);

BUFx3_ASAP7_75t_L g2594 ( 
.A(n_2374),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2409),
.Y(n_2595)
);

AND2x4_ASAP7_75t_L g2596 ( 
.A(n_2314),
.B(n_2035),
.Y(n_2596)
);

HB1xp67_ASAP7_75t_L g2597 ( 
.A(n_2463),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2409),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2301),
.B(n_892),
.Y(n_2599)
);

BUFx2_ASAP7_75t_L g2600 ( 
.A(n_2276),
.Y(n_2600)
);

AOI22xp5_ASAP7_75t_L g2601 ( 
.A1(n_2446),
.A2(n_716),
.B1(n_719),
.B2(n_706),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2259),
.B(n_2091),
.Y(n_2602)
);

AND2x4_ASAP7_75t_L g2603 ( 
.A(n_2276),
.B(n_2091),
.Y(n_2603)
);

BUFx2_ASAP7_75t_L g2604 ( 
.A(n_2276),
.Y(n_2604)
);

AOI21xp5_ASAP7_75t_L g2605 ( 
.A1(n_2219),
.A2(n_1231),
.B(n_1214),
.Y(n_2605)
);

A2O1A1Ixp33_ASAP7_75t_L g2606 ( 
.A1(n_2442),
.A2(n_726),
.B(n_735),
.C(n_733),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2409),
.Y(n_2607)
);

INVx2_ASAP7_75t_SL g2608 ( 
.A(n_2397),
.Y(n_2608)
);

BUFx3_ASAP7_75t_L g2609 ( 
.A(n_2397),
.Y(n_2609)
);

NAND2x1p5_ASAP7_75t_L g2610 ( 
.A(n_2286),
.B(n_1214),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2259),
.B(n_895),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2236),
.Y(n_2612)
);

BUFx4_ASAP7_75t_SL g2613 ( 
.A(n_2379),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2236),
.Y(n_2614)
);

AOI21xp33_ASAP7_75t_L g2615 ( 
.A1(n_2214),
.A2(n_742),
.B(n_736),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2236),
.Y(n_2616)
);

AOI21xp5_ASAP7_75t_L g2617 ( 
.A1(n_2250),
.A2(n_1231),
.B(n_1214),
.Y(n_2617)
);

INVx1_ASAP7_75t_SL g2618 ( 
.A(n_2389),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2235),
.B(n_898),
.Y(n_2619)
);

BUFx2_ASAP7_75t_L g2620 ( 
.A(n_2464),
.Y(n_2620)
);

HB1xp67_ASAP7_75t_L g2621 ( 
.A(n_2235),
.Y(n_2621)
);

NAND2x1_ASAP7_75t_L g2622 ( 
.A(n_2436),
.B(n_2226),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2451),
.Y(n_2623)
);

BUFx8_ASAP7_75t_L g2624 ( 
.A(n_2397),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2451),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2452),
.Y(n_2626)
);

AND2x4_ASAP7_75t_L g2627 ( 
.A(n_2282),
.B(n_325),
.Y(n_2627)
);

HB1xp67_ASAP7_75t_L g2628 ( 
.A(n_2237),
.Y(n_2628)
);

AND2x4_ASAP7_75t_L g2629 ( 
.A(n_2282),
.B(n_2365),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2267),
.Y(n_2630)
);

BUFx6f_ASAP7_75t_L g2631 ( 
.A(n_2223),
.Y(n_2631)
);

OAI21xp5_ASAP7_75t_L g2632 ( 
.A1(n_2225),
.A2(n_899),
.B(n_898),
.Y(n_2632)
);

CKINVDCx8_ASAP7_75t_R g2633 ( 
.A(n_2454),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2322),
.Y(n_2634)
);

AOI21xp5_ASAP7_75t_L g2635 ( 
.A1(n_2269),
.A2(n_1231),
.B(n_996),
.Y(n_2635)
);

A2O1A1Ixp33_ASAP7_75t_L g2636 ( 
.A1(n_2459),
.A2(n_744),
.B(n_747),
.C(n_746),
.Y(n_2636)
);

AOI21xp5_ASAP7_75t_L g2637 ( 
.A1(n_2262),
.A2(n_1231),
.B(n_996),
.Y(n_2637)
);

INVx3_ASAP7_75t_L g2638 ( 
.A(n_2461),
.Y(n_2638)
);

AOI22xp33_ASAP7_75t_L g2639 ( 
.A1(n_2384),
.A2(n_2449),
.B1(n_2360),
.B2(n_2467),
.Y(n_2639)
);

BUFx3_ASAP7_75t_L g2640 ( 
.A(n_2454),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2452),
.Y(n_2641)
);

BUFx3_ASAP7_75t_L g2642 ( 
.A(n_2454),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2237),
.B(n_899),
.Y(n_2643)
);

BUFx3_ASAP7_75t_L g2644 ( 
.A(n_2223),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2338),
.B(n_748),
.Y(n_2645)
);

BUFx10_ASAP7_75t_L g2646 ( 
.A(n_2418),
.Y(n_2646)
);

INVx2_ASAP7_75t_SL g2647 ( 
.A(n_2461),
.Y(n_2647)
);

AO32x1_ASAP7_75t_L g2648 ( 
.A1(n_2360),
.A2(n_723),
.A3(n_757),
.B1(n_919),
.B2(n_7),
.Y(n_2648)
);

AND2x4_ASAP7_75t_L g2649 ( 
.A(n_2344),
.B(n_327),
.Y(n_2649)
);

BUFx4_ASAP7_75t_SL g2650 ( 
.A(n_2290),
.Y(n_2650)
);

AOI21xp5_ASAP7_75t_L g2651 ( 
.A1(n_2293),
.A2(n_996),
.B(n_963),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2253),
.B(n_763),
.Y(n_2652)
);

AND2x4_ASAP7_75t_L g2653 ( 
.A(n_2344),
.B(n_329),
.Y(n_2653)
);

BUFx2_ASAP7_75t_SL g2654 ( 
.A(n_2418),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2253),
.B(n_2227),
.Y(n_2655)
);

AOI22xp33_ASAP7_75t_L g2656 ( 
.A1(n_2449),
.A2(n_765),
.B1(n_766),
.B2(n_764),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2458),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2458),
.Y(n_2658)
);

OAI22xp5_ASAP7_75t_L g2659 ( 
.A1(n_2227),
.A2(n_9),
.B1(n_4),
.B2(n_6),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2329),
.Y(n_2660)
);

BUFx12f_ASAP7_75t_L g2661 ( 
.A(n_2432),
.Y(n_2661)
);

HB1xp67_ASAP7_75t_L g2662 ( 
.A(n_2291),
.Y(n_2662)
);

HB1xp67_ASAP7_75t_L g2663 ( 
.A(n_2299),
.Y(n_2663)
);

AOI21xp5_ASAP7_75t_L g2664 ( 
.A1(n_2385),
.A2(n_996),
.B(n_963),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2411),
.Y(n_2665)
);

BUFx6f_ASAP7_75t_L g2666 ( 
.A(n_2334),
.Y(n_2666)
);

OR2x2_ASAP7_75t_SL g2667 ( 
.A(n_2468),
.B(n_4),
.Y(n_2667)
);

INVx3_ASAP7_75t_L g2668 ( 
.A(n_2411),
.Y(n_2668)
);

NOR2xp67_ASAP7_75t_SL g2669 ( 
.A(n_2263),
.B(n_967),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2231),
.B(n_6),
.Y(n_2670)
);

CKINVDCx20_ASAP7_75t_R g2671 ( 
.A(n_2392),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2432),
.B(n_330),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2310),
.Y(n_2673)
);

NAND2x1p5_ASAP7_75t_L g2674 ( 
.A(n_2222),
.B(n_967),
.Y(n_2674)
);

AOI22xp33_ASAP7_75t_SL g2675 ( 
.A1(n_2443),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_2675)
);

NOR2xp67_ASAP7_75t_SL g2676 ( 
.A(n_2222),
.B(n_967),
.Y(n_2676)
);

AOI21xp5_ASAP7_75t_L g2677 ( 
.A1(n_2315),
.A2(n_996),
.B(n_963),
.Y(n_2677)
);

OAI22xp5_ASAP7_75t_L g2678 ( 
.A1(n_2231),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_2678)
);

AOI21xp5_ASAP7_75t_L g2679 ( 
.A1(n_2340),
.A2(n_996),
.B(n_963),
.Y(n_2679)
);

BUFx12f_ASAP7_75t_L g2680 ( 
.A(n_2334),
.Y(n_2680)
);

BUFx2_ASAP7_75t_L g2681 ( 
.A(n_2299),
.Y(n_2681)
);

AND2x4_ASAP7_75t_L g2682 ( 
.A(n_2345),
.B(n_335),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2310),
.Y(n_2683)
);

BUFx3_ASAP7_75t_L g2684 ( 
.A(n_2427),
.Y(n_2684)
);

AND2x4_ASAP7_75t_L g2685 ( 
.A(n_2287),
.B(n_2295),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2465),
.B(n_336),
.Y(n_2686)
);

OAI22x1_ASAP7_75t_L g2687 ( 
.A1(n_2475),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_2687)
);

BUFx4_ASAP7_75t_SL g2688 ( 
.A(n_2290),
.Y(n_2688)
);

BUFx6f_ASAP7_75t_L g2689 ( 
.A(n_2285),
.Y(n_2689)
);

AND2x2_ASAP7_75t_L g2690 ( 
.A(n_2465),
.B(n_337),
.Y(n_2690)
);

AOI21xp5_ASAP7_75t_L g2691 ( 
.A1(n_2341),
.A2(n_963),
.B(n_930),
.Y(n_2691)
);

OR2x2_ASAP7_75t_L g2692 ( 
.A(n_2423),
.B(n_16),
.Y(n_2692)
);

AND2x4_ASAP7_75t_L g2693 ( 
.A(n_2287),
.B(n_342),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2310),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2324),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2234),
.B(n_18),
.Y(n_2696)
);

INVx2_ASAP7_75t_L g2697 ( 
.A(n_2425),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2465),
.B(n_343),
.Y(n_2698)
);

OR2x2_ASAP7_75t_L g2699 ( 
.A(n_2424),
.B(n_19),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2324),
.Y(n_2700)
);

AND2x4_ASAP7_75t_L g2701 ( 
.A(n_2295),
.B(n_2290),
.Y(n_2701)
);

AOI21xp33_ASAP7_75t_L g2702 ( 
.A1(n_2234),
.A2(n_21),
.B(n_22),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2240),
.Y(n_2703)
);

AND2x4_ASAP7_75t_L g2704 ( 
.A(n_2289),
.B(n_344),
.Y(n_2704)
);

AOI21xp5_ASAP7_75t_L g2705 ( 
.A1(n_2341),
.A2(n_963),
.B(n_930),
.Y(n_2705)
);

INVx2_ASAP7_75t_SL g2706 ( 
.A(n_2422),
.Y(n_2706)
);

INVx3_ASAP7_75t_SL g2707 ( 
.A(n_2289),
.Y(n_2707)
);

OR2x2_ASAP7_75t_L g2708 ( 
.A(n_2284),
.B(n_21),
.Y(n_2708)
);

AOI22xp33_ASAP7_75t_L g2709 ( 
.A1(n_2459),
.A2(n_1431),
.B1(n_1274),
.B2(n_1244),
.Y(n_2709)
);

AND2x4_ASAP7_75t_L g2710 ( 
.A(n_2368),
.B(n_347),
.Y(n_2710)
);

CKINVDCx11_ASAP7_75t_R g2711 ( 
.A(n_2441),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2279),
.B(n_22),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2240),
.Y(n_2713)
);

INVx5_ASAP7_75t_L g2714 ( 
.A(n_2460),
.Y(n_2714)
);

O2A1O1Ixp5_ASAP7_75t_SL g2715 ( 
.A1(n_2441),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_2715)
);

NOR2xp33_ASAP7_75t_L g2716 ( 
.A(n_2387),
.B(n_2455),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2324),
.Y(n_2717)
);

NAND2x1p5_ASAP7_75t_L g2718 ( 
.A(n_2224),
.B(n_967),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2354),
.Y(n_2719)
);

INVx4_ASAP7_75t_L g2720 ( 
.A(n_2285),
.Y(n_2720)
);

BUFx6f_ASAP7_75t_L g2721 ( 
.A(n_2308),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2246),
.Y(n_2722)
);

OAI22xp5_ASAP7_75t_SL g2723 ( 
.A1(n_2300),
.A2(n_27),
.B1(n_23),
.B2(n_26),
.Y(n_2723)
);

INVx4_ASAP7_75t_L g2724 ( 
.A(n_2308),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2279),
.B(n_26),
.Y(n_2725)
);

BUFx2_ASAP7_75t_SL g2726 ( 
.A(n_2266),
.Y(n_2726)
);

INVx3_ASAP7_75t_L g2727 ( 
.A(n_2280),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2302),
.B(n_28),
.Y(n_2728)
);

OA21x2_ASAP7_75t_L g2729 ( 
.A1(n_2213),
.A2(n_1431),
.B(n_1274),
.Y(n_2729)
);

AND2x4_ASAP7_75t_L g2730 ( 
.A(n_2229),
.B(n_349),
.Y(n_2730)
);

INVx5_ASAP7_75t_L g2731 ( 
.A(n_2221),
.Y(n_2731)
);

HB1xp67_ASAP7_75t_L g2732 ( 
.A(n_2246),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2251),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2354),
.Y(n_2734)
);

AOI221x1_ASAP7_75t_L g2735 ( 
.A1(n_2343),
.A2(n_976),
.B1(n_979),
.B2(n_972),
.C(n_967),
.Y(n_2735)
);

AOI21xp33_ASAP7_75t_L g2736 ( 
.A1(n_2376),
.A2(n_29),
.B(n_30),
.Y(n_2736)
);

HB1xp67_ASAP7_75t_L g2737 ( 
.A(n_2251),
.Y(n_2737)
);

AND2x4_ASAP7_75t_L g2738 ( 
.A(n_2468),
.B(n_354),
.Y(n_2738)
);

INVx1_ASAP7_75t_SL g2739 ( 
.A(n_2274),
.Y(n_2739)
);

NAND2x1_ASAP7_75t_L g2740 ( 
.A(n_2296),
.B(n_972),
.Y(n_2740)
);

BUFx6f_ASAP7_75t_L g2741 ( 
.A(n_2369),
.Y(n_2741)
);

BUFx6f_ASAP7_75t_L g2742 ( 
.A(n_2239),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2302),
.B(n_31),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2438),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2354),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2245),
.Y(n_2746)
);

AND2x4_ASAP7_75t_L g2747 ( 
.A(n_2260),
.B(n_355),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2361),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2386),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2482),
.Y(n_2750)
);

OAI21x1_ASAP7_75t_L g2751 ( 
.A1(n_2605),
.A2(n_2218),
.B(n_2241),
.Y(n_2751)
);

OAI21x1_ASAP7_75t_L g2752 ( 
.A1(n_2605),
.A2(n_2216),
.B(n_2264),
.Y(n_2752)
);

INVxp67_ASAP7_75t_L g2753 ( 
.A(n_2522),
.Y(n_2753)
);

A2O1A1Ixp33_ASAP7_75t_L g2754 ( 
.A1(n_2529),
.A2(n_2457),
.B(n_2471),
.C(n_2440),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2496),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2500),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2576),
.B(n_2508),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2739),
.B(n_2348),
.Y(n_2758)
);

AND2x4_ASAP7_75t_L g2759 ( 
.A(n_2523),
.B(n_2233),
.Y(n_2759)
);

INVx2_ASAP7_75t_SL g2760 ( 
.A(n_2483),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2739),
.B(n_2662),
.Y(n_2761)
);

O2A1O1Ixp33_ASAP7_75t_L g2762 ( 
.A1(n_2491),
.A2(n_2382),
.B(n_2480),
.C(n_2440),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2516),
.Y(n_2763)
);

AOI21xp5_ASAP7_75t_L g2764 ( 
.A1(n_2554),
.A2(n_2221),
.B(n_2325),
.Y(n_2764)
);

CKINVDCx8_ASAP7_75t_R g2765 ( 
.A(n_2580),
.Y(n_2765)
);

AOI22xp33_ASAP7_75t_L g2766 ( 
.A1(n_2711),
.A2(n_2529),
.B1(n_2675),
.B2(n_2723),
.Y(n_2766)
);

AOI22xp5_ASAP7_75t_SL g2767 ( 
.A1(n_2497),
.A2(n_2233),
.B1(n_2296),
.B2(n_2348),
.Y(n_2767)
);

BUFx3_ASAP7_75t_L g2768 ( 
.A(n_2624),
.Y(n_2768)
);

NAND3xp33_ASAP7_75t_L g2769 ( 
.A(n_2491),
.B(n_2260),
.C(n_2376),
.Y(n_2769)
);

OAI22xp5_ASAP7_75t_L g2770 ( 
.A1(n_2539),
.A2(n_2332),
.B1(n_2311),
.B2(n_2457),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2521),
.Y(n_2771)
);

OAI21x1_ASAP7_75t_L g2772 ( 
.A1(n_2617),
.A2(n_2337),
.B(n_2277),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2531),
.Y(n_2773)
);

BUFx5_ASAP7_75t_L g2774 ( 
.A(n_2573),
.Y(n_2774)
);

OR2x2_ASAP7_75t_L g2775 ( 
.A(n_2541),
.B(n_2326),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2512),
.B(n_2238),
.Y(n_2776)
);

INVx3_ASAP7_75t_L g2777 ( 
.A(n_2685),
.Y(n_2777)
);

INVx1_ASAP7_75t_SL g2778 ( 
.A(n_2495),
.Y(n_2778)
);

OAI21x1_ASAP7_75t_SL g2779 ( 
.A1(n_2712),
.A2(n_2255),
.B(n_2335),
.Y(n_2779)
);

OR2x6_ASAP7_75t_L g2780 ( 
.A(n_2523),
.B(n_2270),
.Y(n_2780)
);

OAI21x1_ASAP7_75t_L g2781 ( 
.A1(n_2617),
.A2(n_2268),
.B(n_2242),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2542),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2621),
.Y(n_2783)
);

AO21x2_ASAP7_75t_L g2784 ( 
.A1(n_2581),
.A2(n_2238),
.B(n_2335),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2575),
.B(n_2220),
.Y(n_2785)
);

OAI21x1_ASAP7_75t_L g2786 ( 
.A1(n_2651),
.A2(n_2391),
.B(n_2448),
.Y(n_2786)
);

HB1xp67_ASAP7_75t_L g2787 ( 
.A(n_2558),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2498),
.B(n_2311),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2501),
.B(n_2318),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2628),
.Y(n_2790)
);

INVx3_ASAP7_75t_L g2791 ( 
.A(n_2685),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2612),
.Y(n_2792)
);

CKINVDCx6p67_ASAP7_75t_R g2793 ( 
.A(n_2579),
.Y(n_2793)
);

INVxp67_ASAP7_75t_SL g2794 ( 
.A(n_2553),
.Y(n_2794)
);

AND2x2_ASAP7_75t_L g2795 ( 
.A(n_2564),
.B(n_2220),
.Y(n_2795)
);

NOR2xp33_ASAP7_75t_L g2796 ( 
.A(n_2716),
.B(n_2462),
.Y(n_2796)
);

OAI22xp5_ASAP7_75t_L g2797 ( 
.A1(n_2539),
.A2(n_2471),
.B1(n_2318),
.B2(n_2355),
.Y(n_2797)
);

O2A1O1Ixp33_ASAP7_75t_SL g2798 ( 
.A1(n_2736),
.A2(n_2487),
.B(n_2589),
.C(n_2659),
.Y(n_2798)
);

AOI22xp5_ASAP7_75t_L g2799 ( 
.A1(n_2533),
.A2(n_2327),
.B1(n_2367),
.B2(n_2355),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2614),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2509),
.Y(n_2801)
);

NOR2xp33_ASAP7_75t_L g2802 ( 
.A(n_2488),
.B(n_2388),
.Y(n_2802)
);

BUFx2_ASAP7_75t_L g2803 ( 
.A(n_2624),
.Y(n_2803)
);

OAI21x1_ASAP7_75t_L g2804 ( 
.A1(n_2651),
.A2(n_2394),
.B(n_2393),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2518),
.B(n_2220),
.Y(n_2805)
);

OAI21x1_ASAP7_75t_L g2806 ( 
.A1(n_2561),
.A2(n_2372),
.B(n_2473),
.Y(n_2806)
);

OAI21x1_ASAP7_75t_L g2807 ( 
.A1(n_2490),
.A2(n_2383),
.B(n_2331),
.Y(n_2807)
);

INVx3_ASAP7_75t_L g2808 ( 
.A(n_2701),
.Y(n_2808)
);

OAI21x1_ASAP7_75t_L g2809 ( 
.A1(n_2490),
.A2(n_2476),
.B(n_2453),
.Y(n_2809)
);

AND2x2_ASAP7_75t_L g2810 ( 
.A(n_2518),
.B(n_2367),
.Y(n_2810)
);

HB1xp67_ASAP7_75t_L g2811 ( 
.A(n_2557),
.Y(n_2811)
);

AOI22xp33_ASAP7_75t_L g2812 ( 
.A1(n_2675),
.A2(n_2327),
.B1(n_2371),
.B2(n_2361),
.Y(n_2812)
);

AND2x2_ASAP7_75t_L g2813 ( 
.A(n_2511),
.B(n_2417),
.Y(n_2813)
);

AOI22xp33_ASAP7_75t_L g2814 ( 
.A1(n_2615),
.A2(n_2371),
.B1(n_2353),
.B2(n_2336),
.Y(n_2814)
);

OAI21xp5_ASAP7_75t_L g2815 ( 
.A1(n_2615),
.A2(n_2435),
.B(n_2403),
.Y(n_2815)
);

OAI21x1_ASAP7_75t_L g2816 ( 
.A1(n_2561),
.A2(n_2718),
.B(n_2595),
.Y(n_2816)
);

OAI21x1_ASAP7_75t_L g2817 ( 
.A1(n_2718),
.A2(n_2598),
.B(n_2590),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2541),
.B(n_2321),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2732),
.Y(n_2819)
);

AO31x2_ASAP7_75t_L g2820 ( 
.A1(n_2607),
.A2(n_2456),
.A3(n_2419),
.B(n_2430),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2737),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2616),
.Y(n_2822)
);

OR2x2_ASAP7_75t_L g2823 ( 
.A(n_2655),
.B(n_2386),
.Y(n_2823)
);

OAI21x1_ASAP7_75t_L g2824 ( 
.A1(n_2543),
.A2(n_2342),
.B(n_2402),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2719),
.Y(n_2825)
);

NAND2xp33_ASAP7_75t_L g2826 ( 
.A(n_2545),
.B(n_2417),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2511),
.B(n_2386),
.Y(n_2827)
);

CKINVDCx5p33_ASAP7_75t_R g2828 ( 
.A(n_2524),
.Y(n_2828)
);

INVx3_ASAP7_75t_L g2829 ( 
.A(n_2701),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2551),
.Y(n_2830)
);

OAI22x1_ASAP7_75t_L g2831 ( 
.A1(n_2618),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_2831)
);

OR2x2_ASAP7_75t_L g2832 ( 
.A(n_2655),
.B(n_2536),
.Y(n_2832)
);

OAI21x1_ASAP7_75t_L g2833 ( 
.A1(n_2543),
.A2(n_2414),
.B(n_2256),
.Y(n_2833)
);

CKINVDCx12_ASAP7_75t_R g2834 ( 
.A(n_2555),
.Y(n_2834)
);

AND2x4_ASAP7_75t_L g2835 ( 
.A(n_2523),
.B(n_2328),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2734),
.Y(n_2836)
);

NOR2xp33_ASAP7_75t_L g2837 ( 
.A(n_2488),
.B(n_2377),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2484),
.Y(n_2838)
);

AO32x2_ASAP7_75t_L g2839 ( 
.A1(n_2659),
.A2(n_2278),
.A3(n_35),
.B1(n_32),
.B2(n_33),
.Y(n_2839)
);

AOI22xp33_ASAP7_75t_L g2840 ( 
.A1(n_2687),
.A2(n_2364),
.B1(n_2428),
.B2(n_2370),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2492),
.Y(n_2841)
);

CKINVDCx16_ASAP7_75t_R g2842 ( 
.A(n_2671),
.Y(n_2842)
);

OA21x2_ASAP7_75t_L g2843 ( 
.A1(n_2515),
.A2(n_2358),
.B(n_2357),
.Y(n_2843)
);

AO21x2_ASAP7_75t_L g2844 ( 
.A1(n_2749),
.A2(n_2421),
.B(n_2477),
.Y(n_2844)
);

OR2x2_ASAP7_75t_L g2845 ( 
.A(n_2536),
.B(n_2366),
.Y(n_2845)
);

OA21x2_ASAP7_75t_L g2846 ( 
.A1(n_2515),
.A2(n_2352),
.B(n_2428),
.Y(n_2846)
);

AO221x2_ASAP7_75t_L g2847 ( 
.A1(n_2678),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.C(n_39),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2559),
.Y(n_2848)
);

OAI21xp5_ASAP7_75t_L g2849 ( 
.A1(n_2645),
.A2(n_2434),
.B(n_2431),
.Y(n_2849)
);

OAI21x1_ASAP7_75t_L g2850 ( 
.A1(n_2740),
.A2(n_2439),
.B(n_2437),
.Y(n_2850)
);

OAI21xp5_ASAP7_75t_L g2851 ( 
.A1(n_2645),
.A2(n_2406),
.B(n_2466),
.Y(n_2851)
);

AOI21xp5_ASAP7_75t_L g2852 ( 
.A1(n_2679),
.A2(n_2622),
.B(n_2535),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2568),
.B(n_36),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2745),
.Y(n_2854)
);

AND2x4_ASAP7_75t_L g2855 ( 
.A(n_2629),
.B(n_2472),
.Y(n_2855)
);

OAI21xp5_ASAP7_75t_L g2856 ( 
.A1(n_2606),
.A2(n_1274),
.B(n_1244),
.Y(n_2856)
);

OAI22xp5_ASAP7_75t_L g2857 ( 
.A1(n_2639),
.A2(n_40),
.B1(n_37),
.B2(n_38),
.Y(n_2857)
);

OAI21x1_ASAP7_75t_L g2858 ( 
.A1(n_2574),
.A2(n_362),
.B(n_356),
.Y(n_2858)
);

AND2x4_ASAP7_75t_L g2859 ( 
.A(n_2629),
.B(n_363),
.Y(n_2859)
);

OAI21x1_ASAP7_75t_L g2860 ( 
.A1(n_2574),
.A2(n_372),
.B(n_371),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2746),
.Y(n_2861)
);

INVx2_ASAP7_75t_SL g2862 ( 
.A(n_2613),
.Y(n_2862)
);

AND2x2_ASAP7_75t_L g2863 ( 
.A(n_2577),
.B(n_41),
.Y(n_2863)
);

INVx1_ASAP7_75t_SL g2864 ( 
.A(n_2618),
.Y(n_2864)
);

AO21x2_ASAP7_75t_L g2865 ( 
.A1(n_2673),
.A2(n_1274),
.B(n_1244),
.Y(n_2865)
);

A2O1A1Ixp33_ASAP7_75t_L g2866 ( 
.A1(n_2736),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2683),
.Y(n_2867)
);

AO21x2_ASAP7_75t_L g2868 ( 
.A1(n_2694),
.A2(n_1274),
.B(n_1244),
.Y(n_2868)
);

OAI21x1_ASAP7_75t_L g2869 ( 
.A1(n_2549),
.A2(n_378),
.B(n_373),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2527),
.Y(n_2870)
);

OAI21x1_ASAP7_75t_L g2871 ( 
.A1(n_2549),
.A2(n_380),
.B(n_379),
.Y(n_2871)
);

OAI21x1_ASAP7_75t_L g2872 ( 
.A1(n_2695),
.A2(n_383),
.B(n_382),
.Y(n_2872)
);

INVx1_ASAP7_75t_SL g2873 ( 
.A(n_2620),
.Y(n_2873)
);

INVx5_ASAP7_75t_L g2874 ( 
.A(n_2731),
.Y(n_2874)
);

OAI21x1_ASAP7_75t_L g2875 ( 
.A1(n_2700),
.A2(n_387),
.B(n_384),
.Y(n_2875)
);

NAND2x1p5_ASAP7_75t_L g2876 ( 
.A(n_2731),
.B(n_972),
.Y(n_2876)
);

BUFx3_ASAP7_75t_L g2877 ( 
.A(n_2528),
.Y(n_2877)
);

OAI22xp33_ASAP7_75t_L g2878 ( 
.A1(n_2678),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.Y(n_2878)
);

OAI22x1_ASAP7_75t_L g2879 ( 
.A1(n_2525),
.A2(n_48),
.B1(n_44),
.B2(n_46),
.Y(n_2879)
);

OAI21x1_ASAP7_75t_L g2880 ( 
.A1(n_2717),
.A2(n_389),
.B(n_388),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2527),
.Y(n_2881)
);

AO21x2_ASAP7_75t_L g2882 ( 
.A1(n_2712),
.A2(n_1274),
.B(n_1244),
.Y(n_2882)
);

A2O1A1Ixp33_ASAP7_75t_L g2883 ( 
.A1(n_2585),
.A2(n_52),
.B(n_46),
.C(n_51),
.Y(n_2883)
);

OAI21x1_ASAP7_75t_L g2884 ( 
.A1(n_2664),
.A2(n_2677),
.B(n_2507),
.Y(n_2884)
);

OA21x2_ASAP7_75t_L g2885 ( 
.A1(n_2735),
.A2(n_51),
.B(n_52),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2582),
.Y(n_2886)
);

INVx4_ASAP7_75t_L g2887 ( 
.A(n_2707),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2703),
.Y(n_2888)
);

AND2x4_ASAP7_75t_L g2889 ( 
.A(n_2742),
.B(n_392),
.Y(n_2889)
);

OAI21xp5_ASAP7_75t_L g2890 ( 
.A1(n_2585),
.A2(n_394),
.B(n_393),
.Y(n_2890)
);

AND2x4_ASAP7_75t_L g2891 ( 
.A(n_2742),
.B(n_395),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2713),
.Y(n_2892)
);

OAI21x1_ASAP7_75t_L g2893 ( 
.A1(n_2610),
.A2(n_398),
.B(n_396),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2722),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2733),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2519),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2532),
.Y(n_2897)
);

OA21x2_ASAP7_75t_L g2898 ( 
.A1(n_2560),
.A2(n_2502),
.B(n_2544),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2623),
.B(n_53),
.Y(n_2899)
);

AO21x2_ASAP7_75t_L g2900 ( 
.A1(n_2725),
.A2(n_53),
.B(n_54),
.Y(n_2900)
);

NOR2xp33_ASAP7_75t_L g2901 ( 
.A(n_2667),
.B(n_54),
.Y(n_2901)
);

OAI22xp5_ASAP7_75t_L g2902 ( 
.A1(n_2562),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2563),
.Y(n_2903)
);

BUFx3_ASAP7_75t_L g2904 ( 
.A(n_2538),
.Y(n_2904)
);

AOI22xp33_ASAP7_75t_L g2905 ( 
.A1(n_2583),
.A2(n_58),
.B1(n_55),
.B2(n_56),
.Y(n_2905)
);

OA21x2_ASAP7_75t_L g2906 ( 
.A1(n_2560),
.A2(n_58),
.B(n_59),
.Y(n_2906)
);

OA21x2_ASAP7_75t_L g2907 ( 
.A1(n_2502),
.A2(n_59),
.B(n_60),
.Y(n_2907)
);

AO221x2_ASAP7_75t_L g2908 ( 
.A1(n_2725),
.A2(n_63),
.B1(n_60),
.B2(n_62),
.C(n_64),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2587),
.Y(n_2909)
);

CKINVDCx5p33_ASAP7_75t_R g2910 ( 
.A(n_2572),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2630),
.Y(n_2911)
);

NOR2xp33_ASAP7_75t_L g2912 ( 
.A(n_2728),
.B(n_63),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2742),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2625),
.Y(n_2914)
);

CKINVDCx5p33_ASAP7_75t_R g2915 ( 
.A(n_2486),
.Y(n_2915)
);

OA21x2_ASAP7_75t_L g2916 ( 
.A1(n_2544),
.A2(n_64),
.B(n_65),
.Y(n_2916)
);

BUFx6f_ASAP7_75t_L g2917 ( 
.A(n_2489),
.Y(n_2917)
);

INVx2_ASAP7_75t_SL g2918 ( 
.A(n_2546),
.Y(n_2918)
);

AOI22xp5_ASAP7_75t_L g2919 ( 
.A1(n_2706),
.A2(n_976),
.B1(n_979),
.B2(n_972),
.Y(n_2919)
);

OAI22xp5_ASAP7_75t_L g2920 ( 
.A1(n_2592),
.A2(n_70),
.B1(n_67),
.B2(n_68),
.Y(n_2920)
);

BUFx2_ASAP7_75t_L g2921 ( 
.A(n_2584),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2626),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2641),
.Y(n_2923)
);

AO21x2_ASAP7_75t_L g2924 ( 
.A1(n_2493),
.A2(n_67),
.B(n_68),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2657),
.Y(n_2925)
);

O2A1O1Ixp33_ASAP7_75t_L g2926 ( 
.A1(n_2702),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2658),
.Y(n_2927)
);

AO32x2_ASAP7_75t_L g2928 ( 
.A1(n_2724),
.A2(n_71),
.A3(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_2928)
);

OAI21x1_ASAP7_75t_L g2929 ( 
.A1(n_2610),
.A2(n_2664),
.B(n_2677),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2602),
.Y(n_2930)
);

NOR2x1_ASAP7_75t_SL g2931 ( 
.A(n_2731),
.B(n_972),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2634),
.B(n_75),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2602),
.Y(n_2933)
);

INVx4_ASAP7_75t_L g2934 ( 
.A(n_2545),
.Y(n_2934)
);

OAI22xp5_ASAP7_75t_L g2935 ( 
.A1(n_2494),
.A2(n_2545),
.B1(n_2570),
.B2(n_2684),
.Y(n_2935)
);

OA21x2_ASAP7_75t_L g2936 ( 
.A1(n_2744),
.A2(n_76),
.B(n_78),
.Y(n_2936)
);

OAI21x1_ASAP7_75t_L g2937 ( 
.A1(n_2493),
.A2(n_402),
.B(n_399),
.Y(n_2937)
);

OAI21x1_ASAP7_75t_SL g2938 ( 
.A1(n_2670),
.A2(n_76),
.B(n_78),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2567),
.Y(n_2939)
);

AO31x2_ASAP7_75t_L g2940 ( 
.A1(n_2697),
.A2(n_81),
.A3(n_79),
.B(n_80),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2567),
.Y(n_2941)
);

OAI21x1_ASAP7_75t_L g2942 ( 
.A1(n_2526),
.A2(n_407),
.B(n_406),
.Y(n_2942)
);

OAI21x1_ASAP7_75t_L g2943 ( 
.A1(n_2635),
.A2(n_409),
.B(n_408),
.Y(n_2943)
);

OAI22xp33_ASAP7_75t_L g2944 ( 
.A1(n_2545),
.A2(n_83),
.B1(n_80),
.B2(n_82),
.Y(n_2944)
);

HB1xp67_ASAP7_75t_L g2945 ( 
.A(n_2535),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_2714),
.Y(n_2946)
);

AO21x2_ASAP7_75t_L g2947 ( 
.A1(n_2632),
.A2(n_83),
.B(n_84),
.Y(n_2947)
);

AOI21xp5_ASAP7_75t_L g2948 ( 
.A1(n_2679),
.A2(n_976),
.B(n_972),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2600),
.B(n_84),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2670),
.Y(n_2950)
);

OAI21x1_ASAP7_75t_L g2951 ( 
.A1(n_2635),
.A2(n_415),
.B(n_410),
.Y(n_2951)
);

O2A1O1Ixp33_ASAP7_75t_L g2952 ( 
.A1(n_2702),
.A2(n_88),
.B(n_85),
.C(n_87),
.Y(n_2952)
);

OAI21x1_ASAP7_75t_L g2953 ( 
.A1(n_2571),
.A2(n_421),
.B(n_418),
.Y(n_2953)
);

CKINVDCx11_ASAP7_75t_R g2954 ( 
.A(n_2633),
.Y(n_2954)
);

OAI21x1_ASAP7_75t_L g2955 ( 
.A1(n_2571),
.A2(n_423),
.B(n_422),
.Y(n_2955)
);

OAI21x1_ASAP7_75t_L g2956 ( 
.A1(n_2637),
.A2(n_2705),
.B(n_2691),
.Y(n_2956)
);

AOI22x1_ASAP7_75t_L g2957 ( 
.A1(n_2654),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_2957)
);

NOR2x1_ASAP7_75t_SL g2958 ( 
.A(n_2731),
.B(n_976),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2660),
.B(n_89),
.Y(n_2959)
);

AND2x4_ASAP7_75t_L g2960 ( 
.A(n_2714),
.B(n_430),
.Y(n_2960)
);

OA21x2_ASAP7_75t_L g2961 ( 
.A1(n_2632),
.A2(n_91),
.B(n_92),
.Y(n_2961)
);

AND2x4_ASAP7_75t_L g2962 ( 
.A(n_2714),
.B(n_431),
.Y(n_2962)
);

OAI21xp5_ASAP7_75t_L g2963 ( 
.A1(n_2636),
.A2(n_440),
.B(n_438),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2714),
.Y(n_2964)
);

BUFx6f_ASAP7_75t_L g2965 ( 
.A(n_2489),
.Y(n_2965)
);

OAI21x1_ASAP7_75t_L g2966 ( 
.A1(n_2637),
.A2(n_442),
.B(n_441),
.Y(n_2966)
);

AND2x4_ASAP7_75t_L g2967 ( 
.A(n_2681),
.B(n_2663),
.Y(n_2967)
);

HB1xp67_ASAP7_75t_L g2968 ( 
.A(n_2748),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2599),
.B(n_91),
.Y(n_2969)
);

INVx1_ASAP7_75t_SL g2970 ( 
.A(n_2517),
.Y(n_2970)
);

INVx2_ASAP7_75t_SL g2971 ( 
.A(n_2593),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2665),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2696),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2763),
.Y(n_2974)
);

BUFx2_ASAP7_75t_L g2975 ( 
.A(n_2967),
.Y(n_2975)
);

INVxp33_ASAP7_75t_L g2976 ( 
.A(n_2954),
.Y(n_2976)
);

AND2x2_ASAP7_75t_L g2977 ( 
.A(n_2801),
.B(n_2604),
.Y(n_2977)
);

AOI22xp33_ASAP7_75t_L g2978 ( 
.A1(n_2847),
.A2(n_2747),
.B1(n_2738),
.B2(n_2570),
.Y(n_2978)
);

BUFx6f_ASAP7_75t_L g2979 ( 
.A(n_2917),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2763),
.Y(n_2980)
);

AND2x4_ASAP7_75t_L g2981 ( 
.A(n_2967),
.B(n_2550),
.Y(n_2981)
);

AND2x2_ASAP7_75t_L g2982 ( 
.A(n_2921),
.B(n_2514),
.Y(n_2982)
);

NOR3xp33_ASAP7_75t_SL g2983 ( 
.A(n_2915),
.B(n_2506),
.C(n_2696),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2753),
.B(n_2864),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2773),
.Y(n_2985)
);

AND2x2_ASAP7_75t_L g2986 ( 
.A(n_2808),
.B(n_2597),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2773),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2750),
.Y(n_2988)
);

INVx2_ASAP7_75t_SL g2989 ( 
.A(n_2760),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2930),
.B(n_2652),
.Y(n_2990)
);

OAI21x1_ASAP7_75t_L g2991 ( 
.A1(n_2852),
.A2(n_2705),
.B(n_2691),
.Y(n_2991)
);

NAND3xp33_ASAP7_75t_L g2992 ( 
.A(n_2847),
.B(n_2534),
.C(n_2499),
.Y(n_2992)
);

NAND2xp33_ASAP7_75t_R g2993 ( 
.A(n_2915),
.B(n_2699),
.Y(n_2993)
);

AOI21xp5_ASAP7_75t_L g2994 ( 
.A1(n_2754),
.A2(n_2648),
.B(n_2570),
.Y(n_2994)
);

NAND2xp33_ASAP7_75t_R g2995 ( 
.A(n_2828),
.B(n_2692),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2808),
.B(n_2504),
.Y(n_2996)
);

OAI22xp5_ASAP7_75t_L g2997 ( 
.A1(n_2766),
.A2(n_2570),
.B1(n_2747),
.B2(n_2708),
.Y(n_2997)
);

NOR2xp33_ASAP7_75t_L g2998 ( 
.A(n_2842),
.B(n_2540),
.Y(n_2998)
);

AND2x4_ASAP7_75t_L g2999 ( 
.A(n_2967),
.B(n_2586),
.Y(n_2999)
);

INVx1_ASAP7_75t_SL g3000 ( 
.A(n_2778),
.Y(n_3000)
);

AOI22xp33_ASAP7_75t_L g3001 ( 
.A1(n_2847),
.A2(n_2908),
.B1(n_2766),
.B2(n_2963),
.Y(n_3001)
);

OAI22xp5_ASAP7_75t_L g3002 ( 
.A1(n_2866),
.A2(n_2530),
.B1(n_2556),
.B2(n_2552),
.Y(n_3002)
);

AOI221xp5_ASAP7_75t_L g3003 ( 
.A1(n_2878),
.A2(n_2499),
.B1(n_2534),
.B2(n_2548),
.C(n_2601),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2755),
.Y(n_3004)
);

NAND2x1p5_ASAP7_75t_L g3005 ( 
.A(n_2874),
.B(n_2520),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2756),
.Y(n_3006)
);

INVx2_ASAP7_75t_SL g3007 ( 
.A(n_2877),
.Y(n_3007)
);

INVx1_ASAP7_75t_SL g3008 ( 
.A(n_2832),
.Y(n_3008)
);

CKINVDCx5p33_ASAP7_75t_R g3009 ( 
.A(n_2828),
.Y(n_3009)
);

INVx2_ASAP7_75t_SL g3010 ( 
.A(n_2877),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2771),
.Y(n_3011)
);

INVx3_ASAP7_75t_L g3012 ( 
.A(n_2887),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2933),
.B(n_2652),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2782),
.Y(n_3014)
);

INVx4_ASAP7_75t_L g3015 ( 
.A(n_2887),
.Y(n_3015)
);

INVx4_ASAP7_75t_L g3016 ( 
.A(n_2954),
.Y(n_3016)
);

CKINVDCx5p33_ASAP7_75t_R g3017 ( 
.A(n_2910),
.Y(n_3017)
);

HB1xp67_ASAP7_75t_L g3018 ( 
.A(n_2968),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2861),
.Y(n_3019)
);

AOI22xp33_ASAP7_75t_L g3020 ( 
.A1(n_2908),
.A2(n_2738),
.B1(n_2661),
.B2(n_2730),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_2914),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2939),
.B(n_2611),
.Y(n_3022)
);

BUFx6f_ASAP7_75t_L g3023 ( 
.A(n_2917),
.Y(n_3023)
);

AOI22xp5_ASAP7_75t_L g3024 ( 
.A1(n_2908),
.A2(n_2638),
.B1(n_2647),
.B2(n_2485),
.Y(n_3024)
);

AOI21xp33_ASAP7_75t_L g3025 ( 
.A1(n_2878),
.A2(n_2952),
.B(n_2926),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2941),
.B(n_2611),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2783),
.Y(n_3027)
);

INVx6_ASAP7_75t_L g3028 ( 
.A(n_2917),
.Y(n_3028)
);

AND2x4_ASAP7_75t_L g3029 ( 
.A(n_2913),
.B(n_2829),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2790),
.B(n_2552),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_2914),
.Y(n_3031)
);

NAND2x1p5_ASAP7_75t_L g3032 ( 
.A(n_2874),
.B(n_2730),
.Y(n_3032)
);

OAI22xp33_ASAP7_75t_L g3033 ( 
.A1(n_2799),
.A2(n_2556),
.B1(n_2638),
.B2(n_2728),
.Y(n_3033)
);

CKINVDCx5p33_ASAP7_75t_R g3034 ( 
.A(n_2910),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2927),
.Y(n_3035)
);

BUFx6f_ASAP7_75t_L g3036 ( 
.A(n_2917),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2927),
.Y(n_3037)
);

AOI22xp33_ASAP7_75t_L g3038 ( 
.A1(n_2837),
.A2(n_2796),
.B1(n_2890),
.B2(n_2802),
.Y(n_3038)
);

OAI22xp5_ASAP7_75t_L g3039 ( 
.A1(n_2866),
.A2(n_2743),
.B1(n_2690),
.B2(n_2698),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2819),
.B(n_2821),
.Y(n_3040)
);

OAI22xp33_ASAP7_75t_L g3041 ( 
.A1(n_2769),
.A2(n_2797),
.B1(n_2879),
.B2(n_2944),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2968),
.Y(n_3042)
);

OAI221xp5_ASAP7_75t_L g3043 ( 
.A1(n_2905),
.A2(n_2656),
.B1(n_2578),
.B2(n_2743),
.C(n_2565),
.Y(n_3043)
);

AOI21xp33_ASAP7_75t_L g3044 ( 
.A1(n_2924),
.A2(n_2796),
.B(n_2961),
.Y(n_3044)
);

INVx3_ASAP7_75t_L g3045 ( 
.A(n_2946),
.Y(n_3045)
);

AOI22xp33_ASAP7_75t_L g3046 ( 
.A1(n_2837),
.A2(n_2686),
.B1(n_2666),
.B2(n_2680),
.Y(n_3046)
);

AND2x4_ASAP7_75t_L g3047 ( 
.A(n_2913),
.B(n_2829),
.Y(n_3047)
);

OR2x2_ASAP7_75t_L g3048 ( 
.A(n_2898),
.B(n_2619),
.Y(n_3048)
);

OAI22xp33_ASAP7_75t_L g3049 ( 
.A1(n_2944),
.A2(n_2666),
.B1(n_2505),
.B2(n_2643),
.Y(n_3049)
);

INVx1_ASAP7_75t_SL g3050 ( 
.A(n_2761),
.Y(n_3050)
);

AOI22xp33_ASAP7_75t_L g3051 ( 
.A1(n_2802),
.A2(n_2666),
.B1(n_2649),
.B2(n_2653),
.Y(n_3051)
);

AOI22xp33_ASAP7_75t_L g3052 ( 
.A1(n_2901),
.A2(n_2649),
.B1(n_2653),
.B2(n_2682),
.Y(n_3052)
);

BUFx2_ASAP7_75t_L g3053 ( 
.A(n_2777),
.Y(n_3053)
);

CKINVDCx5p33_ASAP7_75t_R g3054 ( 
.A(n_2765),
.Y(n_3054)
);

OAI21x1_ASAP7_75t_L g3055 ( 
.A1(n_2929),
.A2(n_2727),
.B(n_2729),
.Y(n_3055)
);

INVx11_ASAP7_75t_L g3056 ( 
.A(n_2834),
.Y(n_3056)
);

BUFx2_ASAP7_75t_L g3057 ( 
.A(n_2777),
.Y(n_3057)
);

OAI221xp5_ASAP7_75t_L g3058 ( 
.A1(n_2905),
.A2(n_2643),
.B1(n_2619),
.B2(n_2672),
.C(n_2726),
.Y(n_3058)
);

HB1xp67_ASAP7_75t_L g3059 ( 
.A(n_2776),
.Y(n_3059)
);

CKINVDCx14_ASAP7_75t_R g3060 ( 
.A(n_2803),
.Y(n_3060)
);

INVx2_ASAP7_75t_L g3061 ( 
.A(n_2830),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2950),
.B(n_2715),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2922),
.Y(n_3063)
);

BUFx6f_ASAP7_75t_L g3064 ( 
.A(n_2965),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2973),
.B(n_2510),
.Y(n_3065)
);

AOI221xp5_ASAP7_75t_L g3066 ( 
.A1(n_2798),
.A2(n_2682),
.B1(n_2710),
.B2(n_2503),
.C(n_2566),
.Y(n_3066)
);

CKINVDCx16_ASAP7_75t_R g3067 ( 
.A(n_2768),
.Y(n_3067)
);

NAND3xp33_ASAP7_75t_SL g3068 ( 
.A(n_2762),
.B(n_2505),
.C(n_2648),
.Y(n_3068)
);

INVx2_ASAP7_75t_SL g3069 ( 
.A(n_2904),
.Y(n_3069)
);

NAND2x1_ASAP7_75t_L g3070 ( 
.A(n_2906),
.B(n_2835),
.Y(n_3070)
);

BUFx3_ASAP7_75t_L g3071 ( 
.A(n_2862),
.Y(n_3071)
);

A2O1A1Ixp33_ASAP7_75t_L g3072 ( 
.A1(n_2883),
.A2(n_2627),
.B(n_2704),
.C(n_2710),
.Y(n_3072)
);

OAI22xp33_ASAP7_75t_L g3073 ( 
.A1(n_2770),
.A2(n_2503),
.B1(n_2537),
.B2(n_2481),
.Y(n_3073)
);

OAI21xp5_ASAP7_75t_L g3074 ( 
.A1(n_2883),
.A2(n_2754),
.B(n_2798),
.Y(n_3074)
);

AOI22xp33_ASAP7_75t_L g3075 ( 
.A1(n_2901),
.A2(n_2704),
.B1(n_2627),
.B2(n_2693),
.Y(n_3075)
);

AOI22xp33_ASAP7_75t_L g3076 ( 
.A1(n_2759),
.A2(n_2693),
.B1(n_2486),
.B2(n_2646),
.Y(n_3076)
);

BUFx12f_ASAP7_75t_L g3077 ( 
.A(n_2853),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2972),
.Y(n_3078)
);

HB1xp67_ASAP7_75t_L g3079 ( 
.A(n_2787),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_2935),
.B(n_2689),
.Y(n_3080)
);

CKINVDCx20_ASAP7_75t_R g3081 ( 
.A(n_2793),
.Y(n_3081)
);

AOI22xp33_ASAP7_75t_L g3082 ( 
.A1(n_2759),
.A2(n_2646),
.B1(n_2596),
.B2(n_2537),
.Y(n_3082)
);

OR2x2_ASAP7_75t_L g3083 ( 
.A(n_2898),
.B(n_2608),
.Y(n_3083)
);

AOI22xp33_ASAP7_75t_L g3084 ( 
.A1(n_2759),
.A2(n_2596),
.B1(n_2566),
.B2(n_2481),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2972),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2923),
.Y(n_3086)
);

AOI22xp33_ASAP7_75t_L g3087 ( 
.A1(n_2779),
.A2(n_2669),
.B1(n_2644),
.B2(n_2720),
.Y(n_3087)
);

AND2x4_ASAP7_75t_L g3088 ( 
.A(n_2835),
.B(n_2594),
.Y(n_3088)
);

INVx2_ASAP7_75t_L g3089 ( 
.A(n_2870),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2898),
.B(n_2510),
.Y(n_3090)
);

BUFx6f_ASAP7_75t_L g3091 ( 
.A(n_2965),
.Y(n_3091)
);

AOI22xp33_ASAP7_75t_SL g3092 ( 
.A1(n_2957),
.A2(n_2510),
.B1(n_2720),
.B2(n_2688),
.Y(n_3092)
);

INVx2_ASAP7_75t_L g3093 ( 
.A(n_2881),
.Y(n_3093)
);

AND2x6_ASAP7_75t_L g3094 ( 
.A(n_2960),
.B(n_2603),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2925),
.B(n_2888),
.Y(n_3095)
);

AOI22xp33_ASAP7_75t_SL g3096 ( 
.A1(n_2767),
.A2(n_2510),
.B1(n_2688),
.B2(n_2724),
.Y(n_3096)
);

OR2x2_ASAP7_75t_L g3097 ( 
.A(n_2787),
.B(n_2668),
.Y(n_3097)
);

A2O1A1Ixp33_ASAP7_75t_L g3098 ( 
.A1(n_2764),
.A2(n_2603),
.B(n_2648),
.C(n_2547),
.Y(n_3098)
);

AOI22xp33_ASAP7_75t_L g3099 ( 
.A1(n_2912),
.A2(n_2609),
.B1(n_2642),
.B2(n_2640),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2848),
.Y(n_3100)
);

BUFx3_ASAP7_75t_L g3101 ( 
.A(n_2904),
.Y(n_3101)
);

AOI22xp5_ASAP7_75t_L g3102 ( 
.A1(n_2902),
.A2(n_2588),
.B1(n_2547),
.B2(n_2513),
.Y(n_3102)
);

BUFx10_ASAP7_75t_L g3103 ( 
.A(n_2960),
.Y(n_3103)
);

INVxp33_ASAP7_75t_SL g3104 ( 
.A(n_2873),
.Y(n_3104)
);

INVx6_ASAP7_75t_L g3105 ( 
.A(n_2965),
.Y(n_3105)
);

OAI222xp33_ASAP7_75t_L g3106 ( 
.A1(n_2857),
.A2(n_2668),
.B1(n_2650),
.B2(n_2727),
.C1(n_2674),
.C2(n_2676),
.Y(n_3106)
);

AOI21x1_ASAP7_75t_L g3107 ( 
.A1(n_2916),
.A2(n_2729),
.B(n_2588),
.Y(n_3107)
);

BUFx2_ASAP7_75t_L g3108 ( 
.A(n_2791),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2892),
.B(n_2721),
.Y(n_3109)
);

NAND2xp33_ASAP7_75t_R g3110 ( 
.A(n_2791),
.B(n_2916),
.Y(n_3110)
);

AO31x2_ASAP7_75t_L g3111 ( 
.A1(n_2792),
.A2(n_2741),
.A3(n_2674),
.B(n_2689),
.Y(n_3111)
);

CKINVDCx8_ASAP7_75t_R g3112 ( 
.A(n_2965),
.Y(n_3112)
);

INVx4_ASAP7_75t_SL g3113 ( 
.A(n_2940),
.Y(n_3113)
);

INVx1_ASAP7_75t_SL g3114 ( 
.A(n_2845),
.Y(n_3114)
);

NAND2xp33_ASAP7_75t_L g3115 ( 
.A(n_2874),
.B(n_2489),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2838),
.Y(n_3116)
);

OAI22xp5_ASAP7_75t_L g3117 ( 
.A1(n_2912),
.A2(n_2689),
.B1(n_2721),
.B2(n_2569),
.Y(n_3117)
);

INVx4_ASAP7_75t_L g3118 ( 
.A(n_2768),
.Y(n_3118)
);

AOI22xp33_ASAP7_75t_L g3119 ( 
.A1(n_2900),
.A2(n_2721),
.B1(n_2569),
.B2(n_2591),
.Y(n_3119)
);

AOI221xp5_ASAP7_75t_L g3120 ( 
.A1(n_2831),
.A2(n_2631),
.B1(n_2591),
.B2(n_2569),
.C(n_2513),
.Y(n_3120)
);

AND2x4_ASAP7_75t_L g3121 ( 
.A(n_2835),
.B(n_2513),
.Y(n_3121)
);

AND2x2_ASAP7_75t_L g3122 ( 
.A(n_2785),
.B(n_2591),
.Y(n_3122)
);

NOR2xp33_ASAP7_75t_L g3123 ( 
.A(n_2970),
.B(n_2631),
.Y(n_3123)
);

BUFx4_ASAP7_75t_SL g3124 ( 
.A(n_2896),
.Y(n_3124)
);

AND2x6_ASAP7_75t_SL g3125 ( 
.A(n_2863),
.B(n_94),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2841),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2811),
.Y(n_3127)
);

AO21x1_ASAP7_75t_L g3128 ( 
.A1(n_2928),
.A2(n_2899),
.B(n_2827),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2811),
.Y(n_3129)
);

AOI22xp33_ASAP7_75t_L g3130 ( 
.A1(n_2900),
.A2(n_2631),
.B1(n_2741),
.B2(n_2709),
.Y(n_3130)
);

AOI22xp33_ASAP7_75t_L g3131 ( 
.A1(n_2947),
.A2(n_2741),
.B1(n_979),
.B2(n_1004),
.Y(n_3131)
);

AOI22xp33_ASAP7_75t_L g3132 ( 
.A1(n_2947),
.A2(n_2920),
.B1(n_2810),
.B2(n_2859),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2897),
.Y(n_3133)
);

OR2x6_ASAP7_75t_L g3134 ( 
.A(n_2780),
.B(n_976),
.Y(n_3134)
);

BUFx4f_ASAP7_75t_SL g3135 ( 
.A(n_2918),
.Y(n_3135)
);

OR2x2_ASAP7_75t_L g3136 ( 
.A(n_2795),
.B(n_94),
.Y(n_3136)
);

NOR2x1p5_ASAP7_75t_L g3137 ( 
.A(n_2969),
.B(n_1048),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2894),
.Y(n_3138)
);

CKINVDCx20_ASAP7_75t_R g3139 ( 
.A(n_2757),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2895),
.Y(n_3140)
);

AND2x2_ASAP7_75t_L g3141 ( 
.A(n_2805),
.B(n_95),
.Y(n_3141)
);

CKINVDCx5p33_ASAP7_75t_R g3142 ( 
.A(n_2971),
.Y(n_3142)
);

AOI21xp5_ASAP7_75t_L g3143 ( 
.A1(n_2826),
.A2(n_979),
.B(n_976),
.Y(n_3143)
);

AO31x2_ASAP7_75t_L g3144 ( 
.A1(n_2792),
.A2(n_98),
.A3(n_96),
.B(n_97),
.Y(n_3144)
);

INVx2_ASAP7_75t_SL g3145 ( 
.A(n_2946),
.Y(n_3145)
);

OR2x2_ASAP7_75t_L g3146 ( 
.A(n_2818),
.B(n_2775),
.Y(n_3146)
);

AOI22xp33_ASAP7_75t_L g3147 ( 
.A1(n_2859),
.A2(n_1004),
.B1(n_1005),
.B2(n_979),
.Y(n_3147)
);

AOI21xp5_ASAP7_75t_L g3148 ( 
.A1(n_2826),
.A2(n_1004),
.B(n_979),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_2903),
.Y(n_3149)
);

CKINVDCx6p67_ASAP7_75t_R g3150 ( 
.A(n_2949),
.Y(n_3150)
);

BUFx3_ASAP7_75t_L g3151 ( 
.A(n_2859),
.Y(n_3151)
);

NOR3xp33_ASAP7_75t_SL g3152 ( 
.A(n_2849),
.B(n_96),
.C(n_97),
.Y(n_3152)
);

OAI22xp33_ASAP7_75t_L g3153 ( 
.A1(n_2961),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_3153)
);

AOI221xp5_ASAP7_75t_L g3154 ( 
.A1(n_2938),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.C(n_102),
.Y(n_3154)
);

AOI221xp5_ASAP7_75t_L g3155 ( 
.A1(n_2945),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.C(n_108),
.Y(n_3155)
);

OAI221xp5_ASAP7_75t_L g3156 ( 
.A1(n_2851),
.A2(n_104),
.B1(n_106),
.B2(n_108),
.C(n_109),
.Y(n_3156)
);

OAI22xp33_ASAP7_75t_L g3157 ( 
.A1(n_2961),
.A2(n_2874),
.B1(n_2916),
.B2(n_2907),
.Y(n_3157)
);

BUFx2_ASAP7_75t_L g3158 ( 
.A(n_2964),
.Y(n_3158)
);

AND2x4_ASAP7_75t_L g3159 ( 
.A(n_2964),
.B(n_110),
.Y(n_3159)
);

AND2x4_ASAP7_75t_L g3160 ( 
.A(n_2780),
.B(n_112),
.Y(n_3160)
);

OAI22xp33_ASAP7_75t_L g3161 ( 
.A1(n_2907),
.A2(n_116),
.B1(n_113),
.B2(n_114),
.Y(n_3161)
);

BUFx6f_ASAP7_75t_L g3162 ( 
.A(n_2960),
.Y(n_3162)
);

AOI22xp33_ASAP7_75t_L g3163 ( 
.A1(n_2855),
.A2(n_1005),
.B1(n_1007),
.B2(n_1004),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2867),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2867),
.Y(n_3165)
);

BUFx12f_ASAP7_75t_L g3166 ( 
.A(n_2962),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2800),
.Y(n_3167)
);

OAI21x1_ASAP7_75t_L g3168 ( 
.A1(n_2991),
.A2(n_2816),
.B(n_2956),
.Y(n_3168)
);

INVx2_ASAP7_75t_L g3169 ( 
.A(n_3165),
.Y(n_3169)
);

AND2x2_ASAP7_75t_L g3170 ( 
.A(n_2975),
.B(n_2945),
.Y(n_3170)
);

AND2x2_ASAP7_75t_L g3171 ( 
.A(n_3059),
.B(n_2780),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_3167),
.Y(n_3172)
);

AND2x4_ASAP7_75t_L g3173 ( 
.A(n_3113),
.B(n_2934),
.Y(n_3173)
);

INVx3_ASAP7_75t_L g3174 ( 
.A(n_3070),
.Y(n_3174)
);

HB1xp67_ASAP7_75t_L g3175 ( 
.A(n_3079),
.Y(n_3175)
);

OA21x2_ASAP7_75t_L g3176 ( 
.A1(n_3044),
.A2(n_2816),
.B(n_2817),
.Y(n_3176)
);

CKINVDCx5p33_ASAP7_75t_R g3177 ( 
.A(n_3054),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_3127),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_3164),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_3100),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_3129),
.Y(n_3181)
);

HB1xp67_ASAP7_75t_L g3182 ( 
.A(n_3018),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_3019),
.Y(n_3183)
);

INVx5_ASAP7_75t_SL g3184 ( 
.A(n_3134),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_3050),
.B(n_2758),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2974),
.Y(n_3186)
);

BUFx6f_ASAP7_75t_L g3187 ( 
.A(n_3160),
.Y(n_3187)
);

BUFx12f_ASAP7_75t_L g3188 ( 
.A(n_3016),
.Y(n_3188)
);

INVx2_ASAP7_75t_L g3189 ( 
.A(n_3083),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2980),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2985),
.Y(n_3191)
);

BUFx6f_ASAP7_75t_L g3192 ( 
.A(n_3160),
.Y(n_3192)
);

AO21x2_ASAP7_75t_L g3193 ( 
.A1(n_3044),
.A2(n_2924),
.B(n_2794),
.Y(n_3193)
);

AND2x2_ASAP7_75t_L g3194 ( 
.A(n_3008),
.B(n_2906),
.Y(n_3194)
);

BUFx2_ASAP7_75t_L g3195 ( 
.A(n_3158),
.Y(n_3195)
);

AND2x2_ASAP7_75t_L g3196 ( 
.A(n_3008),
.B(n_2906),
.Y(n_3196)
);

AOI22xp33_ASAP7_75t_L g3197 ( 
.A1(n_2992),
.A2(n_2855),
.B1(n_2907),
.B2(n_2815),
.Y(n_3197)
);

INVxp67_ASAP7_75t_SL g3198 ( 
.A(n_3090),
.Y(n_3198)
);

INVx3_ASAP7_75t_L g3199 ( 
.A(n_3121),
.Y(n_3199)
);

HB1xp67_ASAP7_75t_L g3200 ( 
.A(n_3114),
.Y(n_3200)
);

INVx3_ASAP7_75t_L g3201 ( 
.A(n_3121),
.Y(n_3201)
);

INVx2_ASAP7_75t_SL g3202 ( 
.A(n_3045),
.Y(n_3202)
);

AO21x2_ASAP7_75t_L g3203 ( 
.A1(n_3157),
.A2(n_2794),
.B(n_2817),
.Y(n_3203)
);

HB1xp67_ASAP7_75t_L g3204 ( 
.A(n_3114),
.Y(n_3204)
);

NOR2xp33_ASAP7_75t_L g3205 ( 
.A(n_3016),
.B(n_2932),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2987),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_3035),
.Y(n_3207)
);

OAI21x1_ASAP7_75t_L g3208 ( 
.A1(n_3055),
.A2(n_2752),
.B(n_2929),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2988),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3014),
.Y(n_3210)
);

AND2x4_ASAP7_75t_L g3211 ( 
.A(n_3113),
.B(n_2934),
.Y(n_3211)
);

OR2x2_ASAP7_75t_L g3212 ( 
.A(n_3050),
.B(n_2800),
.Y(n_3212)
);

NOR2xp33_ASAP7_75t_L g3213 ( 
.A(n_2976),
.B(n_2959),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3042),
.Y(n_3214)
);

NAND2x1_ASAP7_75t_L g3215 ( 
.A(n_3134),
.B(n_2936),
.Y(n_3215)
);

INVx2_ASAP7_75t_L g3216 ( 
.A(n_3021),
.Y(n_3216)
);

AOI21x1_ASAP7_75t_L g3217 ( 
.A1(n_3062),
.A2(n_2936),
.B(n_2911),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_3031),
.Y(n_3218)
);

INVx2_ASAP7_75t_L g3219 ( 
.A(n_3037),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_3004),
.Y(n_3220)
);

INVx2_ASAP7_75t_L g3221 ( 
.A(n_3006),
.Y(n_3221)
);

BUFx2_ASAP7_75t_SL g3222 ( 
.A(n_3118),
.Y(n_3222)
);

INVx2_ASAP7_75t_L g3223 ( 
.A(n_3078),
.Y(n_3223)
);

AND2x4_ASAP7_75t_L g3224 ( 
.A(n_3113),
.B(n_2822),
.Y(n_3224)
);

HB1xp67_ASAP7_75t_L g3225 ( 
.A(n_3097),
.Y(n_3225)
);

AO21x2_ASAP7_75t_L g3226 ( 
.A1(n_2994),
.A2(n_2822),
.B(n_2909),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3011),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_3085),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_3063),
.Y(n_3229)
);

OR2x2_ASAP7_75t_L g3230 ( 
.A(n_3146),
.B(n_2911),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_3086),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3040),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3040),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_3144),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3116),
.Y(n_3235)
);

INVx4_ASAP7_75t_L g3236 ( 
.A(n_3118),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_3144),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_3126),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_3144),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3133),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_3149),
.Y(n_3241)
);

AND2x2_ASAP7_75t_L g3242 ( 
.A(n_3045),
.B(n_3053),
.Y(n_3242)
);

HB1xp67_ASAP7_75t_L g3243 ( 
.A(n_3110),
.Y(n_3243)
);

AND2x2_ASAP7_75t_L g3244 ( 
.A(n_3057),
.B(n_2825),
.Y(n_3244)
);

AND2x2_ASAP7_75t_L g3245 ( 
.A(n_3108),
.B(n_2986),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3095),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_3048),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_3095),
.Y(n_3248)
);

AO21x2_ASAP7_75t_L g3249 ( 
.A1(n_3062),
.A2(n_2836),
.B(n_2825),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3138),
.Y(n_3250)
);

INVx2_ASAP7_75t_L g3251 ( 
.A(n_3140),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_3027),
.Y(n_3252)
);

HB1xp67_ASAP7_75t_L g3253 ( 
.A(n_3030),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_3107),
.Y(n_3254)
);

OAI21x1_ASAP7_75t_L g3255 ( 
.A1(n_3143),
.A2(n_2751),
.B(n_2884),
.Y(n_3255)
);

INVx3_ASAP7_75t_L g3256 ( 
.A(n_3029),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_3061),
.Y(n_3257)
);

OAI21x1_ASAP7_75t_L g3258 ( 
.A1(n_3148),
.A2(n_2781),
.B(n_2772),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3089),
.Y(n_3259)
);

HB1xp67_ASAP7_75t_L g3260 ( 
.A(n_3030),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_3093),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_3145),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_3109),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_3109),
.Y(n_3264)
);

BUFx2_ASAP7_75t_L g3265 ( 
.A(n_3088),
.Y(n_3265)
);

AOI21xp5_ASAP7_75t_SL g3266 ( 
.A1(n_3074),
.A2(n_2936),
.B(n_2885),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_3038),
.B(n_2788),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2990),
.B(n_3013),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3090),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3128),
.Y(n_3270)
);

INVx5_ASAP7_75t_L g3271 ( 
.A(n_3134),
.Y(n_3271)
);

BUFx3_ASAP7_75t_L g3272 ( 
.A(n_3101),
.Y(n_3272)
);

AND2x2_ASAP7_75t_L g3273 ( 
.A(n_3122),
.B(n_2836),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3065),
.Y(n_3274)
);

INVxp33_ASAP7_75t_L g3275 ( 
.A(n_2998),
.Y(n_3275)
);

OR2x6_ASAP7_75t_L g3276 ( 
.A(n_3074),
.B(n_2855),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_3029),
.B(n_2854),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3065),
.Y(n_3278)
);

HB1xp67_ASAP7_75t_L g3279 ( 
.A(n_3000),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_3111),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2990),
.B(n_2789),
.Y(n_3281)
);

HB1xp67_ASAP7_75t_L g3282 ( 
.A(n_3000),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3047),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_3047),
.Y(n_3284)
);

AND2x2_ASAP7_75t_L g3285 ( 
.A(n_2996),
.B(n_2854),
.Y(n_3285)
);

BUFx2_ASAP7_75t_L g3286 ( 
.A(n_3088),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_3111),
.Y(n_3287)
);

BUFx3_ASAP7_75t_L g3288 ( 
.A(n_3012),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3013),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_3111),
.Y(n_3290)
);

AND2x2_ASAP7_75t_L g3291 ( 
.A(n_2984),
.B(n_2774),
.Y(n_3291)
);

INVx3_ASAP7_75t_L g3292 ( 
.A(n_3005),
.Y(n_3292)
);

HB1xp67_ASAP7_75t_L g3293 ( 
.A(n_2977),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_3022),
.Y(n_3294)
);

NAND2x1p5_ASAP7_75t_L g3295 ( 
.A(n_3080),
.B(n_2885),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3022),
.Y(n_3296)
);

AND2x2_ASAP7_75t_L g3297 ( 
.A(n_2982),
.B(n_2774),
.Y(n_3297)
);

INVx3_ASAP7_75t_L g3298 ( 
.A(n_3005),
.Y(n_3298)
);

AND2x2_ASAP7_75t_L g3299 ( 
.A(n_2981),
.B(n_2774),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_2981),
.B(n_2774),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3026),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3026),
.Y(n_3302)
);

BUFx6f_ASAP7_75t_L g3303 ( 
.A(n_2979),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_2979),
.Y(n_3304)
);

INVx1_ASAP7_75t_SL g3305 ( 
.A(n_3135),
.Y(n_3305)
);

AO21x2_ASAP7_75t_L g3306 ( 
.A1(n_3153),
.A2(n_2886),
.B(n_2844),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_2979),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_3136),
.Y(n_3308)
);

AO21x2_ASAP7_75t_L g3309 ( 
.A1(n_3161),
.A2(n_2886),
.B(n_2844),
.Y(n_3309)
);

AND2x2_ASAP7_75t_L g3310 ( 
.A(n_2999),
.B(n_3007),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_2999),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_3023),
.Y(n_3312)
);

HB1xp67_ASAP7_75t_L g3313 ( 
.A(n_3010),
.Y(n_3313)
);

AND2x2_ASAP7_75t_L g3314 ( 
.A(n_3069),
.B(n_2774),
.Y(n_3314)
);

BUFx6f_ASAP7_75t_L g3315 ( 
.A(n_3023),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3033),
.B(n_2813),
.Y(n_3316)
);

OA21x2_ASAP7_75t_L g3317 ( 
.A1(n_3098),
.A2(n_2781),
.B(n_2806),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3023),
.Y(n_3318)
);

HB1xp67_ASAP7_75t_L g3319 ( 
.A(n_3124),
.Y(n_3319)
);

BUFx2_ASAP7_75t_L g3320 ( 
.A(n_3012),
.Y(n_3320)
);

INVx2_ASAP7_75t_L g3321 ( 
.A(n_3036),
.Y(n_3321)
);

NOR2xp33_ASAP7_75t_L g3322 ( 
.A(n_3015),
.B(n_2889),
.Y(n_3322)
);

OR2x2_ASAP7_75t_L g3323 ( 
.A(n_3002),
.B(n_2823),
.Y(n_3323)
);

INVx3_ASAP7_75t_L g3324 ( 
.A(n_3036),
.Y(n_3324)
);

HB1xp67_ASAP7_75t_L g3325 ( 
.A(n_3036),
.Y(n_3325)
);

AND2x2_ASAP7_75t_L g3326 ( 
.A(n_2989),
.B(n_2774),
.Y(n_3326)
);

AND2x2_ASAP7_75t_L g3327 ( 
.A(n_3311),
.B(n_3067),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_3256),
.Y(n_3328)
);

AOI22xp33_ASAP7_75t_L g3329 ( 
.A1(n_3267),
.A2(n_2992),
.B1(n_3001),
.B2(n_3041),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_3180),
.Y(n_3330)
);

NAND3xp33_ASAP7_75t_SL g3331 ( 
.A(n_3243),
.B(n_3066),
.C(n_3156),
.Y(n_3331)
);

OA21x2_ASAP7_75t_L g3332 ( 
.A1(n_3270),
.A2(n_3025),
.B(n_3119),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3256),
.Y(n_3333)
);

AOI22xp33_ASAP7_75t_L g3334 ( 
.A1(n_3197),
.A2(n_3003),
.B1(n_3025),
.B2(n_3039),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3180),
.Y(n_3335)
);

OAI22xp5_ASAP7_75t_L g3336 ( 
.A1(n_3316),
.A2(n_2978),
.B1(n_3152),
.B2(n_3096),
.Y(n_3336)
);

INVx2_ASAP7_75t_L g3337 ( 
.A(n_3256),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_3180),
.Y(n_3338)
);

A2O1A1Ixp33_ASAP7_75t_L g3339 ( 
.A1(n_3205),
.A2(n_3154),
.B(n_2997),
.C(n_2983),
.Y(n_3339)
);

OAI21x1_ASAP7_75t_L g3340 ( 
.A1(n_3215),
.A2(n_3117),
.B(n_3032),
.Y(n_3340)
);

CKINVDCx12_ASAP7_75t_R g3341 ( 
.A(n_3276),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3251),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_L g3343 ( 
.A(n_3289),
.B(n_3002),
.Y(n_3343)
);

OAI22xp5_ASAP7_75t_L g3344 ( 
.A1(n_3276),
.A2(n_3039),
.B1(n_3020),
.B2(n_3092),
.Y(n_3344)
);

AOI22xp33_ASAP7_75t_L g3345 ( 
.A1(n_3270),
.A2(n_2997),
.B1(n_3155),
.B2(n_3043),
.Y(n_3345)
);

OAI221xp5_ASAP7_75t_L g3346 ( 
.A1(n_3268),
.A2(n_2995),
.B1(n_2993),
.B2(n_3132),
.C(n_3120),
.Y(n_3346)
);

AOI22xp33_ASAP7_75t_L g3347 ( 
.A1(n_3295),
.A2(n_3058),
.B1(n_3068),
.B2(n_3049),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_3256),
.Y(n_3348)
);

OAI211xp5_ASAP7_75t_L g3349 ( 
.A1(n_3266),
.A2(n_3072),
.B(n_3024),
.C(n_3058),
.Y(n_3349)
);

OAI21xp33_ASAP7_75t_L g3350 ( 
.A1(n_3198),
.A2(n_3130),
.B(n_3117),
.Y(n_3350)
);

AO21x2_ASAP7_75t_L g3351 ( 
.A1(n_3254),
.A2(n_3073),
.B(n_3141),
.Y(n_3351)
);

AND2x2_ASAP7_75t_L g3352 ( 
.A(n_3311),
.B(n_3245),
.Y(n_3352)
);

AOI21xp33_ASAP7_75t_L g3353 ( 
.A1(n_3275),
.A2(n_3046),
.B(n_3087),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3251),
.Y(n_3354)
);

AOI21xp33_ASAP7_75t_L g3355 ( 
.A1(n_3323),
.A2(n_3082),
.B(n_3099),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3251),
.Y(n_3356)
);

AOI22xp5_ASAP7_75t_SL g3357 ( 
.A1(n_3319),
.A2(n_3104),
.B1(n_3060),
.B2(n_3081),
.Y(n_3357)
);

OAI22xp33_ASAP7_75t_L g3358 ( 
.A1(n_3295),
.A2(n_3150),
.B1(n_3139),
.B2(n_3151),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_3169),
.Y(n_3359)
);

AOI22xp33_ASAP7_75t_SL g3360 ( 
.A1(n_3295),
.A2(n_3192),
.B1(n_3187),
.B2(n_3276),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_3169),
.Y(n_3361)
);

OR2x6_ASAP7_75t_L g3362 ( 
.A(n_3222),
.B(n_3032),
.Y(n_3362)
);

OAI22xp5_ASAP7_75t_L g3363 ( 
.A1(n_3276),
.A2(n_3052),
.B1(n_3051),
.B2(n_3075),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3183),
.Y(n_3364)
);

BUFx6f_ASAP7_75t_SL g3365 ( 
.A(n_3236),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_3245),
.B(n_3015),
.Y(n_3366)
);

AND2x2_ASAP7_75t_L g3367 ( 
.A(n_3310),
.B(n_3123),
.Y(n_3367)
);

OAI21xp33_ASAP7_75t_SL g3368 ( 
.A1(n_3276),
.A2(n_3056),
.B(n_3084),
.Y(n_3368)
);

AOI22xp33_ASAP7_75t_L g3369 ( 
.A1(n_3306),
.A2(n_3137),
.B1(n_2812),
.B2(n_3131),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3183),
.Y(n_3370)
);

AOI22xp33_ASAP7_75t_L g3371 ( 
.A1(n_3306),
.A2(n_2812),
.B1(n_3159),
.B2(n_3077),
.Y(n_3371)
);

AOI221xp5_ASAP7_75t_L g3372 ( 
.A1(n_3269),
.A2(n_3159),
.B1(n_3106),
.B2(n_2840),
.C(n_3142),
.Y(n_3372)
);

AOI22xp5_ASAP7_75t_SL g3373 ( 
.A1(n_3222),
.A2(n_3009),
.B1(n_3034),
.B2(n_3017),
.Y(n_3373)
);

OR2x2_ASAP7_75t_L g3374 ( 
.A(n_3200),
.B(n_3204),
.Y(n_3374)
);

AOI22xp33_ASAP7_75t_L g3375 ( 
.A1(n_3306),
.A2(n_3166),
.B1(n_2840),
.B2(n_2885),
.Y(n_3375)
);

OAI21x1_ASAP7_75t_L g3376 ( 
.A1(n_3215),
.A2(n_2807),
.B(n_2833),
.Y(n_3376)
);

AO31x2_ASAP7_75t_L g3377 ( 
.A1(n_3234),
.A2(n_3239),
.A3(n_3237),
.B(n_3290),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_3310),
.B(n_3071),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_3265),
.B(n_3162),
.Y(n_3379)
);

OAI22xp5_ASAP7_75t_L g3380 ( 
.A1(n_3187),
.A2(n_3076),
.B1(n_3102),
.B2(n_3162),
.Y(n_3380)
);

INVx3_ASAP7_75t_L g3381 ( 
.A(n_3236),
.Y(n_3381)
);

AOI22xp33_ASAP7_75t_L g3382 ( 
.A1(n_3309),
.A2(n_2814),
.B1(n_3094),
.B2(n_2860),
.Y(n_3382)
);

AOI22xp33_ASAP7_75t_L g3383 ( 
.A1(n_3309),
.A2(n_2814),
.B1(n_3094),
.B2(n_2860),
.Y(n_3383)
);

AOI22xp33_ASAP7_75t_L g3384 ( 
.A1(n_3309),
.A2(n_3094),
.B1(n_2858),
.B2(n_2871),
.Y(n_3384)
);

AOI22xp33_ASAP7_75t_L g3385 ( 
.A1(n_3188),
.A2(n_3094),
.B1(n_2858),
.B2(n_2871),
.Y(n_3385)
);

AOI22xp33_ASAP7_75t_SL g3386 ( 
.A1(n_3187),
.A2(n_3162),
.B1(n_3103),
.B2(n_3125),
.Y(n_3386)
);

AOI222xp33_ASAP7_75t_L g3387 ( 
.A1(n_3188),
.A2(n_3115),
.B1(n_2839),
.B2(n_2928),
.C1(n_2856),
.C2(n_2891),
.Y(n_3387)
);

INVx2_ASAP7_75t_SL g3388 ( 
.A(n_3272),
.Y(n_3388)
);

NAND3xp33_ASAP7_75t_L g3389 ( 
.A(n_3323),
.B(n_3163),
.C(n_3147),
.Y(n_3389)
);

OAI21xp33_ASAP7_75t_L g3390 ( 
.A1(n_3269),
.A2(n_2919),
.B(n_2891),
.Y(n_3390)
);

OAI21x1_ASAP7_75t_L g3391 ( 
.A1(n_3217),
.A2(n_2833),
.B(n_2806),
.Y(n_3391)
);

AOI22xp5_ASAP7_75t_L g3392 ( 
.A1(n_3308),
.A2(n_2891),
.B1(n_2889),
.B2(n_2962),
.Y(n_3392)
);

AND2x4_ASAP7_75t_L g3393 ( 
.A(n_3292),
.B(n_3064),
.Y(n_3393)
);

AOI22xp33_ASAP7_75t_L g3394 ( 
.A1(n_3308),
.A2(n_2869),
.B1(n_2955),
.B2(n_2953),
.Y(n_3394)
);

AOI22xp33_ASAP7_75t_L g3395 ( 
.A1(n_3213),
.A2(n_2869),
.B1(n_2955),
.B2(n_2953),
.Y(n_3395)
);

AOI22xp33_ASAP7_75t_L g3396 ( 
.A1(n_3226),
.A2(n_2937),
.B1(n_2784),
.B2(n_2943),
.Y(n_3396)
);

AOI222xp33_ASAP7_75t_L g3397 ( 
.A1(n_3194),
.A2(n_2839),
.B1(n_2928),
.B2(n_2889),
.C1(n_2962),
.C2(n_2937),
.Y(n_3397)
);

INVx2_ASAP7_75t_L g3398 ( 
.A(n_3169),
.Y(n_3398)
);

AND2x2_ASAP7_75t_L g3399 ( 
.A(n_3265),
.B(n_3103),
.Y(n_3399)
);

AOI22xp33_ASAP7_75t_L g3400 ( 
.A1(n_3226),
.A2(n_2784),
.B1(n_2951),
.B2(n_2943),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3209),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_3254),
.Y(n_3402)
);

OR2x6_ASAP7_75t_L g3403 ( 
.A(n_3266),
.B(n_2872),
.Y(n_3403)
);

AOI22xp33_ASAP7_75t_L g3404 ( 
.A1(n_3226),
.A2(n_2951),
.B1(n_2966),
.B2(n_2875),
.Y(n_3404)
);

INVx2_ASAP7_75t_SL g3405 ( 
.A(n_3272),
.Y(n_3405)
);

OAI22xp5_ASAP7_75t_L g3406 ( 
.A1(n_3187),
.A2(n_3112),
.B1(n_3105),
.B2(n_3028),
.Y(n_3406)
);

AOI22xp33_ASAP7_75t_L g3407 ( 
.A1(n_3193),
.A2(n_2966),
.B1(n_2875),
.B2(n_2880),
.Y(n_3407)
);

INVx3_ASAP7_75t_L g3408 ( 
.A(n_3236),
.Y(n_3408)
);

AND2x2_ASAP7_75t_L g3409 ( 
.A(n_3286),
.B(n_3028),
.Y(n_3409)
);

AND2x4_ASAP7_75t_L g3410 ( 
.A(n_3292),
.B(n_3064),
.Y(n_3410)
);

AND2x2_ASAP7_75t_L g3411 ( 
.A(n_3286),
.B(n_3105),
.Y(n_3411)
);

INVx3_ASAP7_75t_L g3412 ( 
.A(n_3236),
.Y(n_3412)
);

HB1xp67_ASAP7_75t_L g3413 ( 
.A(n_3194),
.Y(n_3413)
);

AOI22xp33_ASAP7_75t_L g3414 ( 
.A1(n_3193),
.A2(n_2880),
.B1(n_2872),
.B2(n_2882),
.Y(n_3414)
);

AOI22xp33_ASAP7_75t_L g3415 ( 
.A1(n_3193),
.A2(n_2882),
.B1(n_2846),
.B2(n_2839),
.Y(n_3415)
);

OAI211xp5_ASAP7_75t_L g3416 ( 
.A1(n_3196),
.A2(n_2928),
.B(n_2839),
.C(n_2948),
.Y(n_3416)
);

INVx2_ASAP7_75t_L g3417 ( 
.A(n_3254),
.Y(n_3417)
);

BUFx6f_ASAP7_75t_L g3418 ( 
.A(n_3303),
.Y(n_3418)
);

BUFx2_ASAP7_75t_L g3419 ( 
.A(n_3279),
.Y(n_3419)
);

OAI211xp5_ASAP7_75t_SL g3420 ( 
.A1(n_3281),
.A2(n_119),
.B(n_116),
.C(n_118),
.Y(n_3420)
);

AND2x4_ASAP7_75t_L g3421 ( 
.A(n_3292),
.B(n_3064),
.Y(n_3421)
);

AOI22xp33_ASAP7_75t_L g3422 ( 
.A1(n_3187),
.A2(n_2846),
.B1(n_2893),
.B2(n_2942),
.Y(n_3422)
);

AOI22xp5_ASAP7_75t_L g3423 ( 
.A1(n_3322),
.A2(n_2893),
.B1(n_3091),
.B2(n_2876),
.Y(n_3423)
);

OR2x2_ASAP7_75t_L g3424 ( 
.A(n_3225),
.B(n_3282),
.Y(n_3424)
);

AOI22xp33_ASAP7_75t_SL g3425 ( 
.A1(n_3187),
.A2(n_2958),
.B1(n_2931),
.B2(n_3091),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3209),
.Y(n_3426)
);

OAI211xp5_ASAP7_75t_L g3427 ( 
.A1(n_3196),
.A2(n_3091),
.B(n_2846),
.C(n_2843),
.Y(n_3427)
);

AO21x2_ASAP7_75t_L g3428 ( 
.A1(n_3280),
.A2(n_2809),
.B(n_2786),
.Y(n_3428)
);

OA21x2_ASAP7_75t_L g3429 ( 
.A1(n_3280),
.A2(n_2824),
.B(n_2850),
.Y(n_3429)
);

INVxp33_ASAP7_75t_SL g3430 ( 
.A(n_3177),
.Y(n_3430)
);

AOI22xp33_ASAP7_75t_L g3431 ( 
.A1(n_3192),
.A2(n_3274),
.B1(n_3278),
.B2(n_3289),
.Y(n_3431)
);

OR2x2_ASAP7_75t_L g3432 ( 
.A(n_3230),
.B(n_2820),
.Y(n_3432)
);

NOR4xp25_ASAP7_75t_L g3433 ( 
.A(n_3274),
.B(n_2940),
.C(n_121),
.D(n_118),
.Y(n_3433)
);

CKINVDCx5p33_ASAP7_75t_R g3434 ( 
.A(n_3305),
.Y(n_3434)
);

BUFx12f_ASAP7_75t_L g3435 ( 
.A(n_3192),
.Y(n_3435)
);

NOR2xp33_ASAP7_75t_L g3436 ( 
.A(n_3192),
.B(n_120),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_3210),
.Y(n_3437)
);

BUFx2_ASAP7_75t_L g3438 ( 
.A(n_3288),
.Y(n_3438)
);

NAND2x1_ASAP7_75t_L g3439 ( 
.A(n_3174),
.B(n_2843),
.Y(n_3439)
);

OAI22xp5_ASAP7_75t_L g3440 ( 
.A1(n_3192),
.A2(n_2876),
.B1(n_2843),
.B2(n_2940),
.Y(n_3440)
);

HB1xp67_ASAP7_75t_L g3441 ( 
.A(n_3182),
.Y(n_3441)
);

AND2x2_ASAP7_75t_L g3442 ( 
.A(n_3291),
.B(n_2820),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3210),
.Y(n_3443)
);

OAI221xp5_ASAP7_75t_L g3444 ( 
.A1(n_3278),
.A2(n_122),
.B1(n_124),
.B2(n_127),
.C(n_128),
.Y(n_3444)
);

OAI221xp5_ASAP7_75t_L g3445 ( 
.A1(n_3192),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.C(n_130),
.Y(n_3445)
);

OAI22xp5_ASAP7_75t_L g3446 ( 
.A1(n_3184),
.A2(n_2940),
.B1(n_2820),
.B2(n_2942),
.Y(n_3446)
);

INVx1_ASAP7_75t_SL g3447 ( 
.A(n_3272),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_3291),
.B(n_2820),
.Y(n_3448)
);

AOI22xp33_ASAP7_75t_L g3449 ( 
.A1(n_3203),
.A2(n_2865),
.B1(n_2868),
.B2(n_2824),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3229),
.Y(n_3450)
);

OAI21x1_ASAP7_75t_SL g3451 ( 
.A1(n_3304),
.A2(n_129),
.B(n_131),
.Y(n_3451)
);

INVx4_ASAP7_75t_R g3452 ( 
.A(n_3288),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3229),
.Y(n_3453)
);

INVx2_ASAP7_75t_L g3454 ( 
.A(n_3202),
.Y(n_3454)
);

OAI221xp5_ASAP7_75t_L g3455 ( 
.A1(n_3185),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.C(n_134),
.Y(n_3455)
);

BUFx2_ASAP7_75t_L g3456 ( 
.A(n_3288),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3231),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3231),
.Y(n_3458)
);

INVx2_ASAP7_75t_L g3459 ( 
.A(n_3179),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3364),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3370),
.Y(n_3461)
);

AOI22xp33_ASAP7_75t_SL g3462 ( 
.A1(n_3349),
.A2(n_3271),
.B1(n_3184),
.B2(n_3203),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3401),
.Y(n_3463)
);

BUFx2_ASAP7_75t_L g3464 ( 
.A(n_3435),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3377),
.Y(n_3465)
);

OAI21xp5_ASAP7_75t_SL g3466 ( 
.A1(n_3334),
.A2(n_3298),
.B(n_3292),
.Y(n_3466)
);

BUFx3_ASAP7_75t_L g3467 ( 
.A(n_3430),
.Y(n_3467)
);

AND2x2_ASAP7_75t_L g3468 ( 
.A(n_3360),
.B(n_3199),
.Y(n_3468)
);

INVx1_ASAP7_75t_SL g3469 ( 
.A(n_3357),
.Y(n_3469)
);

INVx2_ASAP7_75t_L g3470 ( 
.A(n_3377),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3426),
.Y(n_3471)
);

HB1xp67_ASAP7_75t_L g3472 ( 
.A(n_3441),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3351),
.B(n_3199),
.Y(n_3473)
);

AND2x2_ASAP7_75t_L g3474 ( 
.A(n_3351),
.B(n_3199),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3437),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3343),
.B(n_3253),
.Y(n_3476)
);

INVx1_ASAP7_75t_SL g3477 ( 
.A(n_3373),
.Y(n_3477)
);

OR2x2_ASAP7_75t_L g3478 ( 
.A(n_3413),
.B(n_3247),
.Y(n_3478)
);

INVx2_ASAP7_75t_L g3479 ( 
.A(n_3377),
.Y(n_3479)
);

AND2x2_ASAP7_75t_L g3480 ( 
.A(n_3438),
.B(n_3199),
.Y(n_3480)
);

AND2x2_ASAP7_75t_L g3481 ( 
.A(n_3456),
.B(n_3201),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3329),
.B(n_3260),
.Y(n_3482)
);

AND2x2_ASAP7_75t_L g3483 ( 
.A(n_3362),
.B(n_3201),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_3377),
.Y(n_3484)
);

INVxp67_ASAP7_75t_SL g3485 ( 
.A(n_3419),
.Y(n_3485)
);

INVxp67_ASAP7_75t_L g3486 ( 
.A(n_3436),
.Y(n_3486)
);

INVx2_ASAP7_75t_L g3487 ( 
.A(n_3402),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3443),
.Y(n_3488)
);

OR2x2_ASAP7_75t_L g3489 ( 
.A(n_3413),
.B(n_3247),
.Y(n_3489)
);

HB1xp67_ASAP7_75t_L g3490 ( 
.A(n_3441),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_3402),
.Y(n_3491)
);

AOI22xp33_ASAP7_75t_SL g3492 ( 
.A1(n_3346),
.A2(n_3271),
.B1(n_3184),
.B2(n_3203),
.Y(n_3492)
);

AND2x4_ASAP7_75t_L g3493 ( 
.A(n_3381),
.B(n_3174),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3450),
.Y(n_3494)
);

INVxp67_ASAP7_75t_SL g3495 ( 
.A(n_3374),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3329),
.B(n_3296),
.Y(n_3496)
);

AND2x2_ASAP7_75t_L g3497 ( 
.A(n_3362),
.B(n_3201),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3334),
.B(n_3350),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_3417),
.Y(n_3499)
);

NOR2xp67_ASAP7_75t_L g3500 ( 
.A(n_3368),
.B(n_3174),
.Y(n_3500)
);

HB1xp67_ASAP7_75t_L g3501 ( 
.A(n_3424),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3453),
.Y(n_3502)
);

NOR2xp33_ASAP7_75t_L g3503 ( 
.A(n_3434),
.B(n_3201),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3457),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3458),
.Y(n_3505)
);

AND2x4_ASAP7_75t_L g3506 ( 
.A(n_3381),
.B(n_3174),
.Y(n_3506)
);

INVxp67_ASAP7_75t_L g3507 ( 
.A(n_3436),
.Y(n_3507)
);

INVx1_ASAP7_75t_SL g3508 ( 
.A(n_3447),
.Y(n_3508)
);

AND2x2_ASAP7_75t_L g3509 ( 
.A(n_3362),
.B(n_3247),
.Y(n_3509)
);

NOR2xp33_ASAP7_75t_L g3510 ( 
.A(n_3353),
.B(n_3313),
.Y(n_3510)
);

INVx2_ASAP7_75t_L g3511 ( 
.A(n_3417),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3330),
.Y(n_3512)
);

AND2x2_ASAP7_75t_L g3513 ( 
.A(n_3399),
.B(n_3170),
.Y(n_3513)
);

BUFx2_ASAP7_75t_L g3514 ( 
.A(n_3418),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3335),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3338),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3342),
.Y(n_3517)
);

AOI22xp33_ASAP7_75t_L g3518 ( 
.A1(n_3331),
.A2(n_3271),
.B1(n_3184),
.B2(n_3298),
.Y(n_3518)
);

CKINVDCx20_ASAP7_75t_R g3519 ( 
.A(n_3378),
.Y(n_3519)
);

INVx4_ASAP7_75t_L g3520 ( 
.A(n_3365),
.Y(n_3520)
);

HB1xp67_ASAP7_75t_L g3521 ( 
.A(n_3332),
.Y(n_3521)
);

AND2x2_ASAP7_75t_L g3522 ( 
.A(n_3379),
.B(n_3170),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3354),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3356),
.Y(n_3524)
);

INVx2_ASAP7_75t_L g3525 ( 
.A(n_3359),
.Y(n_3525)
);

AND2x2_ASAP7_75t_L g3526 ( 
.A(n_3409),
.B(n_3320),
.Y(n_3526)
);

BUFx2_ASAP7_75t_L g3527 ( 
.A(n_3418),
.Y(n_3527)
);

BUFx3_ASAP7_75t_L g3528 ( 
.A(n_3388),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3359),
.Y(n_3529)
);

HB1xp67_ASAP7_75t_L g3530 ( 
.A(n_3332),
.Y(n_3530)
);

AND2x2_ASAP7_75t_L g3531 ( 
.A(n_3411),
.B(n_3320),
.Y(n_3531)
);

AND2x2_ASAP7_75t_L g3532 ( 
.A(n_3340),
.B(n_3242),
.Y(n_3532)
);

OR2x2_ASAP7_75t_L g3533 ( 
.A(n_3332),
.B(n_3189),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3361),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3361),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3398),
.Y(n_3536)
);

INVxp67_ASAP7_75t_L g3537 ( 
.A(n_3405),
.Y(n_3537)
);

INVxp67_ASAP7_75t_L g3538 ( 
.A(n_3327),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3345),
.B(n_3296),
.Y(n_3539)
);

AND2x2_ASAP7_75t_L g3540 ( 
.A(n_3442),
.B(n_3242),
.Y(n_3540)
);

INVx2_ASAP7_75t_L g3541 ( 
.A(n_3398),
.Y(n_3541)
);

NOR2xp33_ASAP7_75t_L g3542 ( 
.A(n_3386),
.B(n_3283),
.Y(n_3542)
);

INVx3_ASAP7_75t_L g3543 ( 
.A(n_3418),
.Y(n_3543)
);

HB1xp67_ASAP7_75t_L g3544 ( 
.A(n_3418),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3459),
.Y(n_3545)
);

AND2x2_ASAP7_75t_L g3546 ( 
.A(n_3448),
.B(n_3171),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3459),
.Y(n_3547)
);

OR2x2_ASAP7_75t_L g3548 ( 
.A(n_3432),
.B(n_3189),
.Y(n_3548)
);

OR2x2_ASAP7_75t_L g3549 ( 
.A(n_3431),
.B(n_3294),
.Y(n_3549)
);

HB1xp67_ASAP7_75t_L g3550 ( 
.A(n_3408),
.Y(n_3550)
);

AND2x4_ASAP7_75t_L g3551 ( 
.A(n_3408),
.B(n_3298),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3345),
.B(n_3301),
.Y(n_3552)
);

AND2x2_ASAP7_75t_L g3553 ( 
.A(n_3393),
.B(n_3171),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3412),
.Y(n_3554)
);

AND2x2_ASAP7_75t_L g3555 ( 
.A(n_3393),
.B(n_3283),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3412),
.Y(n_3556)
);

HB1xp67_ASAP7_75t_L g3557 ( 
.A(n_3403),
.Y(n_3557)
);

AND2x2_ASAP7_75t_L g3558 ( 
.A(n_3410),
.B(n_3284),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3452),
.Y(n_3559)
);

AND2x2_ASAP7_75t_L g3560 ( 
.A(n_3410),
.B(n_3284),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_3431),
.B(n_3301),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_3328),
.Y(n_3562)
);

NOR2x1_ASAP7_75t_L g3563 ( 
.A(n_3358),
.B(n_3298),
.Y(n_3563)
);

AND2x4_ASAP7_75t_L g3564 ( 
.A(n_3403),
.B(n_3234),
.Y(n_3564)
);

AND2x4_ASAP7_75t_L g3565 ( 
.A(n_3403),
.B(n_3234),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3371),
.B(n_3302),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3333),
.Y(n_3567)
);

BUFx3_ASAP7_75t_L g3568 ( 
.A(n_3451),
.Y(n_3568)
);

AND2x2_ASAP7_75t_L g3569 ( 
.A(n_3421),
.B(n_3299),
.Y(n_3569)
);

INVx2_ASAP7_75t_L g3570 ( 
.A(n_3337),
.Y(n_3570)
);

AND2x2_ASAP7_75t_L g3571 ( 
.A(n_3421),
.B(n_3299),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3454),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3352),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3348),
.Y(n_3574)
);

AND2x2_ASAP7_75t_L g3575 ( 
.A(n_3366),
.B(n_3300),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3439),
.Y(n_3576)
);

OR2x2_ASAP7_75t_L g3577 ( 
.A(n_3427),
.B(n_3294),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_3429),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3371),
.B(n_3302),
.Y(n_3579)
);

INVx2_ASAP7_75t_L g3580 ( 
.A(n_3429),
.Y(n_3580)
);

INVx4_ASAP7_75t_L g3581 ( 
.A(n_3365),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3433),
.B(n_3294),
.Y(n_3582)
);

AND2x4_ASAP7_75t_SL g3583 ( 
.A(n_3367),
.B(n_3293),
.Y(n_3583)
);

HB1xp67_ASAP7_75t_L g3584 ( 
.A(n_3341),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3416),
.Y(n_3585)
);

INVx1_ASAP7_75t_SL g3586 ( 
.A(n_3406),
.Y(n_3586)
);

AOI22xp5_ASAP7_75t_L g3587 ( 
.A1(n_3585),
.A2(n_3344),
.B1(n_3336),
.B2(n_3387),
.Y(n_3587)
);

AND2x2_ASAP7_75t_L g3588 ( 
.A(n_3553),
.B(n_3297),
.Y(n_3588)
);

AOI221xp5_ASAP7_75t_L g3589 ( 
.A1(n_3585),
.A2(n_3455),
.B1(n_3445),
.B2(n_3420),
.C(n_3444),
.Y(n_3589)
);

OAI21xp5_ASAP7_75t_L g3590 ( 
.A1(n_3492),
.A2(n_3339),
.B(n_3347),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3514),
.Y(n_3591)
);

AOI322xp5_ASAP7_75t_L g3592 ( 
.A1(n_3498),
.A2(n_3347),
.A3(n_3339),
.B1(n_3358),
.B2(n_3372),
.C1(n_3369),
.C2(n_3375),
.Y(n_3592)
);

OAI22xp5_ASAP7_75t_L g3593 ( 
.A1(n_3469),
.A2(n_3369),
.B1(n_3375),
.B2(n_3382),
.Y(n_3593)
);

AOI221xp5_ASAP7_75t_L g3594 ( 
.A1(n_3462),
.A2(n_3355),
.B1(n_3383),
.B2(n_3382),
.C(n_3380),
.Y(n_3594)
);

BUFx2_ASAP7_75t_L g3595 ( 
.A(n_3519),
.Y(n_3595)
);

NOR4xp25_ASAP7_75t_SL g3596 ( 
.A(n_3466),
.B(n_3195),
.C(n_3390),
.D(n_3318),
.Y(n_3596)
);

INVx2_ASAP7_75t_L g3597 ( 
.A(n_3514),
.Y(n_3597)
);

OAI211xp5_ASAP7_75t_L g3598 ( 
.A1(n_3563),
.A2(n_3397),
.B(n_3383),
.C(n_3384),
.Y(n_3598)
);

OAI21xp5_ASAP7_75t_SL g3599 ( 
.A1(n_3477),
.A2(n_3363),
.B(n_3384),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3472),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3486),
.B(n_3232),
.Y(n_3601)
);

NAND3xp33_ASAP7_75t_L g3602 ( 
.A(n_3521),
.B(n_3389),
.C(n_3407),
.Y(n_3602)
);

BUFx2_ASAP7_75t_L g3603 ( 
.A(n_3519),
.Y(n_3603)
);

AOI222xp33_ASAP7_75t_L g3604 ( 
.A1(n_3507),
.A2(n_3415),
.B1(n_3440),
.B2(n_3407),
.C1(n_3239),
.C2(n_3237),
.Y(n_3604)
);

AND2x4_ASAP7_75t_SL g3605 ( 
.A(n_3520),
.B(n_3392),
.Y(n_3605)
);

OAI221xp5_ASAP7_75t_L g3606 ( 
.A1(n_3518),
.A2(n_3415),
.B1(n_3385),
.B2(n_3425),
.C(n_3423),
.Y(n_3606)
);

OR2x2_ASAP7_75t_L g3607 ( 
.A(n_3495),
.B(n_3175),
.Y(n_3607)
);

INVx2_ASAP7_75t_L g3608 ( 
.A(n_3527),
.Y(n_3608)
);

OAI221xp5_ASAP7_75t_L g3609 ( 
.A1(n_3584),
.A2(n_3385),
.B1(n_3404),
.B2(n_3395),
.C(n_3396),
.Y(n_3609)
);

NAND4xp25_ASAP7_75t_L g3610 ( 
.A(n_3539),
.B(n_3404),
.C(n_3400),
.D(n_3396),
.Y(n_3610)
);

NAND3xp33_ASAP7_75t_L g3611 ( 
.A(n_3530),
.B(n_3400),
.C(n_3395),
.Y(n_3611)
);

OAI33xp33_ASAP7_75t_L g3612 ( 
.A1(n_3552),
.A2(n_3290),
.A3(n_3232),
.B1(n_3233),
.B2(n_3248),
.B3(n_3246),
.Y(n_3612)
);

OAI221xp5_ASAP7_75t_SL g3613 ( 
.A1(n_3482),
.A2(n_3414),
.B1(n_3394),
.B2(n_3449),
.C(n_3422),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3490),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_SL g3615 ( 
.A(n_3500),
.B(n_3271),
.Y(n_3615)
);

NOR2xp33_ASAP7_75t_R g3616 ( 
.A(n_3467),
.B(n_132),
.Y(n_3616)
);

INVx2_ASAP7_75t_L g3617 ( 
.A(n_3527),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3553),
.B(n_3569),
.Y(n_3618)
);

AO21x2_ASAP7_75t_L g3619 ( 
.A1(n_3473),
.A2(n_3239),
.B(n_3237),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3508),
.B(n_3496),
.Y(n_3620)
);

AOI22xp33_ASAP7_75t_L g3621 ( 
.A1(n_3510),
.A2(n_3317),
.B1(n_3446),
.B2(n_3414),
.Y(n_3621)
);

OAI221xp5_ASAP7_75t_SL g3622 ( 
.A1(n_3566),
.A2(n_3579),
.B1(n_3582),
.B2(n_3568),
.C(n_3586),
.Y(n_3622)
);

BUFx2_ASAP7_75t_L g3623 ( 
.A(n_3485),
.Y(n_3623)
);

INVx2_ASAP7_75t_L g3624 ( 
.A(n_3464),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3460),
.Y(n_3625)
);

NAND4xp25_ASAP7_75t_L g3626 ( 
.A(n_3568),
.B(n_3449),
.C(n_3394),
.D(n_3422),
.Y(n_3626)
);

INVx2_ASAP7_75t_L g3627 ( 
.A(n_3473),
.Y(n_3627)
);

NOR3xp33_ASAP7_75t_L g3628 ( 
.A(n_3520),
.B(n_3376),
.C(n_3391),
.Y(n_3628)
);

AOI222xp33_ASAP7_75t_L g3629 ( 
.A1(n_3561),
.A2(n_3233),
.B1(n_3248),
.B2(n_3246),
.C1(n_3195),
.C2(n_3252),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3460),
.Y(n_3630)
);

OA222x2_ASAP7_75t_L g3631 ( 
.A1(n_3533),
.A2(n_3212),
.B1(n_3287),
.B2(n_3280),
.C1(n_3262),
.C2(n_3324),
.Y(n_3631)
);

AOI221xp5_ASAP7_75t_L g3632 ( 
.A1(n_3501),
.A2(n_3252),
.B1(n_3178),
.B2(n_3181),
.C(n_3214),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3461),
.Y(n_3633)
);

BUFx3_ASAP7_75t_L g3634 ( 
.A(n_3467),
.Y(n_3634)
);

AND2x2_ASAP7_75t_L g3635 ( 
.A(n_3569),
.B(n_3297),
.Y(n_3635)
);

AND2x2_ASAP7_75t_L g3636 ( 
.A(n_3571),
.B(n_3300),
.Y(n_3636)
);

AOI221xp5_ASAP7_75t_L g3637 ( 
.A1(n_3538),
.A2(n_3178),
.B1(n_3181),
.B2(n_3214),
.C(n_3238),
.Y(n_3637)
);

OAI22xp33_ASAP7_75t_L g3638 ( 
.A1(n_3559),
.A2(n_3464),
.B1(n_3581),
.B2(n_3520),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3461),
.Y(n_3639)
);

NOR2xp33_ASAP7_75t_R g3640 ( 
.A(n_3581),
.B(n_134),
.Y(n_3640)
);

HB1xp67_ASAP7_75t_L g3641 ( 
.A(n_3463),
.Y(n_3641)
);

HB1xp67_ASAP7_75t_L g3642 ( 
.A(n_3463),
.Y(n_3642)
);

INVx2_ASAP7_75t_L g3643 ( 
.A(n_3474),
.Y(n_3643)
);

INVxp67_ASAP7_75t_L g3644 ( 
.A(n_3528),
.Y(n_3644)
);

INVx1_ASAP7_75t_SL g3645 ( 
.A(n_3528),
.Y(n_3645)
);

AOI22xp33_ASAP7_75t_L g3646 ( 
.A1(n_3542),
.A2(n_3581),
.B1(n_3476),
.B2(n_3549),
.Y(n_3646)
);

OA21x2_ASAP7_75t_L g3647 ( 
.A1(n_3578),
.A2(n_3287),
.B(n_3208),
.Y(n_3647)
);

NOR2xp33_ASAP7_75t_L g3648 ( 
.A(n_3503),
.B(n_3257),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_3543),
.Y(n_3649)
);

AOI221x1_ASAP7_75t_L g3650 ( 
.A1(n_3543),
.A2(n_3318),
.B1(n_3312),
.B2(n_3303),
.C(n_3315),
.Y(n_3650)
);

HB1xp67_ASAP7_75t_L g3651 ( 
.A(n_3475),
.Y(n_3651)
);

OAI221xp5_ASAP7_75t_L g3652 ( 
.A1(n_3537),
.A2(n_3263),
.B1(n_3264),
.B2(n_3238),
.C(n_3250),
.Y(n_3652)
);

INVxp67_ASAP7_75t_L g3653 ( 
.A(n_3550),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3475),
.Y(n_3654)
);

INVxp67_ASAP7_75t_L g3655 ( 
.A(n_3544),
.Y(n_3655)
);

OAI22xp5_ASAP7_75t_L g3656 ( 
.A1(n_3583),
.A2(n_3271),
.B1(n_3184),
.B2(n_3211),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3571),
.B(n_3326),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3474),
.Y(n_3658)
);

NAND3xp33_ASAP7_75t_L g3659 ( 
.A(n_3533),
.B(n_3317),
.C(n_3176),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_3543),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3494),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3494),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_SL g3663 ( 
.A(n_3468),
.B(n_3271),
.Y(n_3663)
);

OA21x2_ASAP7_75t_L g3664 ( 
.A1(n_3578),
.A2(n_3287),
.B(n_3208),
.Y(n_3664)
);

AND2x2_ASAP7_75t_L g3665 ( 
.A(n_3526),
.B(n_3531),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3465),
.Y(n_3666)
);

OAI33xp33_ASAP7_75t_L g3667 ( 
.A1(n_3502),
.A2(n_3250),
.A3(n_3235),
.B1(n_3212),
.B2(n_3257),
.B3(n_3172),
.Y(n_3667)
);

AOI221xp5_ASAP7_75t_L g3668 ( 
.A1(n_3557),
.A2(n_3235),
.B1(n_3259),
.B2(n_3263),
.C(n_3264),
.Y(n_3668)
);

AND2x2_ASAP7_75t_L g3669 ( 
.A(n_3526),
.B(n_3326),
.Y(n_3669)
);

OR2x2_ASAP7_75t_L g3670 ( 
.A(n_3573),
.B(n_3230),
.Y(n_3670)
);

OAI22xp5_ASAP7_75t_L g3671 ( 
.A1(n_3583),
.A2(n_3211),
.B1(n_3173),
.B2(n_3304),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3573),
.B(n_3285),
.Y(n_3672)
);

NOR2x1_ASAP7_75t_L g3673 ( 
.A(n_3554),
.B(n_3556),
.Y(n_3673)
);

BUFx3_ASAP7_75t_L g3674 ( 
.A(n_3493),
.Y(n_3674)
);

OAI21x1_ASAP7_75t_L g3675 ( 
.A1(n_3576),
.A2(n_3217),
.B(n_3228),
.Y(n_3675)
);

OAI332xp33_ASAP7_75t_L g3676 ( 
.A1(n_3577),
.A2(n_3312),
.A3(n_3321),
.B1(n_3307),
.B2(n_3304),
.B3(n_3172),
.C1(n_3207),
.C2(n_3186),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3465),
.Y(n_3677)
);

INVx1_ASAP7_75t_SL g3678 ( 
.A(n_3531),
.Y(n_3678)
);

OAI321xp33_ASAP7_75t_L g3679 ( 
.A1(n_3468),
.A2(n_3321),
.A3(n_3307),
.B1(n_3303),
.B2(n_3315),
.C(n_3314),
.Y(n_3679)
);

AND2x2_ASAP7_75t_L g3680 ( 
.A(n_3555),
.B(n_3285),
.Y(n_3680)
);

OR2x2_ASAP7_75t_L g3681 ( 
.A(n_3549),
.B(n_3259),
.Y(n_3681)
);

INVx1_ASAP7_75t_SL g3682 ( 
.A(n_3480),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3502),
.Y(n_3683)
);

AND2x2_ASAP7_75t_L g3684 ( 
.A(n_3555),
.B(n_3273),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3504),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3572),
.B(n_3273),
.Y(n_3686)
);

NAND3xp33_ASAP7_75t_L g3687 ( 
.A(n_3572),
.B(n_3317),
.C(n_3176),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3470),
.Y(n_3688)
);

OAI22xp33_ASAP7_75t_L g3689 ( 
.A1(n_3577),
.A2(n_3317),
.B1(n_3315),
.B2(n_3303),
.Y(n_3689)
);

AOI222xp33_ASAP7_75t_L g3690 ( 
.A1(n_3532),
.A2(n_3211),
.B1(n_3173),
.B2(n_3227),
.C1(n_3240),
.C2(n_3241),
.Y(n_3690)
);

INVx2_ASAP7_75t_L g3691 ( 
.A(n_3470),
.Y(n_3691)
);

AOI22xp33_ASAP7_75t_L g3692 ( 
.A1(n_3471),
.A2(n_3488),
.B1(n_3565),
.B2(n_3564),
.Y(n_3692)
);

AOI22xp33_ASAP7_75t_L g3693 ( 
.A1(n_3564),
.A2(n_3176),
.B1(n_3249),
.B2(n_3255),
.Y(n_3693)
);

AND2x2_ASAP7_75t_L g3694 ( 
.A(n_3558),
.B(n_3325),
.Y(n_3694)
);

AOI22xp33_ASAP7_75t_L g3695 ( 
.A1(n_3564),
.A2(n_3176),
.B1(n_3249),
.B2(n_3255),
.Y(n_3695)
);

AOI22xp33_ASAP7_75t_L g3696 ( 
.A1(n_3565),
.A2(n_3249),
.B1(n_3258),
.B2(n_3173),
.Y(n_3696)
);

BUFx3_ASAP7_75t_L g3697 ( 
.A(n_3493),
.Y(n_3697)
);

HB1xp67_ASAP7_75t_L g3698 ( 
.A(n_3504),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3505),
.Y(n_3699)
);

AO21x2_ASAP7_75t_L g3700 ( 
.A1(n_3576),
.A2(n_3321),
.B(n_3307),
.Y(n_3700)
);

AOI22xp33_ASAP7_75t_L g3701 ( 
.A1(n_3565),
.A2(n_3258),
.B1(n_3173),
.B2(n_3211),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3493),
.Y(n_3702)
);

AOI211xp5_ASAP7_75t_L g3703 ( 
.A1(n_3590),
.A2(n_3532),
.B(n_3497),
.C(n_3483),
.Y(n_3703)
);

NOR2xp33_ASAP7_75t_L g3704 ( 
.A(n_3634),
.B(n_3575),
.Y(n_3704)
);

NOR3xp33_ASAP7_75t_L g3705 ( 
.A(n_3622),
.B(n_3491),
.C(n_3487),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3641),
.Y(n_3706)
);

BUFx3_ASAP7_75t_L g3707 ( 
.A(n_3595),
.Y(n_3707)
);

NOR2x1_ASAP7_75t_L g3708 ( 
.A(n_3634),
.B(n_3480),
.Y(n_3708)
);

AOI211xp5_ASAP7_75t_L g3709 ( 
.A1(n_3599),
.A2(n_3497),
.B(n_3483),
.C(n_3509),
.Y(n_3709)
);

OR2x2_ASAP7_75t_L g3710 ( 
.A(n_3620),
.B(n_3505),
.Y(n_3710)
);

OR2x2_ASAP7_75t_L g3711 ( 
.A(n_3607),
.B(n_3478),
.Y(n_3711)
);

AOI221xp5_ASAP7_75t_L g3712 ( 
.A1(n_3589),
.A2(n_3547),
.B1(n_3545),
.B2(n_3499),
.C(n_3511),
.Y(n_3712)
);

NAND3xp33_ASAP7_75t_L g3713 ( 
.A(n_3602),
.B(n_3491),
.C(n_3487),
.Y(n_3713)
);

AOI211xp5_ASAP7_75t_L g3714 ( 
.A1(n_3593),
.A2(n_3509),
.B(n_3481),
.C(n_3506),
.Y(n_3714)
);

OR2x2_ASAP7_75t_L g3715 ( 
.A(n_3623),
.B(n_3624),
.Y(n_3715)
);

OR2x2_ASAP7_75t_L g3716 ( 
.A(n_3678),
.B(n_3478),
.Y(n_3716)
);

NAND3xp33_ASAP7_75t_L g3717 ( 
.A(n_3592),
.B(n_3587),
.C(n_3611),
.Y(n_3717)
);

AO21x2_ASAP7_75t_L g3718 ( 
.A1(n_3640),
.A2(n_3484),
.B(n_3479),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3603),
.B(n_3558),
.Y(n_3719)
);

AND2x2_ASAP7_75t_L g3720 ( 
.A(n_3665),
.B(n_3560),
.Y(n_3720)
);

AND2x2_ASAP7_75t_L g3721 ( 
.A(n_3618),
.B(n_3560),
.Y(n_3721)
);

BUFx2_ASAP7_75t_L g3722 ( 
.A(n_3674),
.Y(n_3722)
);

AND2x4_ASAP7_75t_L g3723 ( 
.A(n_3645),
.B(n_3481),
.Y(n_3723)
);

AOI22xp33_ASAP7_75t_L g3724 ( 
.A1(n_3594),
.A2(n_3610),
.B1(n_3646),
.B2(n_3626),
.Y(n_3724)
);

OAI211xp5_ASAP7_75t_L g3725 ( 
.A1(n_3616),
.A2(n_3489),
.B(n_3511),
.C(n_3499),
.Y(n_3725)
);

INVxp67_ASAP7_75t_L g3726 ( 
.A(n_3591),
.Y(n_3726)
);

NOR2xp33_ASAP7_75t_L g3727 ( 
.A(n_3638),
.B(n_3575),
.Y(n_3727)
);

NAND2x1_ASAP7_75t_L g3728 ( 
.A(n_3679),
.B(n_3673),
.Y(n_3728)
);

AND2x2_ASAP7_75t_L g3729 ( 
.A(n_3644),
.B(n_3522),
.Y(n_3729)
);

OR2x2_ASAP7_75t_L g3730 ( 
.A(n_3682),
.B(n_3489),
.Y(n_3730)
);

NOR2xp33_ASAP7_75t_L g3731 ( 
.A(n_3638),
.B(n_3522),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3605),
.B(n_3513),
.Y(n_3732)
);

AOI22xp5_ASAP7_75t_L g3733 ( 
.A1(n_3598),
.A2(n_3551),
.B1(n_3513),
.B2(n_3506),
.Y(n_3733)
);

NAND4xp75_ASAP7_75t_L g3734 ( 
.A(n_3663),
.B(n_3574),
.C(n_3529),
.D(n_3534),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3605),
.B(n_3546),
.Y(n_3735)
);

AOI22xp33_ASAP7_75t_L g3736 ( 
.A1(n_3646),
.A2(n_3567),
.B1(n_3570),
.B2(n_3562),
.Y(n_3736)
);

NOR2x1_ASAP7_75t_L g3737 ( 
.A(n_3615),
.B(n_3506),
.Y(n_3737)
);

AO21x2_ASAP7_75t_L g3738 ( 
.A1(n_3640),
.A2(n_3484),
.B(n_3479),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3674),
.Y(n_3739)
);

AND2x2_ASAP7_75t_L g3740 ( 
.A(n_3694),
.B(n_3546),
.Y(n_3740)
);

NAND4xp75_ASAP7_75t_L g3741 ( 
.A(n_3663),
.B(n_3574),
.C(n_3529),
.D(n_3534),
.Y(n_3741)
);

INVx2_ASAP7_75t_L g3742 ( 
.A(n_3697),
.Y(n_3742)
);

AOI22xp33_ASAP7_75t_L g3743 ( 
.A1(n_3609),
.A2(n_3567),
.B1(n_3570),
.B2(n_3562),
.Y(n_3743)
);

NOR3xp33_ASAP7_75t_L g3744 ( 
.A(n_3613),
.B(n_3536),
.C(n_3535),
.Y(n_3744)
);

AND2x4_ASAP7_75t_L g3745 ( 
.A(n_3697),
.B(n_3591),
.Y(n_3745)
);

OR2x2_ASAP7_75t_L g3746 ( 
.A(n_3600),
.B(n_3548),
.Y(n_3746)
);

NAND3xp33_ASAP7_75t_L g3747 ( 
.A(n_3604),
.B(n_3541),
.C(n_3525),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3641),
.Y(n_3748)
);

NOR2x1_ASAP7_75t_L g3749 ( 
.A(n_3615),
.B(n_3551),
.Y(n_3749)
);

BUFx3_ASAP7_75t_L g3750 ( 
.A(n_3614),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_3700),
.Y(n_3751)
);

OR2x2_ASAP7_75t_L g3752 ( 
.A(n_3655),
.B(n_3548),
.Y(n_3752)
);

OA211x2_ASAP7_75t_L g3753 ( 
.A1(n_3653),
.A2(n_3551),
.B(n_3315),
.C(n_3303),
.Y(n_3753)
);

AND2x2_ASAP7_75t_L g3754 ( 
.A(n_3684),
.B(n_3540),
.Y(n_3754)
);

OR2x2_ASAP7_75t_L g3755 ( 
.A(n_3601),
.B(n_3512),
.Y(n_3755)
);

NAND4xp75_ASAP7_75t_L g3756 ( 
.A(n_3650),
.B(n_3523),
.C(n_3515),
.D(n_3517),
.Y(n_3756)
);

AND2x2_ASAP7_75t_L g3757 ( 
.A(n_3680),
.B(n_3540),
.Y(n_3757)
);

AND2x2_ASAP7_75t_L g3758 ( 
.A(n_3636),
.B(n_3516),
.Y(n_3758)
);

NOR2xp33_ASAP7_75t_L g3759 ( 
.A(n_3676),
.B(n_3524),
.Y(n_3759)
);

BUFx3_ASAP7_75t_L g3760 ( 
.A(n_3702),
.Y(n_3760)
);

NOR3xp33_ASAP7_75t_L g3761 ( 
.A(n_3606),
.B(n_3580),
.C(n_3541),
.Y(n_3761)
);

INVx3_ASAP7_75t_L g3762 ( 
.A(n_3700),
.Y(n_3762)
);

AOI22xp5_ASAP7_75t_L g3763 ( 
.A1(n_3621),
.A2(n_3523),
.B1(n_3525),
.B2(n_3314),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3642),
.Y(n_3764)
);

NAND3xp33_ASAP7_75t_L g3765 ( 
.A(n_3621),
.B(n_3580),
.C(n_3429),
.Y(n_3765)
);

NOR3xp33_ASAP7_75t_SL g3766 ( 
.A(n_3656),
.B(n_3241),
.C(n_3240),
.Y(n_3766)
);

BUFx12f_ASAP7_75t_L g3767 ( 
.A(n_3616),
.Y(n_3767)
);

NOR3xp33_ASAP7_75t_L g3768 ( 
.A(n_3689),
.B(n_3168),
.C(n_135),
.Y(n_3768)
);

NOR3xp33_ASAP7_75t_L g3769 ( 
.A(n_3689),
.B(n_3612),
.C(n_3608),
.Y(n_3769)
);

AOI22xp33_ASAP7_75t_L g3770 ( 
.A1(n_3629),
.A2(n_3628),
.B1(n_3667),
.B2(n_3692),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3642),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3651),
.Y(n_3772)
);

INVx2_ASAP7_75t_L g3773 ( 
.A(n_3660),
.Y(n_3773)
);

AOI22xp33_ASAP7_75t_SL g3774 ( 
.A1(n_3596),
.A2(n_3315),
.B1(n_3303),
.B2(n_3168),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3597),
.B(n_3608),
.Y(n_3775)
);

NOR2x1_ASAP7_75t_L g3776 ( 
.A(n_3597),
.B(n_3324),
.Y(n_3776)
);

AND2x2_ASAP7_75t_L g3777 ( 
.A(n_3588),
.B(n_3277),
.Y(n_3777)
);

AND2x2_ASAP7_75t_L g3778 ( 
.A(n_3635),
.B(n_3277),
.Y(n_3778)
);

AND2x2_ASAP7_75t_L g3779 ( 
.A(n_3657),
.B(n_3324),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3617),
.B(n_3186),
.Y(n_3780)
);

AOI22xp33_ASAP7_75t_SL g3781 ( 
.A1(n_3659),
.A2(n_3631),
.B1(n_3643),
.B2(n_3627),
.Y(n_3781)
);

AND2x2_ASAP7_75t_L g3782 ( 
.A(n_3669),
.B(n_3324),
.Y(n_3782)
);

OR2x2_ASAP7_75t_L g3783 ( 
.A(n_3672),
.B(n_3261),
.Y(n_3783)
);

AOI221xp5_ASAP7_75t_L g3784 ( 
.A1(n_3692),
.A2(n_3227),
.B1(n_3191),
.B2(n_3206),
.C(n_3207),
.Y(n_3784)
);

AND2x4_ASAP7_75t_SL g3785 ( 
.A(n_3617),
.B(n_3315),
.Y(n_3785)
);

BUFx12f_ASAP7_75t_L g3786 ( 
.A(n_3681),
.Y(n_3786)
);

NAND3xp33_ASAP7_75t_L g3787 ( 
.A(n_3649),
.B(n_3206),
.C(n_3191),
.Y(n_3787)
);

AND2x2_ASAP7_75t_L g3788 ( 
.A(n_3648),
.B(n_3262),
.Y(n_3788)
);

NAND3xp33_ASAP7_75t_L g3789 ( 
.A(n_3625),
.B(n_3261),
.C(n_3218),
.Y(n_3789)
);

OAI22xp5_ASAP7_75t_L g3790 ( 
.A1(n_3696),
.A2(n_3202),
.B1(n_3224),
.B2(n_3221),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3648),
.B(n_3244),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3630),
.B(n_3220),
.Y(n_3792)
);

AND2x4_ASAP7_75t_L g3793 ( 
.A(n_3660),
.B(n_3224),
.Y(n_3793)
);

AND2x2_ASAP7_75t_L g3794 ( 
.A(n_3671),
.B(n_3244),
.Y(n_3794)
);

AND2x2_ASAP7_75t_L g3795 ( 
.A(n_3719),
.B(n_3690),
.Y(n_3795)
);

INVx2_ASAP7_75t_L g3796 ( 
.A(n_3707),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3775),
.Y(n_3797)
);

OAI22xp5_ASAP7_75t_L g3798 ( 
.A1(n_3781),
.A2(n_3701),
.B1(n_3696),
.B2(n_3632),
.Y(n_3798)
);

AOI22xp33_ASAP7_75t_L g3799 ( 
.A1(n_3717),
.A2(n_3724),
.B1(n_3761),
.B2(n_3759),
.Y(n_3799)
);

AND2x2_ASAP7_75t_L g3800 ( 
.A(n_3732),
.B(n_3686),
.Y(n_3800)
);

INVxp67_ASAP7_75t_SL g3801 ( 
.A(n_3767),
.Y(n_3801)
);

INVx2_ASAP7_75t_L g3802 ( 
.A(n_3745),
.Y(n_3802)
);

INVx2_ASAP7_75t_SL g3803 ( 
.A(n_3723),
.Y(n_3803)
);

OR2x2_ASAP7_75t_L g3804 ( 
.A(n_3715),
.B(n_3670),
.Y(n_3804)
);

INVx6_ASAP7_75t_L g3805 ( 
.A(n_3745),
.Y(n_3805)
);

AOI221xp5_ASAP7_75t_L g3806 ( 
.A1(n_3724),
.A2(n_3687),
.B1(n_3695),
.B2(n_3693),
.C(n_3651),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_3723),
.B(n_3633),
.Y(n_3807)
);

INVxp67_ASAP7_75t_L g3808 ( 
.A(n_3718),
.Y(n_3808)
);

INVx4_ASAP7_75t_L g3809 ( 
.A(n_3722),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3775),
.Y(n_3810)
);

AO21x2_ASAP7_75t_L g3811 ( 
.A1(n_3718),
.A2(n_3698),
.B(n_3643),
.Y(n_3811)
);

HB1xp67_ASAP7_75t_L g3812 ( 
.A(n_3738),
.Y(n_3812)
);

OR2x2_ASAP7_75t_L g3813 ( 
.A(n_3711),
.B(n_3627),
.Y(n_3813)
);

BUFx6f_ASAP7_75t_L g3814 ( 
.A(n_3738),
.Y(n_3814)
);

INVx3_ASAP7_75t_L g3815 ( 
.A(n_3785),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3706),
.Y(n_3816)
);

AND2x2_ASAP7_75t_L g3817 ( 
.A(n_3735),
.B(n_3658),
.Y(n_3817)
);

AOI33xp33_ASAP7_75t_L g3818 ( 
.A1(n_3781),
.A2(n_3693),
.A3(n_3695),
.B1(n_3658),
.B2(n_3662),
.B3(n_3699),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3748),
.Y(n_3819)
);

INVx2_ASAP7_75t_L g3820 ( 
.A(n_3762),
.Y(n_3820)
);

AND2x2_ASAP7_75t_L g3821 ( 
.A(n_3720),
.B(n_3639),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3764),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3771),
.Y(n_3823)
);

INVx2_ASAP7_75t_L g3824 ( 
.A(n_3776),
.Y(n_3824)
);

NAND3xp33_ASAP7_75t_SL g3825 ( 
.A(n_3768),
.B(n_3668),
.C(n_3637),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3772),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3726),
.Y(n_3827)
);

CKINVDCx5p33_ASAP7_75t_R g3828 ( 
.A(n_3750),
.Y(n_3828)
);

OAI211xp5_ASAP7_75t_L g3829 ( 
.A1(n_3768),
.A2(n_3701),
.B(n_3698),
.C(n_3654),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3762),
.Y(n_3830)
);

AOI22xp33_ASAP7_75t_L g3831 ( 
.A1(n_3761),
.A2(n_3770),
.B1(n_3769),
.B2(n_3786),
.Y(n_3831)
);

OAI22xp5_ASAP7_75t_L g3832 ( 
.A1(n_3774),
.A2(n_3652),
.B1(n_3683),
.B2(n_3661),
.Y(n_3832)
);

OR2x2_ASAP7_75t_L g3833 ( 
.A(n_3716),
.B(n_3685),
.Y(n_3833)
);

OAI22xp5_ASAP7_75t_L g3834 ( 
.A1(n_3774),
.A2(n_3691),
.B1(n_3666),
.B2(n_3688),
.Y(n_3834)
);

INVx2_ASAP7_75t_L g3835 ( 
.A(n_3708),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3726),
.Y(n_3836)
);

INVxp67_ASAP7_75t_L g3837 ( 
.A(n_3725),
.Y(n_3837)
);

NOR2xp33_ASAP7_75t_R g3838 ( 
.A(n_3704),
.B(n_135),
.Y(n_3838)
);

INVx5_ASAP7_75t_L g3839 ( 
.A(n_3739),
.Y(n_3839)
);

OR2x2_ASAP7_75t_L g3840 ( 
.A(n_3752),
.B(n_3666),
.Y(n_3840)
);

AND2x2_ASAP7_75t_L g3841 ( 
.A(n_3721),
.B(n_3729),
.Y(n_3841)
);

AND2x4_ASAP7_75t_SL g3842 ( 
.A(n_3742),
.B(n_3733),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_3709),
.B(n_3675),
.Y(n_3843)
);

HB1xp67_ASAP7_75t_L g3844 ( 
.A(n_3725),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3731),
.B(n_3619),
.Y(n_3845)
);

HB1xp67_ASAP7_75t_L g3846 ( 
.A(n_3773),
.Y(n_3846)
);

INVx1_ASAP7_75t_SL g3847 ( 
.A(n_3730),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3780),
.Y(n_3848)
);

AND2x2_ASAP7_75t_L g3849 ( 
.A(n_3740),
.B(n_3677),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3780),
.Y(n_3850)
);

OR2x2_ASAP7_75t_L g3851 ( 
.A(n_3746),
.B(n_3677),
.Y(n_3851)
);

INVxp67_ASAP7_75t_SL g3852 ( 
.A(n_3728),
.Y(n_3852)
);

BUFx2_ASAP7_75t_L g3853 ( 
.A(n_3737),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3755),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_3714),
.B(n_3619),
.Y(n_3855)
);

OR2x2_ASAP7_75t_L g3856 ( 
.A(n_3710),
.B(n_3688),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3760),
.B(n_3691),
.Y(n_3857)
);

OR2x2_ASAP7_75t_L g3858 ( 
.A(n_3743),
.B(n_3220),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_3751),
.Y(n_3859)
);

INVx2_ASAP7_75t_L g3860 ( 
.A(n_3749),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3727),
.B(n_3220),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3792),
.Y(n_3862)
);

BUFx2_ASAP7_75t_L g3863 ( 
.A(n_3793),
.Y(n_3863)
);

AOI32xp33_ASAP7_75t_L g3864 ( 
.A1(n_3770),
.A2(n_3703),
.A3(n_3769),
.B1(n_3712),
.B2(n_3744),
.Y(n_3864)
);

AND2x4_ASAP7_75t_L g3865 ( 
.A(n_3793),
.B(n_3221),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3792),
.Y(n_3866)
);

HB1xp67_ASAP7_75t_L g3867 ( 
.A(n_3756),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3713),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3712),
.B(n_3221),
.Y(n_3869)
);

NOR3xp33_ASAP7_75t_SL g3870 ( 
.A(n_3734),
.B(n_3741),
.C(n_3747),
.Y(n_3870)
);

INVx4_ASAP7_75t_L g3871 ( 
.A(n_3758),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3783),
.Y(n_3872)
);

AND2x2_ASAP7_75t_L g3873 ( 
.A(n_3754),
.B(n_3228),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3757),
.Y(n_3874)
);

AND2x4_ASAP7_75t_L g3875 ( 
.A(n_3788),
.B(n_3190),
.Y(n_3875)
);

BUFx3_ASAP7_75t_L g3876 ( 
.A(n_3782),
.Y(n_3876)
);

AOI33xp33_ASAP7_75t_L g3877 ( 
.A1(n_3743),
.A2(n_3218),
.A3(n_137),
.B1(n_138),
.B2(n_139),
.B3(n_140),
.Y(n_3877)
);

AOI33xp33_ASAP7_75t_L g3878 ( 
.A1(n_3736),
.A2(n_136),
.A3(n_140),
.B1(n_141),
.B2(n_142),
.B3(n_144),
.Y(n_3878)
);

AND2x2_ASAP7_75t_L g3879 ( 
.A(n_3791),
.B(n_3228),
.Y(n_3879)
);

HB1xp67_ASAP7_75t_L g3880 ( 
.A(n_3705),
.Y(n_3880)
);

AND2x2_ASAP7_75t_L g3881 ( 
.A(n_3794),
.B(n_3179),
.Y(n_3881)
);

INVx2_ASAP7_75t_L g3882 ( 
.A(n_3753),
.Y(n_3882)
);

OAI31xp33_ASAP7_75t_L g3883 ( 
.A1(n_3765),
.A2(n_3224),
.A3(n_3190),
.B(n_3223),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_3705),
.B(n_3179),
.Y(n_3884)
);

OR2x2_ASAP7_75t_L g3885 ( 
.A(n_3736),
.B(n_3223),
.Y(n_3885)
);

NAND3xp33_ASAP7_75t_L g3886 ( 
.A(n_3744),
.B(n_3763),
.C(n_3766),
.Y(n_3886)
);

INVx1_ASAP7_75t_SL g3887 ( 
.A(n_3805),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3812),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_3809),
.B(n_3777),
.Y(n_3889)
);

NAND2x1p5_ASAP7_75t_L g3890 ( 
.A(n_3809),
.B(n_3779),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_L g3891 ( 
.A(n_3803),
.B(n_3778),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3812),
.Y(n_3892)
);

AOI22xp5_ASAP7_75t_L g3893 ( 
.A1(n_3831),
.A2(n_3790),
.B1(n_3784),
.B2(n_3766),
.Y(n_3893)
);

AOI22xp5_ASAP7_75t_L g3894 ( 
.A1(n_3831),
.A2(n_3790),
.B1(n_3784),
.B2(n_3787),
.Y(n_3894)
);

INVx2_ASAP7_75t_L g3895 ( 
.A(n_3805),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_L g3896 ( 
.A(n_3802),
.B(n_3789),
.Y(n_3896)
);

OAI22xp5_ASAP7_75t_L g3897 ( 
.A1(n_3799),
.A2(n_3852),
.B1(n_3880),
.B2(n_3886),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3846),
.Y(n_3898)
);

OAI33xp33_ASAP7_75t_L g3899 ( 
.A1(n_3837),
.A2(n_3798),
.A3(n_3868),
.B1(n_3808),
.B2(n_3855),
.B3(n_3845),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3846),
.Y(n_3900)
);

INVx2_ASAP7_75t_L g3901 ( 
.A(n_3805),
.Y(n_3901)
);

AO22x1_ASAP7_75t_L g3902 ( 
.A1(n_3852),
.A2(n_3814),
.B1(n_3880),
.B2(n_3844),
.Y(n_3902)
);

BUFx2_ASAP7_75t_L g3903 ( 
.A(n_3801),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3814),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3814),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3814),
.Y(n_3906)
);

INVx2_ASAP7_75t_L g3907 ( 
.A(n_3863),
.Y(n_3907)
);

OAI32xp33_ASAP7_75t_L g3908 ( 
.A1(n_3867),
.A2(n_3219),
.A3(n_3216),
.B1(n_3664),
.B2(n_3647),
.Y(n_3908)
);

AND2x2_ASAP7_75t_L g3909 ( 
.A(n_3801),
.B(n_3647),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3808),
.Y(n_3910)
);

NAND3xp33_ASAP7_75t_L g3911 ( 
.A(n_3864),
.B(n_3664),
.C(n_3647),
.Y(n_3911)
);

INVx2_ASAP7_75t_L g3912 ( 
.A(n_3839),
.Y(n_3912)
);

AOI22xp5_ASAP7_75t_L g3913 ( 
.A1(n_3799),
.A2(n_3664),
.B1(n_3428),
.B2(n_3224),
.Y(n_3913)
);

NOR2xp33_ASAP7_75t_L g3914 ( 
.A(n_3828),
.B(n_3216),
.Y(n_3914)
);

OAI21xp5_ASAP7_75t_L g3915 ( 
.A1(n_3837),
.A2(n_3219),
.B(n_3216),
.Y(n_3915)
);

OAI211xp5_ASAP7_75t_L g3916 ( 
.A1(n_3870),
.A2(n_3219),
.B(n_141),
.C(n_142),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_L g3917 ( 
.A(n_3841),
.B(n_136),
.Y(n_3917)
);

HB1xp67_ASAP7_75t_L g3918 ( 
.A(n_3811),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3859),
.Y(n_3919)
);

NOR2x1_ASAP7_75t_L g3920 ( 
.A(n_3811),
.B(n_145),
.Y(n_3920)
);

OR2x2_ASAP7_75t_L g3921 ( 
.A(n_3804),
.B(n_3847),
.Y(n_3921)
);

INVx2_ASAP7_75t_SL g3922 ( 
.A(n_3839),
.Y(n_3922)
);

INVxp67_ASAP7_75t_L g3923 ( 
.A(n_3853),
.Y(n_3923)
);

NOR2xp33_ASAP7_75t_L g3924 ( 
.A(n_3796),
.B(n_145),
.Y(n_3924)
);

NAND2x1_ASAP7_75t_L g3925 ( 
.A(n_3824),
.B(n_146),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_3839),
.Y(n_3926)
);

NAND3xp33_ASAP7_75t_L g3927 ( 
.A(n_3818),
.B(n_147),
.C(n_148),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3859),
.Y(n_3928)
);

INVx2_ASAP7_75t_L g3929 ( 
.A(n_3839),
.Y(n_3929)
);

OR2x2_ASAP7_75t_L g3930 ( 
.A(n_3874),
.B(n_3813),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_L g3931 ( 
.A(n_3877),
.B(n_147),
.Y(n_3931)
);

AOI22xp5_ASAP7_75t_L g3932 ( 
.A1(n_3825),
.A2(n_3428),
.B1(n_2868),
.B2(n_2865),
.Y(n_3932)
);

INVx2_ASAP7_75t_L g3933 ( 
.A(n_3871),
.Y(n_3933)
);

OAI33xp33_ASAP7_75t_L g3934 ( 
.A1(n_3834),
.A2(n_148),
.A3(n_149),
.B1(n_150),
.B2(n_151),
.B3(n_152),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3827),
.Y(n_3935)
);

NOR2xp67_ASAP7_75t_SL g3936 ( 
.A(n_3867),
.B(n_149),
.Y(n_3936)
);

HB1xp67_ASAP7_75t_L g3937 ( 
.A(n_3835),
.Y(n_3937)
);

INVx2_ASAP7_75t_L g3938 ( 
.A(n_3871),
.Y(n_3938)
);

OA222x2_ASAP7_75t_L g3939 ( 
.A1(n_3835),
.A2(n_150),
.B1(n_152),
.B2(n_154),
.C1(n_155),
.C2(n_156),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3836),
.Y(n_3940)
);

INVx2_ASAP7_75t_SL g3941 ( 
.A(n_3815),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3877),
.B(n_154),
.Y(n_3942)
);

NOR2xp33_ASAP7_75t_L g3943 ( 
.A(n_3854),
.B(n_3842),
.Y(n_3943)
);

INVx1_ASAP7_75t_SL g3944 ( 
.A(n_3838),
.Y(n_3944)
);

OR2x2_ASAP7_75t_L g3945 ( 
.A(n_3807),
.B(n_156),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3820),
.Y(n_3946)
);

AND2x2_ASAP7_75t_L g3947 ( 
.A(n_3842),
.B(n_157),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3820),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3830),
.Y(n_3949)
);

OAI222xp33_ASAP7_75t_L g3950 ( 
.A1(n_3844),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.C1(n_161),
.C2(n_162),
.Y(n_3950)
);

OR2x6_ASAP7_75t_L g3951 ( 
.A(n_3860),
.B(n_160),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3860),
.B(n_161),
.Y(n_3952)
);

OAI211xp5_ASAP7_75t_L g3953 ( 
.A1(n_3870),
.A2(n_162),
.B(n_163),
.C(n_164),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3830),
.Y(n_3954)
);

AND2x4_ASAP7_75t_L g3955 ( 
.A(n_3815),
.B(n_163),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3817),
.B(n_165),
.Y(n_3956)
);

AND2x2_ASAP7_75t_L g3957 ( 
.A(n_3876),
.B(n_169),
.Y(n_3957)
);

AOI22xp5_ASAP7_75t_L g3958 ( 
.A1(n_3825),
.A2(n_3806),
.B1(n_3829),
.B2(n_3832),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3840),
.Y(n_3959)
);

INVx2_ASAP7_75t_L g3960 ( 
.A(n_3876),
.Y(n_3960)
);

XOR2xp5_ASAP7_75t_L g3961 ( 
.A(n_3843),
.B(n_170),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3851),
.Y(n_3962)
);

AND2x4_ASAP7_75t_L g3963 ( 
.A(n_3821),
.B(n_171),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3833),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3856),
.Y(n_3965)
);

A2O1A1Ixp33_ASAP7_75t_L g3966 ( 
.A1(n_3818),
.A2(n_172),
.B(n_175),
.C(n_176),
.Y(n_3966)
);

AND2x2_ASAP7_75t_L g3967 ( 
.A(n_3800),
.B(n_172),
.Y(n_3967)
);

NAND4xp75_ASAP7_75t_L g3968 ( 
.A(n_3882),
.B(n_176),
.C(n_178),
.D(n_180),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3816),
.Y(n_3969)
);

NOR2xp33_ASAP7_75t_L g3970 ( 
.A(n_3797),
.B(n_178),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3819),
.Y(n_3971)
);

AND2x4_ASAP7_75t_L g3972 ( 
.A(n_3822),
.B(n_182),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3823),
.Y(n_3973)
);

AOI22xp5_ASAP7_75t_L g3974 ( 
.A1(n_3795),
.A2(n_2850),
.B1(n_184),
.B2(n_185),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3826),
.Y(n_3975)
);

INVx2_ASAP7_75t_L g3976 ( 
.A(n_3918),
.Y(n_3976)
);

AOI21xp33_ASAP7_75t_SL g3977 ( 
.A1(n_3927),
.A2(n_3897),
.B(n_3958),
.Y(n_3977)
);

INVxp67_ASAP7_75t_L g3978 ( 
.A(n_3903),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3898),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3900),
.Y(n_3980)
);

AOI21xp33_ASAP7_75t_L g3981 ( 
.A1(n_3958),
.A2(n_3882),
.B(n_3810),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3937),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3921),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_3944),
.B(n_3878),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3920),
.Y(n_3985)
);

AND2x2_ASAP7_75t_L g3986 ( 
.A(n_3941),
.B(n_3849),
.Y(n_3986)
);

AND2x2_ASAP7_75t_L g3987 ( 
.A(n_3887),
.B(n_3872),
.Y(n_3987)
);

NOR2xp33_ASAP7_75t_R g3988 ( 
.A(n_3947),
.B(n_3838),
.Y(n_3988)
);

AOI22xp5_ASAP7_75t_L g3989 ( 
.A1(n_3899),
.A2(n_3861),
.B1(n_3869),
.B2(n_3857),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3920),
.Y(n_3990)
);

AND2x2_ASAP7_75t_L g3991 ( 
.A(n_3907),
.B(n_3848),
.Y(n_3991)
);

CKINVDCx5p33_ASAP7_75t_R g3992 ( 
.A(n_3951),
.Y(n_3992)
);

INVx5_ASAP7_75t_L g3993 ( 
.A(n_3951),
.Y(n_3993)
);

AND2x2_ASAP7_75t_L g3994 ( 
.A(n_3890),
.B(n_3850),
.Y(n_3994)
);

INVxp67_ASAP7_75t_SL g3995 ( 
.A(n_3902),
.Y(n_3995)
);

AOI221xp5_ASAP7_75t_L g3996 ( 
.A1(n_3966),
.A2(n_3884),
.B1(n_3883),
.B2(n_3862),
.C(n_3866),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_L g3997 ( 
.A(n_3895),
.B(n_3878),
.Y(n_3997)
);

NOR3xp33_ASAP7_75t_L g3998 ( 
.A(n_3953),
.B(n_3858),
.C(n_3885),
.Y(n_3998)
);

AOI21xp5_ASAP7_75t_L g3999 ( 
.A1(n_3916),
.A2(n_3865),
.B(n_3875),
.Y(n_3999)
);

AND2x2_ASAP7_75t_L g4000 ( 
.A(n_3901),
.B(n_3875),
.Y(n_4000)
);

AOI22xp5_ASAP7_75t_L g4001 ( 
.A1(n_3893),
.A2(n_3894),
.B1(n_3943),
.B2(n_3961),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3955),
.B(n_3865),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3904),
.Y(n_4003)
);

AND2x2_ASAP7_75t_L g4004 ( 
.A(n_3960),
.B(n_3873),
.Y(n_4004)
);

OR2x6_ASAP7_75t_L g4005 ( 
.A(n_3933),
.B(n_3881),
.Y(n_4005)
);

INVx1_ASAP7_75t_SL g4006 ( 
.A(n_3955),
.Y(n_4006)
);

INVx1_ASAP7_75t_SL g4007 ( 
.A(n_3930),
.Y(n_4007)
);

OR2x2_ASAP7_75t_L g4008 ( 
.A(n_3923),
.B(n_3959),
.Y(n_4008)
);

OR2x2_ASAP7_75t_L g4009 ( 
.A(n_3889),
.B(n_3879),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_SL g4010 ( 
.A(n_3893),
.B(n_183),
.Y(n_4010)
);

INVx2_ASAP7_75t_SL g4011 ( 
.A(n_3922),
.Y(n_4011)
);

AND2x4_ASAP7_75t_L g4012 ( 
.A(n_3912),
.B(n_185),
.Y(n_4012)
);

INVx2_ASAP7_75t_L g4013 ( 
.A(n_3888),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3905),
.Y(n_4014)
);

INVx1_ASAP7_75t_SL g4015 ( 
.A(n_3957),
.Y(n_4015)
);

AND2x2_ASAP7_75t_L g4016 ( 
.A(n_3967),
.B(n_186),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3906),
.Y(n_4017)
);

BUFx2_ASAP7_75t_L g4018 ( 
.A(n_3938),
.Y(n_4018)
);

AND2x4_ASAP7_75t_L g4019 ( 
.A(n_3926),
.B(n_187),
.Y(n_4019)
);

AND2x2_ASAP7_75t_L g4020 ( 
.A(n_3962),
.B(n_188),
.Y(n_4020)
);

INVx2_ASAP7_75t_L g4021 ( 
.A(n_3892),
.Y(n_4021)
);

AND2x2_ASAP7_75t_L g4022 ( 
.A(n_3964),
.B(n_189),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_3936),
.B(n_189),
.Y(n_4023)
);

AND2x2_ASAP7_75t_L g4024 ( 
.A(n_3965),
.B(n_190),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_L g4025 ( 
.A(n_3963),
.B(n_190),
.Y(n_4025)
);

CKINVDCx16_ASAP7_75t_R g4026 ( 
.A(n_3963),
.Y(n_4026)
);

AND2x2_ASAP7_75t_L g4027 ( 
.A(n_3891),
.B(n_191),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_L g4028 ( 
.A(n_3925),
.B(n_3968),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3929),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_3970),
.B(n_191),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_3946),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3924),
.B(n_192),
.Y(n_4032)
);

INVx2_ASAP7_75t_L g4033 ( 
.A(n_3910),
.Y(n_4033)
);

INVx2_ASAP7_75t_L g4034 ( 
.A(n_3909),
.Y(n_4034)
);

OAI31xp33_ASAP7_75t_L g4035 ( 
.A1(n_3950),
.A2(n_192),
.A3(n_193),
.B(n_195),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3917),
.B(n_193),
.Y(n_4036)
);

NOR3xp33_ASAP7_75t_SL g4037 ( 
.A(n_3935),
.B(n_195),
.C(n_196),
.Y(n_4037)
);

INVx3_ASAP7_75t_L g4038 ( 
.A(n_3972),
.Y(n_4038)
);

INVx2_ASAP7_75t_L g4039 ( 
.A(n_3972),
.Y(n_4039)
);

INVx3_ASAP7_75t_L g4040 ( 
.A(n_3919),
.Y(n_4040)
);

INVx1_ASAP7_75t_SL g4041 ( 
.A(n_3945),
.Y(n_4041)
);

AND2x2_ASAP7_75t_L g4042 ( 
.A(n_3940),
.B(n_196),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_3931),
.B(n_198),
.Y(n_4043)
);

INVx2_ASAP7_75t_L g4044 ( 
.A(n_3948),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_L g4045 ( 
.A(n_3942),
.B(n_198),
.Y(n_4045)
);

AND2x2_ASAP7_75t_L g4046 ( 
.A(n_3914),
.B(n_199),
.Y(n_4046)
);

AO21x2_ASAP7_75t_L g4047 ( 
.A1(n_3952),
.A2(n_3911),
.B(n_3894),
.Y(n_4047)
);

NOR2x1_ASAP7_75t_L g4048 ( 
.A(n_3928),
.B(n_199),
.Y(n_4048)
);

BUFx2_ASAP7_75t_L g4049 ( 
.A(n_3956),
.Y(n_4049)
);

AND2x2_ASAP7_75t_L g4050 ( 
.A(n_3896),
.B(n_200),
.Y(n_4050)
);

AND2x2_ASAP7_75t_L g4051 ( 
.A(n_3939),
.B(n_3949),
.Y(n_4051)
);

AND2x2_ASAP7_75t_L g4052 ( 
.A(n_3954),
.B(n_200),
.Y(n_4052)
);

AND2x4_ASAP7_75t_L g4053 ( 
.A(n_3969),
.B(n_201),
.Y(n_4053)
);

HB1xp67_ASAP7_75t_L g4054 ( 
.A(n_3971),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3973),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3975),
.Y(n_4056)
);

NAND2xp33_ASAP7_75t_R g4057 ( 
.A(n_3939),
.B(n_201),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3915),
.Y(n_4058)
);

OR2x2_ASAP7_75t_L g4059 ( 
.A(n_4026),
.B(n_3974),
.Y(n_4059)
);

AOI22xp5_ASAP7_75t_L g4060 ( 
.A1(n_4010),
.A2(n_3998),
.B1(n_4001),
.B2(n_4047),
.Y(n_4060)
);

AND2x2_ASAP7_75t_L g4061 ( 
.A(n_3986),
.B(n_3974),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_L g4062 ( 
.A(n_3993),
.B(n_3995),
.Y(n_4062)
);

OAI21xp33_ASAP7_75t_L g4063 ( 
.A1(n_3977),
.A2(n_3932),
.B(n_3913),
.Y(n_4063)
);

OAI22xp5_ASAP7_75t_L g4064 ( 
.A1(n_3995),
.A2(n_3913),
.B1(n_3934),
.B2(n_3908),
.Y(n_4064)
);

AOI22xp33_ASAP7_75t_L g4065 ( 
.A1(n_3998),
.A2(n_2786),
.B1(n_2804),
.B2(n_1048),
.Y(n_4065)
);

AND2x2_ASAP7_75t_L g4066 ( 
.A(n_4006),
.B(n_202),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3993),
.B(n_202),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_L g4068 ( 
.A(n_3992),
.B(n_203),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3993),
.Y(n_4069)
);

AND3x2_ASAP7_75t_L g4070 ( 
.A(n_3978),
.B(n_203),
.C(n_204),
.Y(n_4070)
);

INVx1_ASAP7_75t_SL g4071 ( 
.A(n_3988),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_3992),
.B(n_205),
.Y(n_4072)
);

OR2x2_ASAP7_75t_L g4073 ( 
.A(n_4039),
.B(n_4007),
.Y(n_4073)
);

NOR3xp33_ASAP7_75t_SL g4074 ( 
.A(n_4010),
.B(n_206),
.C(n_207),
.Y(n_4074)
);

INVx2_ASAP7_75t_L g4075 ( 
.A(n_3993),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_4040),
.Y(n_4076)
);

INVx1_ASAP7_75t_SL g4077 ( 
.A(n_3988),
.Y(n_4077)
);

AND2x2_ASAP7_75t_L g4078 ( 
.A(n_3987),
.B(n_4004),
.Y(n_4078)
);

OAI211xp5_ASAP7_75t_L g4079 ( 
.A1(n_3989),
.A2(n_206),
.B(n_207),
.C(n_208),
.Y(n_4079)
);

AND3x1_ASAP7_75t_L g4080 ( 
.A(n_4035),
.B(n_4037),
.C(n_4028),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_4040),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_4038),
.B(n_208),
.Y(n_4082)
);

HB1xp67_ASAP7_75t_L g4083 ( 
.A(n_3978),
.Y(n_4083)
);

NOR2xp33_ASAP7_75t_L g4084 ( 
.A(n_4015),
.B(n_209),
.Y(n_4084)
);

OR2x2_ASAP7_75t_L g4085 ( 
.A(n_4039),
.B(n_210),
.Y(n_4085)
);

INVxp67_ASAP7_75t_L g4086 ( 
.A(n_4057),
.Y(n_4086)
);

OAI21xp33_ASAP7_75t_L g4087 ( 
.A1(n_3984),
.A2(n_210),
.B(n_211),
.Y(n_4087)
);

NAND2xp5_ASAP7_75t_L g4088 ( 
.A(n_4038),
.B(n_212),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_4040),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_3985),
.B(n_212),
.Y(n_4090)
);

AND3x2_ASAP7_75t_L g4091 ( 
.A(n_3990),
.B(n_213),
.C(n_214),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_4048),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_4034),
.B(n_214),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_4038),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_4034),
.B(n_215),
.Y(n_4095)
);

AND2x2_ASAP7_75t_L g4096 ( 
.A(n_3983),
.B(n_216),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_4029),
.Y(n_4097)
);

NAND2xp67_ASAP7_75t_L g4098 ( 
.A(n_4052),
.B(n_216),
.Y(n_4098)
);

AND2x2_ASAP7_75t_L g4099 ( 
.A(n_4000),
.B(n_4018),
.Y(n_4099)
);

AND5x1_ASAP7_75t_L g4100 ( 
.A(n_3996),
.B(n_217),
.C(n_218),
.D(n_219),
.E(n_221),
.Y(n_4100)
);

NAND2xp33_ASAP7_75t_L g4101 ( 
.A(n_4037),
.B(n_4051),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_4011),
.B(n_217),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_4000),
.B(n_221),
.Y(n_4103)
);

INVx2_ASAP7_75t_L g4104 ( 
.A(n_4011),
.Y(n_4104)
);

INVx3_ASAP7_75t_L g4105 ( 
.A(n_4012),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_L g4106 ( 
.A(n_4047),
.B(n_222),
.Y(n_4106)
);

HB1xp67_ASAP7_75t_L g4107 ( 
.A(n_4005),
.Y(n_4107)
);

AND2x4_ASAP7_75t_L g4108 ( 
.A(n_3982),
.B(n_223),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_3999),
.B(n_223),
.Y(n_4109)
);

OR2x2_ASAP7_75t_L g4110 ( 
.A(n_3997),
.B(n_224),
.Y(n_4110)
);

NOR2xp33_ASAP7_75t_L g4111 ( 
.A(n_4041),
.B(n_224),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_4029),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_4012),
.Y(n_4113)
);

NAND2xp67_ASAP7_75t_SL g4114 ( 
.A(n_3994),
.B(n_4052),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_4022),
.B(n_225),
.Y(n_4115)
);

OAI21xp33_ASAP7_75t_SL g4116 ( 
.A1(n_3981),
.A2(n_225),
.B(n_226),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_SL g4117 ( 
.A(n_4002),
.B(n_227),
.Y(n_4117)
);

INVx3_ASAP7_75t_L g4118 ( 
.A(n_4012),
.Y(n_4118)
);

OR2x2_ASAP7_75t_L g4119 ( 
.A(n_4008),
.B(n_227),
.Y(n_4119)
);

HB1xp67_ASAP7_75t_L g4120 ( 
.A(n_4005),
.Y(n_4120)
);

AND2x2_ASAP7_75t_L g4121 ( 
.A(n_4027),
.B(n_228),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_4019),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_4019),
.Y(n_4123)
);

AOI21xp33_ASAP7_75t_L g4124 ( 
.A1(n_4086),
.A2(n_4057),
.B(n_4009),
.Y(n_4124)
);

OR2x2_ASAP7_75t_L g4125 ( 
.A(n_4105),
.B(n_4005),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_4105),
.Y(n_4126)
);

AOI22xp5_ASAP7_75t_L g4127 ( 
.A1(n_4060),
.A2(n_4050),
.B1(n_3991),
.B2(n_4049),
.Y(n_4127)
);

AOI22xp33_ASAP7_75t_SL g4128 ( 
.A1(n_4079),
.A2(n_4058),
.B1(n_4054),
.B2(n_3976),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_L g4129 ( 
.A(n_4099),
.B(n_4022),
.Y(n_4129)
);

AOI221xp5_ASAP7_75t_L g4130 ( 
.A1(n_4064),
.A2(n_3979),
.B1(n_3980),
.B2(n_4054),
.C(n_3976),
.Y(n_4130)
);

AOI221xp5_ASAP7_75t_L g4131 ( 
.A1(n_4064),
.A2(n_4033),
.B1(n_4013),
.B2(n_4021),
.C(n_4017),
.Y(n_4131)
);

OAI322xp33_ASAP7_75t_L g4132 ( 
.A1(n_4106),
.A2(n_4033),
.A3(n_4013),
.B1(n_4021),
.B2(n_4056),
.C1(n_4055),
.C2(n_4031),
.Y(n_4132)
);

INVx2_ASAP7_75t_L g4133 ( 
.A(n_4118),
.Y(n_4133)
);

AOI31xp33_ASAP7_75t_L g4134 ( 
.A1(n_4107),
.A2(n_4003),
.A3(n_4014),
.B(n_4044),
.Y(n_4134)
);

A2O1A1Ixp33_ASAP7_75t_L g4135 ( 
.A1(n_4106),
.A2(n_4045),
.B(n_4043),
.C(n_4042),
.Y(n_4135)
);

OAI211xp5_ASAP7_75t_SL g4136 ( 
.A1(n_4063),
.A2(n_4044),
.B(n_4030),
.C(n_4032),
.Y(n_4136)
);

AOI21xp5_ASAP7_75t_L g4137 ( 
.A1(n_4101),
.A2(n_4023),
.B(n_4020),
.Y(n_4137)
);

OAI31xp33_ASAP7_75t_L g4138 ( 
.A1(n_4092),
.A2(n_4042),
.A3(n_4024),
.B(n_4019),
.Y(n_4138)
);

AOI211xp5_ASAP7_75t_SL g4139 ( 
.A1(n_4120),
.A2(n_4046),
.B(n_4025),
.C(n_4036),
.Y(n_4139)
);

AOI22xp33_ASAP7_75t_SL g4140 ( 
.A1(n_4078),
.A2(n_4016),
.B1(n_4053),
.B2(n_232),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_4118),
.Y(n_4141)
);

AND2x2_ASAP7_75t_SL g4142 ( 
.A(n_4080),
.B(n_4053),
.Y(n_4142)
);

OAI21xp5_ASAP7_75t_L g4143 ( 
.A1(n_4116),
.A2(n_4053),
.B(n_230),
.Y(n_4143)
);

AO22x1_ASAP7_75t_L g4144 ( 
.A1(n_4113),
.A2(n_229),
.B1(n_230),
.B2(n_233),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_4062),
.Y(n_4145)
);

INVx2_ASAP7_75t_L g4146 ( 
.A(n_4122),
.Y(n_4146)
);

INVx2_ASAP7_75t_L g4147 ( 
.A(n_4123),
.Y(n_4147)
);

NOR2xp33_ASAP7_75t_L g4148 ( 
.A(n_4071),
.B(n_229),
.Y(n_4148)
);

OAI22xp33_ASAP7_75t_L g4149 ( 
.A1(n_4109),
.A2(n_234),
.B1(n_235),
.B2(n_237),
.Y(n_4149)
);

AOI211xp5_ASAP7_75t_L g4150 ( 
.A1(n_4062),
.A2(n_234),
.B(n_235),
.C(n_237),
.Y(n_4150)
);

O2A1O1Ixp33_ASAP7_75t_L g4151 ( 
.A1(n_4083),
.A2(n_238),
.B(n_240),
.C(n_241),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_4070),
.B(n_240),
.Y(n_4152)
);

INVx2_ASAP7_75t_L g4153 ( 
.A(n_4076),
.Y(n_4153)
);

OAI32xp33_ASAP7_75t_L g4154 ( 
.A1(n_4059),
.A2(n_242),
.A3(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_4154)
);

NOR2xp33_ASAP7_75t_L g4155 ( 
.A(n_4071),
.B(n_4077),
.Y(n_4155)
);

INVx1_ASAP7_75t_SL g4156 ( 
.A(n_4073),
.Y(n_4156)
);

INVx2_ASAP7_75t_SL g4157 ( 
.A(n_4104),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_4091),
.B(n_244),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_L g4159 ( 
.A(n_4077),
.B(n_246),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_4094),
.B(n_247),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_4098),
.B(n_248),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4081),
.Y(n_4162)
);

OAI221xp5_ASAP7_75t_L g4163 ( 
.A1(n_4100),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.C(n_252),
.Y(n_4163)
);

AOI22xp5_ASAP7_75t_L g4164 ( 
.A1(n_4061),
.A2(n_250),
.B1(n_253),
.B2(n_255),
.Y(n_4164)
);

XNOR2x1_ASAP7_75t_L g4165 ( 
.A(n_4110),
.B(n_253),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_4089),
.Y(n_4166)
);

AOI21xp33_ASAP7_75t_L g4167 ( 
.A1(n_4069),
.A2(n_255),
.B(n_256),
.Y(n_4167)
);

AOI211xp5_ASAP7_75t_SL g4168 ( 
.A1(n_4097),
.A2(n_4112),
.B(n_4067),
.C(n_4111),
.Y(n_4168)
);

NOR2xp33_ASAP7_75t_L g4169 ( 
.A(n_4087),
.B(n_257),
.Y(n_4169)
);

AND2x2_ASAP7_75t_L g4170 ( 
.A(n_4066),
.B(n_257),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_4067),
.Y(n_4171)
);

OAI22xp33_ASAP7_75t_L g4172 ( 
.A1(n_4068),
.A2(n_258),
.B1(n_259),
.B2(n_262),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4075),
.Y(n_4173)
);

NAND2xp5_ASAP7_75t_L g4174 ( 
.A(n_4103),
.B(n_258),
.Y(n_4174)
);

OR2x2_ASAP7_75t_L g4175 ( 
.A(n_4072),
.B(n_4119),
.Y(n_4175)
);

BUFx2_ASAP7_75t_L g4176 ( 
.A(n_4114),
.Y(n_4176)
);

AOI21xp33_ASAP7_75t_L g4177 ( 
.A1(n_4082),
.A2(n_259),
.B(n_262),
.Y(n_4177)
);

OAI21xp33_ASAP7_75t_L g4178 ( 
.A1(n_4074),
.A2(n_263),
.B(n_264),
.Y(n_4178)
);

A2O1A1Ixp33_ASAP7_75t_L g4179 ( 
.A1(n_4084),
.A2(n_263),
.B(n_264),
.C(n_265),
.Y(n_4179)
);

AOI21xp5_ASAP7_75t_L g4180 ( 
.A1(n_4090),
.A2(n_4117),
.B(n_4088),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_4102),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_4085),
.Y(n_4182)
);

NAND3xp33_ASAP7_75t_SL g4183 ( 
.A(n_4096),
.B(n_266),
.C(n_268),
.Y(n_4183)
);

AND2x2_ASAP7_75t_L g4184 ( 
.A(n_4142),
.B(n_4121),
.Y(n_4184)
);

OR2x2_ASAP7_75t_L g4185 ( 
.A(n_4125),
.B(n_4093),
.Y(n_4185)
);

INVx2_ASAP7_75t_L g4186 ( 
.A(n_4133),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4129),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4126),
.Y(n_4188)
);

OR2x6_ASAP7_75t_L g4189 ( 
.A(n_4141),
.B(n_4090),
.Y(n_4189)
);

INVx1_ASAP7_75t_SL g4190 ( 
.A(n_4156),
.Y(n_4190)
);

AOI31xp33_ASAP7_75t_L g4191 ( 
.A1(n_4140),
.A2(n_4095),
.A3(n_4093),
.B(n_4115),
.Y(n_4191)
);

INVx2_ASAP7_75t_L g4192 ( 
.A(n_4146),
.Y(n_4192)
);

HB1xp67_ASAP7_75t_L g4193 ( 
.A(n_4156),
.Y(n_4193)
);

NAND2xp5_ASAP7_75t_L g4194 ( 
.A(n_4144),
.B(n_4108),
.Y(n_4194)
);

INVx2_ASAP7_75t_SL g4195 ( 
.A(n_4147),
.Y(n_4195)
);

AOI221xp5_ASAP7_75t_L g4196 ( 
.A1(n_4130),
.A2(n_4065),
.B1(n_4095),
.B2(n_4108),
.C(n_271),
.Y(n_4196)
);

AND2x2_ASAP7_75t_L g4197 ( 
.A(n_4157),
.B(n_266),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_4138),
.B(n_4176),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4170),
.Y(n_4199)
);

NAND2x1p5_ASAP7_75t_L g4200 ( 
.A(n_4145),
.B(n_268),
.Y(n_4200)
);

AND2x2_ASAP7_75t_L g4201 ( 
.A(n_4139),
.B(n_4155),
.Y(n_4201)
);

OAI21xp5_ASAP7_75t_SL g4202 ( 
.A1(n_4128),
.A2(n_270),
.B(n_271),
.Y(n_4202)
);

OR2x2_ASAP7_75t_L g4203 ( 
.A(n_4159),
.B(n_270),
.Y(n_4203)
);

OAI22xp5_ASAP7_75t_L g4204 ( 
.A1(n_4127),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_4204)
);

AOI21xp33_ASAP7_75t_SL g4205 ( 
.A1(n_4138),
.A2(n_272),
.B(n_273),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_4158),
.Y(n_4206)
);

NOR2xp33_ASAP7_75t_L g4207 ( 
.A(n_4124),
.B(n_274),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4161),
.Y(n_4208)
);

AOI31xp33_ASAP7_75t_L g4209 ( 
.A1(n_4143),
.A2(n_275),
.A3(n_276),
.B(n_277),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_4134),
.Y(n_4210)
);

NAND2x1p5_ASAP7_75t_L g4211 ( 
.A(n_4182),
.B(n_275),
.Y(n_4211)
);

INVx2_ASAP7_75t_L g4212 ( 
.A(n_4175),
.Y(n_4212)
);

AND2x4_ASAP7_75t_L g4213 ( 
.A(n_4173),
.B(n_277),
.Y(n_4213)
);

O2A1O1Ixp33_ASAP7_75t_L g4214 ( 
.A1(n_4132),
.A2(n_278),
.B(n_279),
.C(n_280),
.Y(n_4214)
);

OAI22xp33_ASAP7_75t_L g4215 ( 
.A1(n_4168),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_L g4216 ( 
.A(n_4131),
.B(n_281),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_4152),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_4174),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_L g4219 ( 
.A(n_4137),
.B(n_281),
.Y(n_4219)
);

AOI21xp5_ASAP7_75t_L g4220 ( 
.A1(n_4180),
.A2(n_283),
.B(n_284),
.Y(n_4220)
);

NOR2xp33_ASAP7_75t_L g4221 ( 
.A(n_4178),
.B(n_284),
.Y(n_4221)
);

INVxp67_ASAP7_75t_L g4222 ( 
.A(n_4148),
.Y(n_4222)
);

NOR2xp33_ASAP7_75t_L g4223 ( 
.A(n_4163),
.B(n_285),
.Y(n_4223)
);

NAND2xp5_ASAP7_75t_L g4224 ( 
.A(n_4150),
.B(n_286),
.Y(n_4224)
);

INVx2_ASAP7_75t_L g4225 ( 
.A(n_4153),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4171),
.Y(n_4226)
);

BUFx2_ASAP7_75t_SL g4227 ( 
.A(n_4162),
.Y(n_4227)
);

INVx1_ASAP7_75t_SL g4228 ( 
.A(n_4165),
.Y(n_4228)
);

HB1xp67_ASAP7_75t_L g4229 ( 
.A(n_4166),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_SL g4230 ( 
.A(n_4149),
.B(n_286),
.Y(n_4230)
);

OAI322xp33_ASAP7_75t_L g4231 ( 
.A1(n_4160),
.A2(n_287),
.A3(n_288),
.B1(n_293),
.B2(n_295),
.C1(n_296),
.C2(n_298),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_SL g4232 ( 
.A(n_4151),
.B(n_288),
.Y(n_4232)
);

AOI32xp33_ASAP7_75t_L g4233 ( 
.A1(n_4136),
.A2(n_293),
.A3(n_295),
.B1(n_299),
.B2(n_301),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_4193),
.Y(n_4234)
);

NOR4xp25_ASAP7_75t_SL g4235 ( 
.A(n_4202),
.B(n_4181),
.C(n_4135),
.D(n_4167),
.Y(n_4235)
);

INVx2_ASAP7_75t_L g4236 ( 
.A(n_4211),
.Y(n_4236)
);

AND2x2_ASAP7_75t_L g4237 ( 
.A(n_4184),
.B(n_4169),
.Y(n_4237)
);

NAND3xp33_ASAP7_75t_SL g4238 ( 
.A(n_4190),
.B(n_4150),
.C(n_4164),
.Y(n_4238)
);

NAND2x1_ASAP7_75t_L g4239 ( 
.A(n_4189),
.B(n_4213),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_L g4240 ( 
.A(n_4205),
.B(n_4179),
.Y(n_4240)
);

AOI22xp5_ASAP7_75t_L g4241 ( 
.A1(n_4210),
.A2(n_4183),
.B1(n_4172),
.B2(n_4177),
.Y(n_4241)
);

NAND2xp5_ASAP7_75t_SL g4242 ( 
.A(n_4194),
.B(n_4132),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_4211),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_4200),
.Y(n_4244)
);

XOR2x2_ASAP7_75t_L g4245 ( 
.A(n_4228),
.B(n_4154),
.Y(n_4245)
);

NOR3xp33_ASAP7_75t_SL g4246 ( 
.A(n_4202),
.B(n_299),
.C(n_301),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4200),
.Y(n_4247)
);

AND2x2_ASAP7_75t_L g4248 ( 
.A(n_4201),
.B(n_4228),
.Y(n_4248)
);

OR2x2_ASAP7_75t_L g4249 ( 
.A(n_4198),
.B(n_302),
.Y(n_4249)
);

OAI22xp5_ASAP7_75t_L g4250 ( 
.A1(n_4186),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4197),
.Y(n_4251)
);

OR2x2_ASAP7_75t_L g4252 ( 
.A(n_4189),
.B(n_303),
.Y(n_4252)
);

AND2x2_ASAP7_75t_SL g4253 ( 
.A(n_4185),
.B(n_304),
.Y(n_4253)
);

NAND2xp33_ASAP7_75t_SL g4254 ( 
.A(n_4195),
.B(n_305),
.Y(n_4254)
);

AND2x2_ASAP7_75t_L g4255 ( 
.A(n_4199),
.B(n_306),
.Y(n_4255)
);

AOI31xp33_ASAP7_75t_L g4256 ( 
.A1(n_4222),
.A2(n_307),
.A3(n_308),
.B(n_310),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_SL g4257 ( 
.A(n_4215),
.B(n_308),
.Y(n_4257)
);

NOR3xp33_ASAP7_75t_SL g4258 ( 
.A(n_4216),
.B(n_310),
.C(n_311),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_4213),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_4233),
.B(n_311),
.Y(n_4260)
);

OR2x2_ASAP7_75t_L g4261 ( 
.A(n_4189),
.B(n_312),
.Y(n_4261)
);

AND2x2_ASAP7_75t_SL g4262 ( 
.A(n_4192),
.B(n_313),
.Y(n_4262)
);

OAI22xp33_ASAP7_75t_SL g4263 ( 
.A1(n_4219),
.A2(n_4224),
.B1(n_4232),
.B2(n_4188),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4229),
.Y(n_4264)
);

O2A1O1Ixp33_ASAP7_75t_L g4265 ( 
.A1(n_4214),
.A2(n_313),
.B(n_314),
.C(n_315),
.Y(n_4265)
);

NOR2xp33_ASAP7_75t_R g4266 ( 
.A(n_4206),
.B(n_314),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_4227),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4203),
.Y(n_4268)
);

NOR3xp33_ASAP7_75t_SL g4269 ( 
.A(n_4207),
.B(n_315),
.C(n_316),
.Y(n_4269)
);

OR2x2_ASAP7_75t_L g4270 ( 
.A(n_4225),
.B(n_317),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4209),
.Y(n_4271)
);

NOR2xp33_ASAP7_75t_L g4272 ( 
.A(n_4191),
.B(n_317),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_L g4273 ( 
.A(n_4223),
.B(n_318),
.Y(n_4273)
);

NOR2xp33_ASAP7_75t_L g4274 ( 
.A(n_4217),
.B(n_319),
.Y(n_4274)
);

AOI21xp5_ASAP7_75t_L g4275 ( 
.A1(n_4239),
.A2(n_4230),
.B(n_4220),
.Y(n_4275)
);

AOI22xp5_ASAP7_75t_SL g4276 ( 
.A1(n_4243),
.A2(n_4221),
.B1(n_4204),
.B2(n_4212),
.Y(n_4276)
);

OA22x2_ASAP7_75t_L g4277 ( 
.A1(n_4241),
.A2(n_4208),
.B1(n_4226),
.B2(n_4187),
.Y(n_4277)
);

NOR3xp33_ASAP7_75t_L g4278 ( 
.A(n_4242),
.B(n_4218),
.C(n_4196),
.Y(n_4278)
);

NOR2x1_ASAP7_75t_L g4279 ( 
.A(n_4244),
.B(n_4247),
.Y(n_4279)
);

OAI22xp5_ASAP7_75t_SL g4280 ( 
.A1(n_4234),
.A2(n_4231),
.B1(n_321),
.B2(n_322),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_4252),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4261),
.Y(n_4282)
);

AOI21xp5_ASAP7_75t_L g4283 ( 
.A1(n_4257),
.A2(n_4231),
.B(n_322),
.Y(n_4283)
);

AOI221x1_ASAP7_75t_SL g4284 ( 
.A1(n_4267),
.A2(n_320),
.B1(n_443),
.B2(n_445),
.C(n_448),
.Y(n_4284)
);

AO22x1_ASAP7_75t_L g4285 ( 
.A1(n_4236),
.A2(n_450),
.B1(n_451),
.B2(n_452),
.Y(n_4285)
);

OAI21xp5_ASAP7_75t_L g4286 ( 
.A1(n_4248),
.A2(n_453),
.B(n_455),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_4259),
.Y(n_4287)
);

NOR2x1p5_ASAP7_75t_L g4288 ( 
.A(n_4238),
.B(n_457),
.Y(n_4288)
);

NOR3xp33_ASAP7_75t_L g4289 ( 
.A(n_4263),
.B(n_458),
.C(n_460),
.Y(n_4289)
);

AOI22xp5_ASAP7_75t_L g4290 ( 
.A1(n_4272),
.A2(n_463),
.B1(n_464),
.B2(n_465),
.Y(n_4290)
);

AOI21xp5_ASAP7_75t_L g4291 ( 
.A1(n_4254),
.A2(n_1005),
.B(n_1044),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_L g4292 ( 
.A(n_4253),
.B(n_466),
.Y(n_4292)
);

INVx2_ASAP7_75t_L g4293 ( 
.A(n_4262),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4255),
.Y(n_4294)
);

XNOR2xp5_ASAP7_75t_L g4295 ( 
.A(n_4245),
.B(n_468),
.Y(n_4295)
);

NAND3xp33_ASAP7_75t_L g4296 ( 
.A(n_4246),
.B(n_1048),
.C(n_1007),
.Y(n_4296)
);

AND2x2_ASAP7_75t_L g4297 ( 
.A(n_4237),
.B(n_1007),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_SL g4298 ( 
.A(n_4264),
.B(n_1007),
.Y(n_4298)
);

INVxp67_ASAP7_75t_SL g4299 ( 
.A(n_4279),
.Y(n_4299)
);

INVxp67_ASAP7_75t_L g4300 ( 
.A(n_4280),
.Y(n_4300)
);

A2O1A1Ixp33_ASAP7_75t_L g4301 ( 
.A1(n_4284),
.A2(n_4265),
.B(n_4275),
.C(n_4283),
.Y(n_4301)
);

OR2x2_ASAP7_75t_L g4302 ( 
.A(n_4287),
.B(n_4249),
.Y(n_4302)
);

BUFx2_ASAP7_75t_L g4303 ( 
.A(n_4293),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4295),
.Y(n_4304)
);

AOI221xp5_ASAP7_75t_L g4305 ( 
.A1(n_4278),
.A2(n_4263),
.B1(n_4271),
.B2(n_4240),
.C(n_4289),
.Y(n_4305)
);

NAND2xp5_ASAP7_75t_L g4306 ( 
.A(n_4281),
.B(n_4251),
.Y(n_4306)
);

INVx1_ASAP7_75t_SL g4307 ( 
.A(n_4292),
.Y(n_4307)
);

INVxp67_ASAP7_75t_L g4308 ( 
.A(n_4282),
.Y(n_4308)
);

OR2x2_ASAP7_75t_L g4309 ( 
.A(n_4294),
.B(n_4260),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4277),
.Y(n_4310)
);

NAND3xp33_ASAP7_75t_L g4311 ( 
.A(n_4276),
.B(n_4269),
.C(n_4258),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4288),
.Y(n_4312)
);

NAND3xp33_ASAP7_75t_L g4313 ( 
.A(n_4296),
.B(n_4235),
.C(n_4241),
.Y(n_4313)
);

INVx2_ASAP7_75t_SL g4314 ( 
.A(n_4285),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_SL g4315 ( 
.A(n_4299),
.B(n_4266),
.Y(n_4315)
);

AOI31xp33_ASAP7_75t_L g4316 ( 
.A1(n_4300),
.A2(n_4268),
.A3(n_4273),
.B(n_4270),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_L g4317 ( 
.A(n_4310),
.B(n_4274),
.Y(n_4317)
);

NOR2x1_ASAP7_75t_L g4318 ( 
.A(n_4311),
.B(n_4256),
.Y(n_4318)
);

OA22x2_ASAP7_75t_L g4319 ( 
.A1(n_4314),
.A2(n_4286),
.B1(n_4290),
.B2(n_4250),
.Y(n_4319)
);

NAND3xp33_ASAP7_75t_L g4320 ( 
.A(n_4305),
.B(n_4235),
.C(n_4291),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_4303),
.Y(n_4321)
);

AOI22xp33_ASAP7_75t_L g4322 ( 
.A1(n_4313),
.A2(n_4297),
.B1(n_4298),
.B2(n_4290),
.Y(n_4322)
);

OAI22xp33_ASAP7_75t_L g4323 ( 
.A1(n_4306),
.A2(n_4308),
.B1(n_4302),
.B2(n_4312),
.Y(n_4323)
);

NOR2x1_ASAP7_75t_L g4324 ( 
.A(n_4301),
.B(n_1007),
.Y(n_4324)
);

AO22x2_ASAP7_75t_L g4325 ( 
.A1(n_4304),
.A2(n_1007),
.B1(n_1044),
.B2(n_1040),
.Y(n_4325)
);

OR2x2_ASAP7_75t_L g4326 ( 
.A(n_4321),
.B(n_4309),
.Y(n_4326)
);

AOI22xp5_ASAP7_75t_L g4327 ( 
.A1(n_4318),
.A2(n_4307),
.B1(n_1016),
.B2(n_1033),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_4323),
.B(n_1016),
.Y(n_4328)
);

NAND4xp25_ASAP7_75t_L g4329 ( 
.A(n_4317),
.B(n_1016),
.C(n_1044),
.D(n_1040),
.Y(n_4329)
);

AOI22xp33_ASAP7_75t_L g4330 ( 
.A1(n_4315),
.A2(n_1016),
.B1(n_1044),
.B2(n_1040),
.Y(n_4330)
);

AOI221xp5_ASAP7_75t_SL g4331 ( 
.A1(n_4316),
.A2(n_1016),
.B1(n_1044),
.B2(n_1040),
.C(n_1004),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4319),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_4326),
.Y(n_4333)
);

AOI22xp5_ASAP7_75t_L g4334 ( 
.A1(n_4332),
.A2(n_4320),
.B1(n_4322),
.B2(n_4324),
.Y(n_4334)
);

OR2x2_ASAP7_75t_L g4335 ( 
.A(n_4328),
.B(n_4325),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_L g4336 ( 
.A(n_4327),
.B(n_1016),
.Y(n_4336)
);

OAI22xp33_ASAP7_75t_L g4337 ( 
.A1(n_4329),
.A2(n_1005),
.B1(n_1044),
.B2(n_1040),
.Y(n_4337)
);

AOI22xp5_ASAP7_75t_L g4338 ( 
.A1(n_4333),
.A2(n_4331),
.B1(n_4330),
.B2(n_1033),
.Y(n_4338)
);

O2A1O1Ixp5_ASAP7_75t_SL g4339 ( 
.A1(n_4336),
.A2(n_4334),
.B(n_4337),
.C(n_4335),
.Y(n_4339)
);

NAND3x1_ASAP7_75t_L g4340 ( 
.A(n_4338),
.B(n_1005),
.C(n_1040),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_4339),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_4341),
.Y(n_4342)
);

NAND4xp25_ASAP7_75t_L g4343 ( 
.A(n_4342),
.B(n_4340),
.C(n_1005),
.D(n_1004),
.Y(n_4343)
);

BUFx2_ASAP7_75t_L g4344 ( 
.A(n_4343),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_L g4345 ( 
.A(n_4344),
.B(n_1033),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4345),
.Y(n_4346)
);

AOI21xp5_ASAP7_75t_L g4347 ( 
.A1(n_4346),
.A2(n_1033),
.B(n_1048),
.Y(n_4347)
);

INVx2_ASAP7_75t_L g4348 ( 
.A(n_4347),
.Y(n_4348)
);

AOI21xp33_ASAP7_75t_L g4349 ( 
.A1(n_4348),
.A2(n_1033),
.B(n_1048),
.Y(n_4349)
);

AOI22xp33_ASAP7_75t_SL g4350 ( 
.A1(n_4349),
.A2(n_1033),
.B1(n_1048),
.B2(n_955),
.Y(n_4350)
);

OAI221xp5_ASAP7_75t_R g4351 ( 
.A1(n_4349),
.A2(n_927),
.B1(n_930),
.B2(n_955),
.C(n_4334),
.Y(n_4351)
);

AOI221x1_ASAP7_75t_L g4352 ( 
.A1(n_4351),
.A2(n_927),
.B1(n_930),
.B2(n_955),
.C(n_4350),
.Y(n_4352)
);

AOI221xp5_ASAP7_75t_L g4353 ( 
.A1(n_4352),
.A2(n_927),
.B1(n_930),
.B2(n_955),
.C(n_4323),
.Y(n_4353)
);

AOI211xp5_ASAP7_75t_L g4354 ( 
.A1(n_4353),
.A2(n_955),
.B(n_927),
.C(n_930),
.Y(n_4354)
);


endmodule