module fake_netlist_6_734_n_954 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_954);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_954;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_671;
wire n_607;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_842;
wire n_758;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_184;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_880;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g184 ( 
.A(n_5),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_171),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_134),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_101),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_23),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_35),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_53),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_43),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_96),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_69),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_119),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_85),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_90),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_54),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_100),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_42),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_130),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_16),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_124),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_1),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_158),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_6),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_136),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_71),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_99),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_7),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_88),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_176),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_95),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_155),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_20),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_60),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_156),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_116),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_165),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_129),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_182),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_169),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_86),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_17),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_163),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_78),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_3),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_70),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_181),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_117),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_111),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_175),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_13),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_140),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_180),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_104),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_16),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_29),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_146),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_128),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_68),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_44),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_57),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_150),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_56),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_178),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_30),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_110),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_25),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_252),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_191),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_250),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_193),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_184),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_205),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_210),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_208),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_207),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_207),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_L g270 ( 
.A(n_219),
.B(n_0),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_203),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_220),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_229),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_238),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_254),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_240),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_219),
.B(n_0),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_212),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_232),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_189),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_189),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_219),
.B(n_1),
.Y(n_282)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_202),
.Y(n_283)
);

INVxp33_ASAP7_75t_SL g284 ( 
.A(n_187),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_218),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_240),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_246),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_246),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_202),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_247),
.Y(n_290)
);

INVxp33_ASAP7_75t_SL g291 ( 
.A(n_188),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_242),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_247),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_248),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_248),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_185),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_253),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_199),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_197),
.Y(n_299)
);

INVxp33_ASAP7_75t_SL g300 ( 
.A(n_194),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_199),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_198),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_186),
.Y(n_303)
);

INVxp33_ASAP7_75t_SL g304 ( 
.A(n_201),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_L g305 ( 
.A(n_231),
.B(n_2),
.Y(n_305)
);

INVxp33_ASAP7_75t_SL g306 ( 
.A(n_204),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_242),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_298),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_284),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_255),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_258),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_291),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_259),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_260),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_261),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_268),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_263),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_263),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_271),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_269),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_269),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_283),
.B(n_280),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_267),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_303),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_267),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_262),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_264),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_281),
.B(n_289),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_300),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_304),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_265),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_278),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_270),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_306),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_286),
.B(n_2),
.Y(n_340)
);

INVxp33_ASAP7_75t_L g341 ( 
.A(n_279),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_305),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_277),
.B(n_206),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_256),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_299),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_257),
.B(n_231),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_299),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_285),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_266),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_302),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_302),
.A2(n_224),
.B1(n_251),
.B2(n_249),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_282),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_266),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_274),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_276),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_272),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_273),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_274),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_297),
.B(n_253),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_275),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_276),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_275),
.B(n_190),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_296),
.B(n_192),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_287),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_292),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_290),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_317),
.Y(n_367)
);

BUFx10_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_330),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_356),
.B(n_287),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_309),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_309),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_352),
.B(n_343),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_356),
.B(n_288),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_343),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_343),
.B(n_209),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_307),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_360),
.B(n_288),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_312),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_338),
.B(n_195),
.Y(n_380)
);

INVx5_ASAP7_75t_L g381 ( 
.A(n_332),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_307),
.Y(n_382)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_332),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_312),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_343),
.B(n_211),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_332),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_332),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_332),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_327),
.B(n_253),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_308),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_332),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_360),
.B(n_294),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_338),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_346),
.A2(n_199),
.B1(n_196),
.B2(n_200),
.Y(n_395)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_341),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_358),
.B(n_294),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_365),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_330),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_313),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_327),
.B(n_215),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_357),
.B(n_295),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_333),
.B(n_221),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_333),
.B(n_225),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_365),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_330),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_313),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_362),
.A2(n_199),
.B1(n_230),
.B2(n_245),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_323),
.Y(n_409)
);

AND2x2_ASAP7_75t_SL g410 ( 
.A(n_358),
.B(n_3),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_315),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_314),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_314),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_331),
.A2(n_233),
.B1(n_216),
.B2(n_241),
.Y(n_414)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_329),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_355),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_315),
.Y(n_417)
);

AND2x2_ASAP7_75t_SL g418 ( 
.A(n_311),
.B(n_33),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_320),
.Y(n_419)
);

AND2x6_ASAP7_75t_L g420 ( 
.A(n_344),
.B(n_34),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_331),
.A2(n_228),
.B1(n_217),
.B2(n_239),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_363),
.B(n_295),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_357),
.B(n_213),
.Y(n_423)
);

INVx5_ASAP7_75t_L g424 ( 
.A(n_320),
.Y(n_424)
);

INVxp33_ASAP7_75t_L g425 ( 
.A(n_349),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_318),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_318),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_336),
.B(n_222),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_319),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_319),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_324),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_329),
.Y(n_432)
);

OAI22xp33_ASAP7_75t_SL g433 ( 
.A1(n_359),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_324),
.B(n_234),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_328),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_351),
.B(n_293),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_342),
.B(n_235),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_344),
.B(n_236),
.Y(n_438)
);

BUFx8_ASAP7_75t_SL g439 ( 
.A(n_337),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_325),
.B(n_237),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_415),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_373),
.B(n_344),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_438),
.B(n_344),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_405),
.B(n_353),
.Y(n_444)
);

AND2x6_ASAP7_75t_SL g445 ( 
.A(n_436),
.B(n_340),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_375),
.B(n_353),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_435),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_376),
.A2(n_354),
.B1(n_353),
.B2(n_334),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_390),
.B(n_353),
.Y(n_449)
);

A2O1A1Ixp33_ASAP7_75t_SL g450 ( 
.A1(n_406),
.A2(n_354),
.B(n_336),
.C(n_326),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_415),
.B(n_354),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_422),
.A2(n_354),
.B1(n_311),
.B2(n_347),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_415),
.B(n_316),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_335),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_411),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g456 ( 
.A1(n_410),
.A2(n_328),
.B1(n_325),
.B2(n_326),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_411),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g458 ( 
.A1(n_410),
.A2(n_342),
.B1(n_322),
.B2(n_321),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_401),
.B(n_339),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_390),
.B(n_345),
.Y(n_460)
);

OR2x6_ASAP7_75t_L g461 ( 
.A(n_377),
.B(n_366),
.Y(n_461)
);

NOR2xp67_ASAP7_75t_L g462 ( 
.A(n_378),
.B(n_350),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_417),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_377),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_384),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_398),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_417),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_401),
.B(n_321),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_369),
.B(n_322),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_369),
.B(n_361),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_394),
.B(n_364),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_387),
.B(n_36),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_387),
.B(n_366),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_382),
.B(n_340),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_418),
.A2(n_348),
.B1(n_5),
.B2(n_6),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_418),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_SL g477 ( 
.A(n_388),
.B(n_389),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_397),
.B(n_4),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_418),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_399),
.B(n_37),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_399),
.B(n_38),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_394),
.B(n_9),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_382),
.B(n_10),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_433),
.B(n_11),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_384),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_385),
.B(n_431),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_388),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_393),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_423),
.B(n_11),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_423),
.B(n_12),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_434),
.B(n_12),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_371),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_428),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_403),
.B(n_39),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_403),
.B(n_40),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_404),
.B(n_41),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_404),
.B(n_45),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_440),
.B(n_13),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_431),
.B(n_46),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_395),
.A2(n_94),
.B1(n_179),
.B2(n_177),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_428),
.A2(n_92),
.B1(n_174),
.B2(n_173),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_430),
.B(n_47),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_430),
.Y(n_503)
);

AND2x6_ASAP7_75t_SL g504 ( 
.A(n_380),
.B(n_437),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_412),
.B(n_48),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_412),
.B(n_432),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_437),
.B(n_14),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_371),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_372),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_412),
.B(n_49),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_408),
.A2(n_93),
.B1(n_172),
.B2(n_170),
.Y(n_511)
);

A2O1A1Ixp33_ASAP7_75t_L g512 ( 
.A1(n_380),
.A2(n_14),
.B(n_15),
.C(n_17),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_380),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_372),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_383),
.A2(n_97),
.B(n_167),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_432),
.B(n_50),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_426),
.B(n_51),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_428),
.B(n_414),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_379),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_421),
.B(n_15),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_379),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_426),
.B(n_52),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_461),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_447),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_455),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_492),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_473),
.Y(n_527)
);

A2O1A1Ixp33_ASAP7_75t_L g528 ( 
.A1(n_475),
.A2(n_429),
.B(n_427),
.C(n_425),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_508),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_441),
.B(n_416),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_457),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_488),
.B(n_370),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_449),
.A2(n_420),
.B1(n_374),
.B2(n_402),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_463),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_446),
.B(n_427),
.Y(n_535)
);

INVx6_ASAP7_75t_L g536 ( 
.A(n_504),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_467),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_461),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_441),
.B(n_429),
.Y(n_539)
);

CKINVDCx14_ASAP7_75t_R g540 ( 
.A(n_461),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_R g541 ( 
.A(n_474),
.B(n_367),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_503),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_466),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_469),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_473),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_442),
.A2(n_420),
.B1(n_386),
.B2(n_419),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_473),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_459),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_464),
.Y(n_549)
);

NOR3xp33_ASAP7_75t_SL g550 ( 
.A(n_460),
.B(n_409),
.C(n_367),
.Y(n_550)
);

AOI21xp33_ASAP7_75t_L g551 ( 
.A1(n_507),
.A2(n_396),
.B(n_409),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_493),
.B(n_420),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_443),
.B(n_419),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_509),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_483),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_445),
.Y(n_556)
);

NAND3xp33_ASAP7_75t_SL g557 ( 
.A(n_475),
.B(n_368),
.C(n_439),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_513),
.B(n_420),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_514),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_487),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_487),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_471),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_519),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_521),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_468),
.B(n_420),
.Y(n_565)
);

NOR3xp33_ASAP7_75t_SL g566 ( 
.A(n_448),
.B(n_439),
.C(n_368),
.Y(n_566)
);

OR2x2_ASAP7_75t_SL g567 ( 
.A(n_454),
.B(n_368),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_465),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_473),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_494),
.B(n_388),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_452),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_442),
.B(n_413),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_485),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_513),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_473),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_471),
.B(n_391),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_506),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_486),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_507),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_518),
.A2(n_420),
.B1(n_386),
.B2(n_413),
.Y(n_580)
);

CKINVDCx6p67_ASAP7_75t_R g581 ( 
.A(n_484),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_486),
.B(n_386),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_444),
.B(n_413),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_526),
.Y(n_584)
);

OAI21x1_ASAP7_75t_L g585 ( 
.A1(n_582),
.A2(n_480),
.B(n_472),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_524),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_544),
.B(n_456),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_574),
.B(n_453),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_560),
.Y(n_589)
);

AO31x2_ASAP7_75t_L g590 ( 
.A1(n_572),
.A2(n_490),
.A3(n_489),
.B(n_498),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_525),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_577),
.B(n_456),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_531),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_538),
.B(n_470),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_565),
.A2(n_451),
.B(n_497),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_572),
.A2(n_496),
.B(n_495),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_548),
.B(n_462),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_534),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_562),
.B(n_476),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_526),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_555),
.B(n_489),
.Y(n_601)
);

AOI221x1_ASAP7_75t_L g602 ( 
.A1(n_528),
.A2(n_490),
.B1(n_491),
.B2(n_498),
.C(n_511),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_570),
.A2(n_505),
.B(n_510),
.Y(n_603)
);

AO21x1_ASAP7_75t_L g604 ( 
.A1(n_570),
.A2(n_491),
.B(n_478),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_577),
.B(n_458),
.Y(n_605)
);

BUFx4f_ASAP7_75t_SL g606 ( 
.A(n_543),
.Y(n_606)
);

AOI31xp67_ASAP7_75t_L g607 ( 
.A1(n_580),
.A2(n_502),
.A3(n_481),
.B(n_499),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_578),
.B(n_458),
.Y(n_608)
);

OA22x2_ASAP7_75t_L g609 ( 
.A1(n_571),
.A2(n_579),
.B1(n_549),
.B2(n_533),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_543),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_538),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_532),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_523),
.B(n_558),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_578),
.B(n_476),
.Y(n_614)
);

NAND2x1p5_ASAP7_75t_L g615 ( 
.A(n_558),
.B(n_477),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_539),
.A2(n_450),
.B(n_481),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_535),
.A2(n_553),
.B(n_576),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_546),
.A2(n_450),
.B(n_520),
.Y(n_618)
);

BUFx12f_ASAP7_75t_L g619 ( 
.A(n_536),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_530),
.A2(n_522),
.B(n_517),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_L g621 ( 
.A1(n_528),
.A2(n_479),
.B(n_516),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_551),
.Y(n_622)
);

OAI21x1_ASAP7_75t_L g623 ( 
.A1(n_573),
.A2(n_515),
.B(n_501),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_567),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_530),
.A2(n_383),
.B(n_479),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_L g626 ( 
.A1(n_583),
.A2(n_500),
.B(n_482),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_579),
.A2(n_512),
.B1(n_400),
.B2(n_407),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_537),
.B(n_407),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_542),
.A2(n_392),
.B1(n_389),
.B2(n_388),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_536),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g631 ( 
.A1(n_529),
.A2(n_383),
.B(n_392),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_557),
.A2(n_413),
.B1(n_392),
.B2(n_389),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_554),
.Y(n_633)
);

OAI21x1_ASAP7_75t_L g634 ( 
.A1(n_631),
.A2(n_560),
.B(n_561),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_606),
.Y(n_635)
);

NOR2xp67_ASAP7_75t_L g636 ( 
.A(n_597),
.B(n_612),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_586),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_587),
.B(n_532),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_591),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_613),
.B(n_558),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_596),
.A2(n_569),
.B(n_552),
.Y(n_641)
);

O2A1O1Ixp33_ASAP7_75t_L g642 ( 
.A1(n_599),
.A2(n_564),
.B(n_559),
.C(n_563),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_593),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_622),
.B(n_581),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_601),
.B(n_536),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_619),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_584),
.Y(n_647)
);

NAND2x1p5_ASAP7_75t_L g648 ( 
.A(n_589),
.B(n_569),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_598),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_600),
.Y(n_650)
);

INVx6_ASAP7_75t_L g651 ( 
.A(n_613),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_595),
.A2(n_552),
.B(n_583),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_588),
.B(n_568),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_589),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_623),
.A2(n_575),
.B(n_527),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_630),
.B(n_556),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_595),
.A2(n_552),
.B(n_527),
.Y(n_657)
);

OAI21xp33_ASAP7_75t_SL g658 ( 
.A1(n_621),
.A2(n_545),
.B(n_547),
.Y(n_658)
);

O2A1O1Ixp5_ASAP7_75t_L g659 ( 
.A1(n_604),
.A2(n_566),
.B(n_550),
.C(n_545),
.Y(n_659)
);

AOI21xp33_ASAP7_75t_SL g660 ( 
.A1(n_609),
.A2(n_556),
.B(n_541),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_633),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_588),
.B(n_540),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_628),
.Y(n_663)
);

NAND2x1p5_ASAP7_75t_L g664 ( 
.A(n_594),
.B(n_527),
.Y(n_664)
);

OAI22xp33_ASAP7_75t_L g665 ( 
.A1(n_614),
.A2(n_541),
.B1(n_575),
.B2(n_527),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_611),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_615),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_628),
.Y(n_668)
);

OAI211xp5_ASAP7_75t_L g669 ( 
.A1(n_602),
.A2(n_540),
.B(n_547),
.C(n_575),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_615),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_608),
.Y(n_671)
);

OAI21x1_ASAP7_75t_L g672 ( 
.A1(n_603),
.A2(n_575),
.B(n_392),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_608),
.Y(n_673)
);

NOR2xp67_ASAP7_75t_SL g674 ( 
.A(n_610),
.B(n_388),
.Y(n_674)
);

OAI221xp5_ASAP7_75t_SL g675 ( 
.A1(n_614),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.C(n_21),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_594),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_587),
.B(n_413),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_617),
.B(n_389),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_627),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_609),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_627),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_592),
.A2(n_392),
.B1(n_389),
.B2(n_424),
.Y(n_682)
);

AND2x6_ASAP7_75t_L g683 ( 
.A(n_592),
.B(n_55),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_R g684 ( 
.A(n_646),
.B(n_605),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_636),
.A2(n_624),
.B1(n_626),
.B2(n_605),
.Y(n_685)
);

AOI222xp33_ASAP7_75t_L g686 ( 
.A1(n_645),
.A2(n_618),
.B1(n_590),
.B2(n_629),
.C1(n_22),
.C2(n_23),
.Y(n_686)
);

OR2x6_ASAP7_75t_L g687 ( 
.A(n_657),
.B(n_641),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_679),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_644),
.A2(n_638),
.B1(n_680),
.B2(n_676),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_637),
.Y(n_690)
);

AOI21x1_ASAP7_75t_L g691 ( 
.A1(n_652),
.A2(n_616),
.B(n_678),
.Y(n_691)
);

AOI222xp33_ASAP7_75t_L g692 ( 
.A1(n_638),
.A2(n_590),
.B1(n_629),
.B2(n_21),
.C1(n_22),
.C2(n_24),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_SL g693 ( 
.A1(n_680),
.A2(n_625),
.B1(n_617),
.B2(n_590),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_673),
.B(n_671),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_666),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_R g696 ( 
.A(n_662),
.B(n_625),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_640),
.B(n_632),
.Y(n_697)
);

AOI221xp5_ASAP7_75t_L g698 ( 
.A1(n_675),
.A2(n_660),
.B1(n_681),
.B2(n_643),
.C(n_639),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_665),
.A2(n_616),
.B1(n_620),
.B2(n_585),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_647),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_649),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_663),
.B(n_668),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_665),
.A2(n_620),
.B1(n_424),
.B2(n_381),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_661),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_R g705 ( 
.A(n_640),
.B(n_667),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_667),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_641),
.A2(n_607),
.B(n_381),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_657),
.A2(n_381),
.B(n_424),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_653),
.B(n_18),
.Y(n_709)
);

BUFx10_ASAP7_75t_L g710 ( 
.A(n_651),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_652),
.A2(n_424),
.B(n_381),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_651),
.B(n_19),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_651),
.B(n_58),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_650),
.B(n_24),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_654),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_664),
.B(n_670),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_683),
.A2(n_658),
.B1(n_677),
.B2(n_654),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_L g718 ( 
.A1(n_656),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_642),
.Y(n_719)
);

NAND3xp33_ASAP7_75t_SL g720 ( 
.A(n_659),
.B(n_26),
.C(n_27),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_669),
.A2(n_424),
.B1(n_381),
.B2(n_30),
.Y(n_721)
);

AOI221xp5_ASAP7_75t_L g722 ( 
.A1(n_675),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.C(n_32),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_642),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_635),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_669),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_664),
.B(n_59),
.Y(n_726)
);

OAI21x1_ASAP7_75t_L g727 ( 
.A1(n_672),
.A2(n_61),
.B(n_62),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_648),
.A2(n_678),
.B1(n_682),
.B2(n_659),
.Y(n_728)
);

AOI221xp5_ASAP7_75t_L g729 ( 
.A1(n_682),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.C(n_66),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_683),
.A2(n_67),
.B1(n_72),
.B2(n_73),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_683),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_731)
);

OR2x6_ASAP7_75t_L g732 ( 
.A(n_648),
.B(n_77),
.Y(n_732)
);

OAI22xp33_ASAP7_75t_L g733 ( 
.A1(n_683),
.A2(n_674),
.B1(n_655),
.B2(n_634),
.Y(n_733)
);

NAND3xp33_ASAP7_75t_SL g734 ( 
.A(n_683),
.B(n_79),
.C(n_80),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_679),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_647),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_680),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_638),
.B(n_84),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_647),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_637),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_689),
.B(n_87),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_695),
.Y(n_742)
);

AOI211xp5_ASAP7_75t_L g743 ( 
.A1(n_718),
.A2(n_722),
.B(n_725),
.C(n_720),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_SL g744 ( 
.A1(n_721),
.A2(n_89),
.B1(n_91),
.B2(n_98),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_690),
.B(n_102),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_724),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_701),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_686),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_702),
.B(n_107),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_711),
.A2(n_108),
.B(n_109),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_692),
.A2(n_720),
.B1(n_718),
.B2(n_734),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_710),
.Y(n_752)
);

OA21x2_ASAP7_75t_L g753 ( 
.A1(n_707),
.A2(n_112),
.B(n_113),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_706),
.B(n_115),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_704),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_740),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_688),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_712),
.B(n_118),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_684),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_688),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_735),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_710),
.Y(n_762)
);

OAI21x1_ASAP7_75t_L g763 ( 
.A1(n_707),
.A2(n_123),
.B(n_125),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_697),
.B(n_126),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_735),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_SL g766 ( 
.A1(n_732),
.A2(n_127),
.B(n_131),
.Y(n_766)
);

NAND3xp33_ASAP7_75t_L g767 ( 
.A(n_685),
.B(n_132),
.C(n_133),
.Y(n_767)
);

AO31x2_ASAP7_75t_L g768 ( 
.A1(n_728),
.A2(n_135),
.A3(n_137),
.B(n_138),
.Y(n_768)
);

A2O1A1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_729),
.A2(n_139),
.B(n_141),
.C(n_142),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_709),
.B(n_144),
.Y(n_770)
);

AOI221xp5_ASAP7_75t_L g771 ( 
.A1(n_698),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.C(n_151),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_687),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_734),
.A2(n_731),
.B(n_730),
.C(n_693),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_700),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_706),
.B(n_716),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_691),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_715),
.B(n_732),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_713),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_737),
.A2(n_152),
.B1(n_153),
.B2(n_157),
.Y(n_779)
);

BUFx12f_ASAP7_75t_L g780 ( 
.A(n_732),
.Y(n_780)
);

OAI21x1_ASAP7_75t_L g781 ( 
.A1(n_708),
.A2(n_160),
.B(n_161),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_738),
.B(n_694),
.Y(n_782)
);

AOI221xp5_ASAP7_75t_L g783 ( 
.A1(n_693),
.A2(n_162),
.B1(n_164),
.B2(n_166),
.C(n_183),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_736),
.B(n_739),
.Y(n_784)
);

BUFx10_ASAP7_75t_L g785 ( 
.A(n_719),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_715),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_726),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_747),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_757),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_776),
.B(n_687),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_747),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_776),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_757),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_763),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_785),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_785),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_761),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_755),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_760),
.Y(n_799)
);

INVxp67_ASAP7_75t_SL g800 ( 
.A(n_760),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_756),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_765),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_772),
.B(n_768),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_780),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_772),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_774),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_784),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_775),
.B(n_777),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_768),
.Y(n_809)
);

NAND2x1p5_ASAP7_75t_L g810 ( 
.A(n_753),
.B(n_723),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_768),
.B(n_699),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_768),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_775),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_782),
.B(n_717),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_787),
.B(n_714),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_753),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_777),
.B(n_727),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_753),
.B(n_703),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_782),
.B(n_733),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_773),
.B(n_786),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_741),
.B(n_745),
.Y(n_821)
);

NOR2x1_ASAP7_75t_L g822 ( 
.A(n_795),
.B(n_752),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_813),
.B(n_746),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_814),
.A2(n_748),
.B1(n_751),
.B2(n_771),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_803),
.B(n_786),
.Y(n_825)
);

AND2x4_ASAP7_75t_SL g826 ( 
.A(n_796),
.B(n_752),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_813),
.B(n_762),
.Y(n_827)
);

INVx1_ASAP7_75t_SL g828 ( 
.A(n_808),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_804),
.Y(n_829)
);

AO21x2_ASAP7_75t_L g830 ( 
.A1(n_809),
.A2(n_812),
.B(n_803),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_814),
.A2(n_748),
.B1(n_751),
.B2(n_743),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_820),
.A2(n_780),
.B1(n_773),
.B2(n_696),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_805),
.B(n_762),
.Y(n_833)
);

NOR4xp25_ASAP7_75t_SL g834 ( 
.A(n_809),
.B(n_705),
.C(n_812),
.D(n_783),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_821),
.A2(n_759),
.B1(n_744),
.B2(n_769),
.Y(n_835)
);

NAND4xp25_ASAP7_75t_L g836 ( 
.A(n_815),
.B(n_819),
.C(n_820),
.D(n_803),
.Y(n_836)
);

NOR3xp33_ASAP7_75t_L g837 ( 
.A(n_815),
.B(n_767),
.C(n_769),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_R g838 ( 
.A(n_804),
.B(n_742),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_788),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_798),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_839),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_827),
.B(n_819),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_828),
.B(n_808),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_825),
.B(n_805),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_825),
.B(n_807),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_833),
.B(n_807),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_823),
.B(n_808),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_839),
.B(n_805),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_840),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_836),
.B(n_806),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_830),
.B(n_790),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_830),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_832),
.B(n_806),
.Y(n_853)
);

CKINVDCx6p67_ASAP7_75t_R g854 ( 
.A(n_838),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_849),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_849),
.Y(n_856)
);

INVxp33_ASAP7_75t_L g857 ( 
.A(n_853),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_850),
.B(n_820),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_846),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_842),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_851),
.A2(n_831),
.B(n_824),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_848),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_844),
.B(n_822),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_845),
.B(n_811),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_851),
.B(n_799),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_861),
.B(n_844),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_855),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_863),
.B(n_860),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_863),
.B(n_843),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_859),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_856),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_857),
.B(n_847),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_858),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_857),
.B(n_854),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_864),
.B(n_848),
.Y(n_875)
);

NOR4xp25_ASAP7_75t_L g876 ( 
.A(n_874),
.B(n_824),
.C(n_835),
.D(n_852),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_869),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_870),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_866),
.B(n_854),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_873),
.B(n_862),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_878),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_877),
.Y(n_882)
);

OAI22xp33_ASAP7_75t_L g883 ( 
.A1(n_880),
.A2(n_873),
.B1(n_872),
.B2(n_868),
.Y(n_883)
);

INVx3_ASAP7_75t_SL g884 ( 
.A(n_881),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_882),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_883),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_881),
.B(n_876),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_884),
.B(n_879),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_887),
.B(n_868),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_885),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_887),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_886),
.B(n_871),
.Y(n_892)
);

NOR3x1_ASAP7_75t_L g893 ( 
.A(n_887),
.B(n_867),
.C(n_838),
.Y(n_893)
);

NOR4xp25_ASAP7_75t_L g894 ( 
.A(n_887),
.B(n_865),
.C(n_770),
.D(n_869),
.Y(n_894)
);

AOI21x1_ASAP7_75t_L g895 ( 
.A1(n_887),
.A2(n_875),
.B(n_865),
.Y(n_895)
);

AOI221xp5_ASAP7_75t_SL g896 ( 
.A1(n_891),
.A2(n_778),
.B1(n_811),
.B2(n_796),
.C(n_750),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_889),
.A2(n_829),
.B1(n_837),
.B2(n_804),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_888),
.Y(n_898)
);

AOI222xp33_ASAP7_75t_L g899 ( 
.A1(n_892),
.A2(n_811),
.B1(n_778),
.B2(n_829),
.C1(n_826),
.C2(n_818),
.Y(n_899)
);

OAI21xp33_ASAP7_75t_SL g900 ( 
.A1(n_894),
.A2(n_890),
.B(n_892),
.Y(n_900)
);

AOI211xp5_ASAP7_75t_L g901 ( 
.A1(n_893),
.A2(n_766),
.B(n_779),
.C(n_758),
.Y(n_901)
);

AOI21xp33_ASAP7_75t_L g902 ( 
.A1(n_895),
.A2(n_749),
.B(n_764),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_898),
.A2(n_899),
.B1(n_900),
.B2(n_897),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_901),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_896),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_902),
.A2(n_834),
.B1(n_826),
.B2(n_841),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_898),
.B(n_841),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_898),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_898),
.B(n_797),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_R g910 ( 
.A(n_898),
.B(n_795),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_898),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_908),
.B(n_808),
.Y(n_912)
);

NAND4xp25_ASAP7_75t_L g913 ( 
.A(n_903),
.B(n_821),
.C(n_754),
.D(n_795),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_911),
.Y(n_914)
);

XOR2xp5_ASAP7_75t_L g915 ( 
.A(n_904),
.B(n_754),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_907),
.B(n_802),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_907),
.B(n_905),
.Y(n_917)
);

NAND3xp33_ASAP7_75t_SL g918 ( 
.A(n_910),
.B(n_909),
.C(n_906),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_903),
.A2(n_796),
.B1(n_795),
.B2(n_802),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_911),
.Y(n_920)
);

NAND4xp25_ASAP7_75t_L g921 ( 
.A(n_913),
.B(n_808),
.C(n_817),
.D(n_790),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_914),
.Y(n_922)
);

OR4x1_ASAP7_75t_L g923 ( 
.A(n_920),
.B(n_797),
.C(n_789),
.D(n_781),
.Y(n_923)
);

NOR2x2_ASAP7_75t_L g924 ( 
.A(n_919),
.B(n_801),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_917),
.B(n_796),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_912),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_915),
.Y(n_927)
);

NOR2x1_ASAP7_75t_L g928 ( 
.A(n_918),
.B(n_796),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_916),
.B(n_796),
.Y(n_929)
);

OAI211xp5_ASAP7_75t_L g930 ( 
.A1(n_917),
.A2(n_796),
.B(n_816),
.C(n_799),
.Y(n_930)
);

AND3x2_ASAP7_75t_L g931 ( 
.A(n_922),
.B(n_800),
.C(n_817),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_926),
.Y(n_932)
);

NOR3xp33_ASAP7_75t_SL g933 ( 
.A(n_925),
.B(n_708),
.C(n_733),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_928),
.B(n_817),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_927),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_924),
.Y(n_936)
);

OAI221xp5_ASAP7_75t_L g937 ( 
.A1(n_921),
.A2(n_929),
.B1(n_930),
.B2(n_923),
.C(n_810),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_922),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_938),
.Y(n_939)
);

NOR2xp67_ASAP7_75t_L g940 ( 
.A(n_932),
.B(n_816),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_936),
.B(n_806),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_931),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_939),
.A2(n_935),
.B1(n_934),
.B2(n_937),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_941),
.A2(n_933),
.B(n_817),
.Y(n_944)
);

NOR4xp25_ASAP7_75t_SL g945 ( 
.A(n_943),
.B(n_942),
.C(n_940),
.D(n_933),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_944),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_945),
.B(n_798),
.Y(n_947)
);

XNOR2xp5_ASAP7_75t_L g948 ( 
.A(n_946),
.B(n_810),
.Y(n_948)
);

OA21x2_ASAP7_75t_L g949 ( 
.A1(n_946),
.A2(n_800),
.B(n_801),
.Y(n_949)
);

OAI321xp33_ASAP7_75t_L g950 ( 
.A1(n_947),
.A2(n_810),
.A3(n_794),
.B1(n_786),
.B2(n_789),
.C(n_801),
.Y(n_950)
);

AOI222xp33_ASAP7_75t_SL g951 ( 
.A1(n_948),
.A2(n_816),
.B1(n_798),
.B2(n_793),
.C1(n_792),
.C2(n_791),
.Y(n_951)
);

AOI222xp33_ASAP7_75t_L g952 ( 
.A1(n_950),
.A2(n_949),
.B1(n_794),
.B2(n_816),
.C1(n_786),
.C2(n_818),
.Y(n_952)
);

OAI221xp5_ASAP7_75t_R g953 ( 
.A1(n_952),
.A2(n_951),
.B1(n_949),
.B2(n_794),
.C(n_810),
.Y(n_953)
);

AOI211xp5_ASAP7_75t_L g954 ( 
.A1(n_953),
.A2(n_794),
.B(n_818),
.C(n_790),
.Y(n_954)
);


endmodule