module fake_jpeg_10921_n_432 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_432);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_432;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_5),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_10),
.B(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_57),
.A2(n_109),
.B1(n_42),
.B2(n_44),
.Y(n_165)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_9),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_59),
.B(n_89),
.Y(n_129)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_62),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_63),
.B(n_75),
.Y(n_121)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_64),
.Y(n_173)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_65),
.Y(n_164)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_21),
.B(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_86),
.Y(n_127)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_16),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_73),
.B(n_104),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_74),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_20),
.B(n_13),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_76),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_78),
.Y(n_179)
);

NAND2xp33_ASAP7_75t_SL g79 ( 
.A(n_35),
.B(n_0),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_48),
.Y(n_125)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_81),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_20),
.B(n_10),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_84),
.B(n_92),
.Y(n_144)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_100),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_36),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_91),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_24),
.B(n_11),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_24),
.B(n_11),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_93),
.B(n_99),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_94),
.Y(n_168)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g126 ( 
.A(n_97),
.Y(n_126)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_18),
.B(n_0),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_102),
.Y(n_169)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_105),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_108),
.Y(n_135)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_107),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_36),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_112),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_49),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_125),
.B(n_141),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_54),
.A2(n_23),
.B1(n_46),
.B2(n_26),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g215 ( 
.A1(n_131),
.A2(n_133),
.B1(n_153),
.B2(n_148),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_99),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_132),
.B(n_162),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_67),
.A2(n_23),
.B1(n_46),
.B2(n_26),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_75),
.B(n_18),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_134),
.B(n_136),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_84),
.B(n_52),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_52),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_138),
.B(n_151),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_56),
.A2(n_48),
.B1(n_49),
.B2(n_33),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_140),
.A2(n_175),
.B(n_183),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_59),
.A2(n_17),
.B(n_19),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_22),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_63),
.B(n_22),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_152),
.B(n_161),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_71),
.A2(n_19),
.B1(n_45),
.B2(n_44),
.Y(n_153)
);

AND2x6_ASAP7_75t_L g157 ( 
.A(n_91),
.B(n_1),
.Y(n_157)
);

AOI32xp33_ASAP7_75t_L g242 ( 
.A1(n_157),
.A2(n_132),
.A3(n_79),
.B1(n_73),
.B2(n_182),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_109),
.A2(n_49),
.B1(n_39),
.B2(n_28),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_160),
.A2(n_139),
.B(n_124),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_108),
.B(n_39),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_72),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_74),
.B(n_42),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_163),
.B(n_170),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_141),
.B1(n_129),
.B2(n_121),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_111),
.B(n_29),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_104),
.B(n_29),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_106),
.A2(n_33),
.B1(n_43),
.B2(n_45),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_112),
.B(n_43),
.Y(n_177)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_82),
.B(n_4),
.Y(n_178)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_83),
.A2(n_4),
.B1(n_6),
.B2(n_88),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_125),
.A2(n_94),
.B1(n_97),
.B2(n_165),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_185),
.A2(n_229),
.B1(n_242),
.B2(n_201),
.Y(n_282)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_157),
.A2(n_160),
.B1(n_150),
.B2(n_171),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_187),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_117),
.A2(n_166),
.B1(n_181),
.B2(n_143),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_188),
.Y(n_267)
);

BUFx4f_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_189),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_190),
.B(n_215),
.Y(n_243)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_126),
.Y(n_193)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_193),
.Y(n_266)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_195),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_175),
.A2(n_183),
.B1(n_171),
.B2(n_140),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_196),
.A2(n_228),
.B1(n_238),
.B2(n_236),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_122),
.A2(n_129),
.B1(n_139),
.B2(n_135),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_197),
.A2(n_225),
.B1(n_237),
.B2(n_203),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_182),
.A2(n_145),
.B1(n_176),
.B2(n_144),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_198),
.A2(n_220),
.B1(n_215),
.B2(n_230),
.Y(n_251)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_200),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_127),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_201),
.B(n_202),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_128),
.B(n_158),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_181),
.A2(n_142),
.B1(n_117),
.B2(n_155),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_203),
.A2(n_234),
.B(n_236),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_156),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_217),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_205),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_166),
.A2(n_143),
.B1(n_154),
.B2(n_155),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_206),
.A2(n_239),
.B1(n_205),
.B2(n_233),
.Y(n_277)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_207),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_114),
.B(n_158),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_208),
.B(n_213),
.Y(n_263)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_210),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_115),
.Y(n_211)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_212),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_114),
.B(n_120),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_216),
.Y(n_270)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_154),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_123),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_212),
.Y(n_245)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_222),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_145),
.A2(n_176),
.B1(n_115),
.B2(n_146),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_120),
.B(n_146),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_221),
.B(n_241),
.Y(n_268)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_137),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_113),
.B(n_116),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_223),
.B(n_193),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_130),
.A2(n_159),
.B1(n_147),
.B2(n_167),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_156),
.A2(n_118),
.B(n_113),
.C(n_126),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_230),
.B(n_190),
.C(n_223),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_147),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_227),
.B(n_232),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_130),
.A2(n_159),
.B1(n_137),
.B2(n_169),
.Y(n_229)
);

O2A1O1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_118),
.A2(n_116),
.B(n_148),
.C(n_119),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_231),
.Y(n_265)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

INVx11_ASAP7_75t_L g233 ( 
.A(n_119),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_180),
.A2(n_125),
.B(n_79),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_180),
.A2(n_125),
.B(n_79),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_180),
.A2(n_165),
.B1(n_122),
.B2(n_129),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_132),
.A2(n_25),
.B1(n_55),
.B2(n_58),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_122),
.B(n_63),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_244),
.B(n_261),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g286 ( 
.A(n_245),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_251),
.A2(n_253),
.B1(n_255),
.B2(n_259),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_252),
.B(n_246),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_198),
.B1(n_209),
.B2(n_237),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_209),
.C(n_197),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_257),
.B(n_258),
.C(n_271),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_185),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_187),
.A2(n_194),
.B1(n_234),
.B2(n_238),
.Y(n_259)
);

NAND3xp33_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_283),
.C(n_262),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_187),
.A2(n_220),
.B1(n_240),
.B2(n_221),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_269),
.A2(n_281),
.B1(n_285),
.B2(n_267),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_186),
.B(n_187),
.C(n_202),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_224),
.A2(n_208),
.B1(n_213),
.B2(n_225),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_243),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_282),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_224),
.A2(n_214),
.B1(n_192),
.B2(n_226),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_199),
.B(n_191),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_195),
.B(n_218),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_284),
.B(n_274),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_211),
.A2(n_210),
.B1(n_231),
.B2(n_189),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_276),
.A2(n_189),
.B(n_253),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_287),
.Y(n_334)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_254),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_291),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_276),
.A2(n_249),
.B(n_264),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_290),
.A2(n_306),
.B(n_273),
.Y(n_341)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_263),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_293),
.Y(n_320)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_263),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_262),
.B(n_268),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_296),
.Y(n_321)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_250),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_257),
.B(n_268),
.Y(n_297)
);

XNOR2x1_ASAP7_75t_L g337 ( 
.A(n_297),
.B(n_308),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_259),
.B(n_258),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_299),
.Y(n_323)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_265),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_300),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_271),
.B(n_264),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_304),
.Y(n_327)
);

INVx8_ASAP7_75t_L g304 ( 
.A(n_265),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_307),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_249),
.A2(n_281),
.B(n_255),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_247),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_243),
.B(n_261),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_309),
.B(n_285),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_248),
.B(n_270),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_313),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_243),
.B(n_269),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_312),
.A2(n_280),
.B(n_266),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_245),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_244),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_251),
.B(n_248),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_316),
.A2(n_265),
.B1(n_279),
.B2(n_272),
.Y(n_342)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_317),
.B(n_318),
.Y(n_340)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_278),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_287),
.A2(n_267),
.B(n_245),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_324),
.A2(n_333),
.B(n_338),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_315),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_325),
.B(n_328),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_288),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_256),
.Y(n_329)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_329),
.Y(n_356)
);

XOR2x1_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_331),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_295),
.B(n_266),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_308),
.A2(n_265),
.B1(n_280),
.B2(n_279),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_336),
.A2(n_342),
.B1(n_313),
.B2(n_296),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_314),
.A2(n_272),
.B(n_273),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_309),
.A2(n_293),
.B1(n_298),
.B2(n_308),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_339),
.A2(n_312),
.B1(n_301),
.B2(n_311),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_341),
.A2(n_301),
.B(n_286),
.Y(n_361)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_340),
.Y(n_344)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_344),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_337),
.B(n_297),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_350),
.Y(n_364)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_340),
.Y(n_347)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_347),
.Y(n_373)
);

NAND3xp33_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_332),
.C(n_323),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_355),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_335),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_349),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_337),
.B(n_294),
.C(n_290),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_294),
.C(n_311),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_351),
.B(n_352),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_307),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_353),
.A2(n_358),
.B1(n_325),
.B2(n_341),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_354),
.A2(n_339),
.B1(n_334),
.B2(n_302),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_301),
.C(n_306),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_319),
.B(n_303),
.Y(n_357)
);

NOR3xp33_ASAP7_75t_SL g378 ( 
.A(n_357),
.B(n_331),
.C(n_329),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_325),
.A2(n_316),
.B1(n_312),
.B2(n_302),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_327),
.B(n_339),
.C(n_323),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_359),
.B(n_363),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_361),
.A2(n_362),
.B(n_324),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_324),
.A2(n_302),
.B(n_318),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_329),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_343),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_365),
.Y(n_383)
);

XNOR2x2_ASAP7_75t_SL g366 ( 
.A(n_346),
.B(n_322),
.Y(n_366)
);

AOI21xp33_ASAP7_75t_L g384 ( 
.A1(n_366),
.A2(n_380),
.B(n_351),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_367),
.A2(n_368),
.B1(n_354),
.B2(n_343),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_358),
.A2(n_363),
.B1(n_356),
.B2(n_353),
.Y(n_368)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_369),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_371),
.A2(n_374),
.B(n_361),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_355),
.A2(n_341),
.B(n_322),
.Y(n_374)
);

OAI221xp5_ASAP7_75t_L g375 ( 
.A1(n_356),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.C(n_335),
.Y(n_375)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_375),
.Y(n_385)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_378),
.Y(n_391)
);

AOI322xp5_ASAP7_75t_L g380 ( 
.A1(n_362),
.A2(n_338),
.A3(n_320),
.B1(n_321),
.B2(n_330),
.C1(n_333),
.C2(n_342),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_381),
.B(n_384),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_350),
.C(n_359),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_386),
.B(n_393),
.C(n_377),
.Y(n_398)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_370),
.Y(n_387)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_387),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_388),
.A2(n_369),
.B1(n_365),
.B2(n_379),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_376),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_389),
.Y(n_399)
);

INVx6_ASAP7_75t_L g390 ( 
.A(n_378),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_390),
.A2(n_392),
.B1(n_375),
.B2(n_373),
.Y(n_401)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_370),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_364),
.B(n_360),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_383),
.A2(n_371),
.B(n_345),
.Y(n_394)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_394),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_383),
.A2(n_381),
.B(n_385),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_397),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_398),
.B(n_401),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_386),
.B(n_379),
.C(n_374),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_402),
.B(n_403),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_393),
.B(n_366),
.C(n_372),
.Y(n_403)
);

AO221x1_ASAP7_75t_L g404 ( 
.A1(n_396),
.A2(n_385),
.B1(n_373),
.B2(n_391),
.C(n_392),
.Y(n_404)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_404),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_402),
.B(n_368),
.C(n_382),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_407),
.B(n_408),
.Y(n_413)
);

OAI321xp33_ASAP7_75t_L g408 ( 
.A1(n_395),
.A2(n_390),
.A3(n_382),
.B1(n_387),
.B2(n_360),
.C(n_388),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_398),
.B(n_400),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_SL g415 ( 
.A(n_410),
.B(n_400),
.Y(n_415)
);

AO21x1_ASAP7_75t_L g414 ( 
.A1(n_406),
.A2(n_394),
.B(n_397),
.Y(n_414)
);

HAxp5_ASAP7_75t_L g421 ( 
.A(n_414),
.B(n_411),
.CON(n_421),
.SN(n_421)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_415),
.B(n_416),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_409),
.B(n_403),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_399),
.C(n_396),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_417),
.B(n_418),
.Y(n_422)
);

INVxp33_ASAP7_75t_L g418 ( 
.A(n_407),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_413),
.B(n_411),
.C(n_326),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_420),
.A2(n_421),
.B(n_418),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_289),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_423),
.B(n_338),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_424),
.A2(n_426),
.B(n_414),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_425),
.B(n_345),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_419),
.A2(n_422),
.B(n_421),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_427),
.B(n_428),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_429),
.A2(n_326),
.B(n_333),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_430),
.B(n_342),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_431),
.B(n_336),
.Y(n_432)
);


endmodule