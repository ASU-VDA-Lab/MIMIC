module fake_jpeg_15368_n_178 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_14),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_44),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_20),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_20),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_14),
.B1(n_16),
.B2(n_24),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_26),
.B1(n_16),
.B2(n_18),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_21),
.C(n_23),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_57),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_21),
.C(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_32),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_37),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_32),
.B1(n_36),
.B2(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_65),
.Y(n_78)
);

OA22x2_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_28),
.B1(n_18),
.B2(n_19),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_19),
.B1(n_28),
.B2(n_25),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_28),
.B1(n_22),
.B2(n_25),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_38),
.B1(n_37),
.B2(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_33),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_38),
.B1(n_48),
.B2(n_43),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_69),
.A2(n_74),
.B1(n_37),
.B2(n_40),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_75),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_68),
.B1(n_67),
.B2(n_51),
.Y(n_98)
);

AND2x4_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_56),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_79),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_40),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_15),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_51),
.B(n_49),
.Y(n_86)
);

A2O1A1O1Ixp25_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_53),
.B(n_33),
.C(n_17),
.D(n_63),
.Y(n_104)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_15),
.B1(n_23),
.B2(n_17),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_58),
.B1(n_66),
.B2(n_55),
.Y(n_101)
);

INVxp33_ASAP7_75t_SL g91 ( 
.A(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

AOI22x1_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_71),
.B1(n_62),
.B2(n_86),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_74),
.B1(n_71),
.B2(n_88),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_95),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_101),
.B1(n_0),
.B2(n_1),
.Y(n_122)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_105),
.B(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_89),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_108),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_109),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_112),
.A3(n_109),
.B1(n_115),
.B2(n_116),
.C1(n_106),
.C2(n_123),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_73),
.B1(n_88),
.B2(n_81),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_118),
.B1(n_122),
.B2(n_124),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_78),
.A3(n_70),
.B1(n_87),
.B2(n_40),
.Y(n_118)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_105),
.B(n_107),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_136),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_118),
.A2(n_104),
.B1(n_90),
.B2(n_101),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_137),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_103),
.B(n_94),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_116),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_131),
.C(n_130),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_144),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_146),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_120),
.C(n_111),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_111),
.Y(n_149)
);

NOR2xp67_ASAP7_75t_SL g154 ( 
.A(n_149),
.B(n_138),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_SL g150 ( 
.A(n_142),
.B(n_138),
.C(n_128),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_151),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_148),
.Y(n_151)
);

XNOR2x1_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_150),
.Y(n_162)
);

FAx1_ASAP7_75t_SL g155 ( 
.A(n_149),
.B(n_127),
.CI(n_126),
.CON(n_155),
.SN(n_155)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_142),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_156),
.B(n_9),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_145),
.A2(n_3),
.B(n_4),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_147),
.B(n_5),
.Y(n_158)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_141),
.C(n_143),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_160),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_162),
.A2(n_155),
.B1(n_157),
.B2(n_156),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_11),
.C(n_5),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_4),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_169),
.Y(n_172)
);

AOI31xp33_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_155),
.A3(n_5),
.B(n_8),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_8),
.B1(n_166),
.B2(n_168),
.Y(n_171)
);

OAI21x1_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_163),
.B(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_171),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_166),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_8),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

BUFx24_ASAP7_75t_SL g177 ( 
.A(n_176),
.Y(n_177)
);

XNOR2x2_ASAP7_75t_SL g178 ( 
.A(n_177),
.B(n_174),
.Y(n_178)
);


endmodule