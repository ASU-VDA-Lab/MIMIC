module fake_ariane_563_n_3010 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_345, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_15, n_23, n_87, n_279, n_207, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_221, n_321, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_155, n_127, n_3010);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_345;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_221;
input n_321;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_155;
input n_127;

output n_3010;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_2866;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_416;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_1837;
wire n_817;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_524;
wire n_2731;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_1298;
wire n_737;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_2976;
wire n_1835;
wire n_1457;
wire n_377;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_520;
wire n_870;
wire n_2547;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_1761;
wire n_829;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_557;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_2233;
wire n_2370;
wire n_2663;
wire n_495;
wire n_2914;
wire n_1988;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_2782;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_2950;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_432;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_2885;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_533;
wire n_2867;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_2739;
wire n_376;
wire n_512;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_491;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_461;
wire n_1416;
wire n_2909;
wire n_490;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2271;
wire n_2116;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2926;
wire n_482;
wire n_2620;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_2549;
wire n_2499;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_2791;
wire n_555;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_2970;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_514;
wire n_2748;
wire n_418;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2952;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_2922;
wire n_436;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_2628;
wire n_619;
wire n_967;
wire n_1083;
wire n_437;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2601;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_470;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_477;
wire n_650;
wire n_2388;
wire n_425;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_382;
wire n_489;
wire n_2294;
wire n_2274;
wire n_2895;
wire n_2903;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_397;
wire n_2467;
wire n_2768;
wire n_471;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_2924;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_404;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_2223;
wire n_836;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_370;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_466;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_552;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_379;
wire n_2834;
wire n_2483;
wire n_441;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_1592;
wire n_637;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_2811;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_405;
wire n_1611;
wire n_2122;
wire n_2975;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2998;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_481;
wire n_1609;
wire n_1053;
wire n_600;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_2937;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2783;
wire n_2599;
wire n_699;
wire n_590;
wire n_727;
wire n_1726;
wire n_2075;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_545;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_2853;
wire n_427;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_887;
wire n_729;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_390;
wire n_1156;
wire n_2741;
wire n_501;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2894;
wire n_2300;
wire n_2949;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_551;
wire n_417;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_2994;
wire n_534;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_451;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_2946;
wire n_1734;
wire n_1860;
wire n_403;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_2959;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_704;
wire n_2958;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2468;
wire n_2171;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_2992;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_1191;
wire n_618;
wire n_2492;
wire n_2939;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_1786;
wire n_2627;
wire n_480;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_642;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_602;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_2991;
wire n_1305;
wire n_2785;
wire n_730;
wire n_386;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_463;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_2928;
wire n_943;
wire n_1118;
wire n_678;
wire n_2905;
wire n_2884;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_649;
wire n_2412;
wire n_2720;
wire n_374;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_2907;
wire n_2386;
wire n_819;
wire n_1971;
wire n_2945;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_2936;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2986;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_2796;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_2947;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_368;
wire n_1958;
wire n_2747;
wire n_467;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2820;
wire n_2613;
wire n_497;
wire n_1165;
wire n_2934;
wire n_1641;
wire n_538;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_2647;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_413;
wire n_2401;
wire n_2935;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_685;
wire n_911;
wire n_361;
wire n_2658;
wire n_623;
wire n_2608;
wire n_2920;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_464;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_3008;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_2963;
wire n_519;
wire n_384;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_540;
wire n_2624;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_2938;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_2931;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2977;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_2828;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_2927;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_2180;
wire n_1942;
wire n_2951;
wire n_580;
wire n_1579;
wire n_494;
wire n_2809;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_2974;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_2858;
wire n_972;
wire n_2251;
wire n_2923;
wire n_2843;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2872;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_556;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_541;
wire n_499;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_2630;
wire n_591;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_1720;
wire n_663;
wire n_2409;
wire n_2966;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_385;
wire n_2395;
wire n_917;
wire n_2868;
wire n_2723;
wire n_1271;
wire n_372;
wire n_2440;
wire n_2556;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_399;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_363;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_2967;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_2948;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_2897;
wire n_1322;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_2973;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_369;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_3001;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2577;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2372;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2552;
wire n_2105;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2933;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_459;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_2846;
wire n_1781;
wire n_709;
wire n_2917;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_371;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_2513;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_2957;
wire n_865;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_450;
wire n_1923;
wire n_2955;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_2673;
wire n_1591;
wire n_664;
wire n_2585;
wire n_2995;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_537;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_389;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_719;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1252;
wire n_2239;
wire n_1129;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2940;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_2915;
wire n_431;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_2851;
wire n_2823;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_14),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_338),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_47),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_138),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_350),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_233),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_225),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_318),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_49),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_5),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_234),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_205),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_264),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_52),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_335),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_103),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_152),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_67),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_121),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_84),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_220),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_143),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_114),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_232),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_2),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_23),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_326),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_56),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_164),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_45),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_63),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_131),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_113),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_30),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_81),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_300),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_151),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_29),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_157),
.Y(n_397)
);

BUFx10_ASAP7_75t_L g398 ( 
.A(n_242),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_79),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_356),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_288),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_229),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_347),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_321),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_124),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_302),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_358),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_26),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_304),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_281),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_159),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_172),
.Y(n_412)
);

BUFx8_ASAP7_75t_SL g413 ( 
.A(n_227),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_128),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_27),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_333),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_278),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_263),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_219),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_87),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_103),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_125),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_116),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_248),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_355),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_322),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_206),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_23),
.Y(n_428)
);

INVxp33_ASAP7_75t_SL g429 ( 
.A(n_92),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_113),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_72),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_89),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_76),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_213),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_295),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_186),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_59),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_222),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_334),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_199),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_307),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_90),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_330),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_336),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_43),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_77),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_311),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_158),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_178),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_306),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_292),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_205),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_312),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_161),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_61),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_197),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_192),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_184),
.Y(n_458)
);

INVxp33_ASAP7_75t_SL g459 ( 
.A(n_308),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_186),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_324),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_115),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_31),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_174),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_101),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_293),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_178),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_343),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_320),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_121),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_6),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_291),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_109),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_212),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_353),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_237),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_245),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_38),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_253),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_172),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_211),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_349),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_174),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_108),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_150),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_239),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_298),
.Y(n_487)
);

BUFx10_ASAP7_75t_L g488 ( 
.A(n_228),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_95),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_93),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_86),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_331),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_244),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_45),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_327),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_284),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_269),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_200),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_348),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_257),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_11),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_3),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_195),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_143),
.Y(n_504)
);

INVxp33_ASAP7_75t_R g505 ( 
.A(n_251),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_351),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_272),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_132),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_139),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_12),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_133),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_117),
.Y(n_512)
);

CKINVDCx14_ASAP7_75t_R g513 ( 
.A(n_256),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_79),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_4),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_58),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_199),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_2),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_122),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_207),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_275),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_168),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_276),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_139),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_16),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_22),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_134),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_266),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_71),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_26),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_323),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_153),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_254),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_102),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_259),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_58),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_357),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_260),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_118),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_305),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_165),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_297),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_78),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_129),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_231),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_119),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_176),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_175),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_329),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_211),
.Y(n_550)
);

INVx1_ASAP7_75t_SL g551 ( 
.A(n_319),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_62),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_316),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_314),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_250),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_317),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_142),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_148),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_344),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_207),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_133),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_181),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_36),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_69),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_96),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_252),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_197),
.Y(n_567)
);

BUFx10_ASAP7_75t_L g568 ( 
.A(n_217),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_183),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_287),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_198),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_235),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_196),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_328),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_99),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_203),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_30),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_146),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_93),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_104),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_132),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_86),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_73),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_352),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_5),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_43),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_4),
.Y(n_587)
);

BUFx10_ASAP7_75t_L g588 ( 
.A(n_184),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_299),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_29),
.Y(n_590)
);

CKINVDCx14_ASAP7_75t_R g591 ( 
.A(n_52),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_125),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_273),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_70),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_57),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_44),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_145),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_17),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_309),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_296),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_34),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_44),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_53),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_32),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_7),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_301),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_310),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_313),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_354),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_325),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_95),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_20),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_111),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_315),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_339),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_37),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_337),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_303),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_200),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_78),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_188),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_160),
.Y(n_622)
);

BUFx10_ASAP7_75t_L g623 ( 
.A(n_27),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_277),
.Y(n_624)
);

BUFx8_ASAP7_75t_SL g625 ( 
.A(n_47),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_38),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_12),
.Y(n_627)
);

BUFx5_ASAP7_75t_L g628 ( 
.A(n_294),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_162),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_92),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_154),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_14),
.Y(n_632)
);

INVxp67_ASAP7_75t_SL g633 ( 
.A(n_215),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_345),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_7),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_161),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_346),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_332),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_163),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_255),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_36),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_53),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_194),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_70),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_127),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_49),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_63),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_138),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_124),
.Y(n_649)
);

INVxp67_ASAP7_75t_SL g650 ( 
.A(n_341),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_97),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_122),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_61),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_80),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_342),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_1),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_96),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_218),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_340),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_89),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_17),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_31),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_46),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_19),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_213),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_456),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_456),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_456),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_456),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_383),
.Y(n_670)
);

INVxp33_ASAP7_75t_SL g671 ( 
.A(n_421),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_591),
.Y(n_672)
);

INVxp33_ASAP7_75t_SL g673 ( 
.A(n_383),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_367),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_466),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_367),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_625),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_367),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_466),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_449),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_380),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_364),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_380),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_528),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_380),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_420),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_420),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_420),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_457),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_457),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_382),
.Y(n_691)
);

INVxp67_ASAP7_75t_SL g692 ( 
.A(n_457),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_382),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_385),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_612),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_385),
.Y(n_696)
);

INVxp33_ASAP7_75t_SL g697 ( 
.A(n_612),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_402),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_402),
.Y(n_699)
);

INVxp67_ASAP7_75t_L g700 ( 
.A(n_647),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_528),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_406),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_406),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_410),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_647),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_410),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_438),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_438),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_439),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_533),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_439),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_533),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_443),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_443),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_368),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_449),
.Y(n_716)
);

CKINVDCx16_ASAP7_75t_R g717 ( 
.A(n_370),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_444),
.Y(n_718)
);

INVxp67_ASAP7_75t_SL g719 ( 
.A(n_491),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_398),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_553),
.Y(n_721)
);

INVxp33_ASAP7_75t_SL g722 ( 
.A(n_359),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_370),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_491),
.Y(n_724)
);

INVxp67_ASAP7_75t_SL g725 ( 
.A(n_491),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_578),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_578),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_578),
.Y(n_728)
);

INVxp33_ASAP7_75t_SL g729 ( 
.A(n_361),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_368),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_636),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_636),
.Y(n_732)
);

CKINVDCx16_ASAP7_75t_R g733 ( 
.A(n_372),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_398),
.Y(n_734)
);

CKINVDCx16_ASAP7_75t_R g735 ( 
.A(n_372),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_398),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_636),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_398),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_651),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_488),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_387),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_379),
.Y(n_742)
);

CKINVDCx20_ASAP7_75t_R g743 ( 
.A(n_447),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_387),
.Y(n_744)
);

INVxp33_ASAP7_75t_SL g745 ( 
.A(n_362),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_488),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_651),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_651),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_572),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_660),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_488),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_660),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_488),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_396),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_660),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_661),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_661),
.Y(n_757)
);

INVxp67_ASAP7_75t_SL g758 ( 
.A(n_661),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_378),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_378),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_378),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_384),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_399),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_399),
.Y(n_764)
);

CKINVDCx16_ASAP7_75t_R g765 ( 
.A(n_384),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_413),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_399),
.Y(n_767)
);

INVxp67_ASAP7_75t_SL g768 ( 
.A(n_427),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_427),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_414),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_427),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_390),
.Y(n_772)
);

INVxp33_ASAP7_75t_L g773 ( 
.A(n_390),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_513),
.Y(n_774)
);

BUFx2_ASAP7_75t_SL g775 ( 
.A(n_401),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_432),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_432),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_432),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_470),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_374),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_470),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_375),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_470),
.Y(n_783)
);

INVxp67_ASAP7_75t_SL g784 ( 
.A(n_565),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_565),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_376),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_377),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_565),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_381),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_386),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_627),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_388),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_408),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_389),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_444),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_469),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_469),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_476),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_391),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_392),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_393),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_395),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_476),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_553),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_477),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_477),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_627),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_666),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_666),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_680),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_684),
.A2(n_455),
.B1(n_557),
.B2(n_509),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_667),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_721),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_680),
.Y(n_814)
);

INVxp33_ASAP7_75t_SL g815 ( 
.A(n_675),
.Y(n_815)
);

INVx4_ASAP7_75t_L g816 ( 
.A(n_721),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_721),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_667),
.Y(n_818)
);

INVx5_ASAP7_75t_L g819 ( 
.A(n_721),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_692),
.B(n_627),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_668),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_719),
.B(n_631),
.Y(n_822)
);

INVx5_ASAP7_75t_L g823 ( 
.A(n_721),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_668),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_804),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_725),
.B(n_631),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_758),
.B(n_631),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_762),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_716),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_728),
.B(n_412),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_804),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_684),
.A2(n_630),
.B1(n_429),
.B2(n_567),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_728),
.B(n_568),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_669),
.Y(n_834)
);

NAND2x1p5_ASAP7_75t_L g835 ( 
.A(n_691),
.B(n_409),
.Y(n_835)
);

INVx5_ASAP7_75t_L g836 ( 
.A(n_804),
.Y(n_836)
);

OA21x2_ASAP7_75t_L g837 ( 
.A1(n_716),
.A2(n_486),
.B(n_482),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_804),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_804),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_759),
.Y(n_840)
);

CKINVDCx6p67_ASAP7_75t_R g841 ( 
.A(n_717),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_701),
.A2(n_552),
.B1(n_604),
.B2(n_548),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_691),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_760),
.Y(n_844)
);

AOI22x1_ASAP7_75t_SL g845 ( 
.A1(n_677),
.A2(n_552),
.B1(n_405),
.B2(n_422),
.Y(n_845)
);

OAI21x1_ASAP7_75t_L g846 ( 
.A1(n_693),
.A2(n_805),
.B(n_803),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_710),
.B(n_412),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_776),
.B(n_568),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_693),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_694),
.B(n_449),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_694),
.Y(n_851)
);

INVx4_ASAP7_75t_L g852 ( 
.A(n_720),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_696),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_767),
.Y(n_854)
);

BUFx12f_ASAP7_75t_L g855 ( 
.A(n_766),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_768),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_761),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_762),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_701),
.A2(n_643),
.B1(n_423),
.B2(n_428),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_784),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_763),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_674),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_764),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_676),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_712),
.A2(n_586),
.B1(n_431),
.B2(n_433),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_769),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_712),
.A2(n_434),
.B1(n_440),
.B2(n_397),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_771),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_710),
.B(n_586),
.Y(n_869)
);

OA21x2_ASAP7_75t_L g870 ( 
.A1(n_696),
.A2(n_486),
.B(n_482),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_777),
.Y(n_871)
);

INVx5_ASAP7_75t_L g872 ( 
.A(n_776),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_733),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_735),
.Y(n_874)
);

NAND2xp33_ASAP7_75t_L g875 ( 
.A(n_698),
.B(n_449),
.Y(n_875)
);

INVx4_ASAP7_75t_L g876 ( 
.A(n_720),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_698),
.B(n_449),
.Y(n_877)
);

AND2x6_ASAP7_75t_L g878 ( 
.A(n_699),
.B(n_453),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_699),
.B(n_449),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_SL g880 ( 
.A1(n_754),
.A2(n_448),
.B1(n_452),
.B2(n_446),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_778),
.Y(n_881)
);

OA21x2_ASAP7_75t_L g882 ( 
.A1(n_702),
.A2(n_493),
.B(n_487),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_779),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_702),
.B(n_703),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_673),
.A2(n_458),
.B1(n_462),
.B2(n_454),
.Y(n_885)
);

BUFx12f_ASAP7_75t_L g886 ( 
.A(n_766),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_775),
.B(n_394),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_678),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_781),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_783),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_785),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_774),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_770),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_788),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_791),
.Y(n_895)
);

OA21x2_ASAP7_75t_L g896 ( 
.A1(n_703),
.A2(n_493),
.B(n_487),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_807),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_697),
.A2(n_465),
.B1(n_467),
.B2(n_464),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_765),
.Y(n_899)
);

INVx4_ASAP7_75t_L g900 ( 
.A(n_734),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_704),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_704),
.Y(n_902)
);

OAI22x1_ASAP7_75t_L g903 ( 
.A1(n_700),
.A2(n_705),
.B1(n_695),
.B2(n_670),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_706),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_706),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_707),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_707),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_773),
.B(n_568),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_708),
.Y(n_909)
);

AND2x6_ASAP7_75t_L g910 ( 
.A(n_708),
.B(n_453),
.Y(n_910)
);

BUFx8_ASAP7_75t_L g911 ( 
.A(n_709),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_734),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_774),
.B(n_640),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_709),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_711),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_711),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_713),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_775),
.B(n_496),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_681),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_671),
.A2(n_474),
.B1(n_483),
.B2(n_473),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_736),
.B(n_496),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_736),
.B(n_753),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_713),
.B(n_714),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_714),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_738),
.B(n_531),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_738),
.Y(n_926)
);

AO22x1_ASAP7_75t_L g927 ( 
.A1(n_718),
.A2(n_633),
.B1(n_796),
.B2(n_795),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_740),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_715),
.B(n_568),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_740),
.B(n_409),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_675),
.A2(n_485),
.B1(n_490),
.B2(n_484),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_718),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_855),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_843),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_843),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_884),
.B(n_795),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_855),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_873),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_893),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_886),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_886),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_849),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_893),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_874),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_892),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_892),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_841),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_810),
.Y(n_948)
);

BUFx2_ASAP7_75t_SL g949 ( 
.A(n_912),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_810),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_905),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_841),
.Y(n_952)
);

CKINVDCx16_ASAP7_75t_R g953 ( 
.A(n_899),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_911),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_828),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_911),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_849),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_851),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_911),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_814),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_SL g961 ( 
.A(n_815),
.B(n_679),
.Y(n_961)
);

CKINVDCx20_ASAP7_75t_R g962 ( 
.A(n_828),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_858),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_814),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_815),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_R g966 ( 
.A(n_912),
.B(n_679),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_858),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_851),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_909),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_909),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_922),
.B(n_672),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_916),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_829),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_926),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_930),
.A2(n_751),
.B1(n_753),
.B2(n_746),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_R g976 ( 
.A(n_926),
.B(n_682),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_916),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_880),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_811),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_852),
.B(n_876),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_852),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_852),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_932),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_876),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_876),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_829),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_932),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_908),
.Y(n_988)
);

NOR2x1p5_ASAP7_75t_L g989 ( 
.A(n_900),
.B(n_746),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_832),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_900),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_809),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_900),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_928),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_872),
.B(n_751),
.Y(n_995)
);

NOR2xp67_ASAP7_75t_L g996 ( 
.A(n_928),
.B(n_872),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_809),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_928),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_931),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_862),
.Y(n_1000)
);

OA21x2_ASAP7_75t_L g1001 ( 
.A1(n_846),
.A2(n_797),
.B(n_796),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_905),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_812),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_812),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_862),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_846),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_R g1007 ( 
.A(n_853),
.B(n_742),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_816),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_919),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_818),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_919),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_867),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_840),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_R g1014 ( 
.A(n_853),
.B(n_743),
.Y(n_1014)
);

CKINVDCx16_ASAP7_75t_R g1015 ( 
.A(n_908),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_818),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_840),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_905),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_845),
.Y(n_1019)
);

CKINVDCx16_ASAP7_75t_R g1020 ( 
.A(n_833),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_845),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_920),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_885),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_898),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_913),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_859),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_905),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_816),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_833),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_865),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_835),
.B(n_722),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_927),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_848),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_R g1034 ( 
.A(n_848),
.B(n_780),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_905),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_927),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_872),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_929),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_872),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_921),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_821),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_906),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_R g1043 ( 
.A(n_853),
.B(n_749),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_925),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_887),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_872),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_929),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_854),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_856),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_884),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_860),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_918),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_842),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_903),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_884),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_906),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_903),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_821),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_820),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_820),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_906),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_R g1062 ( 
.A(n_902),
.B(n_672),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_820),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_816),
.Y(n_1064)
);

NAND2xp33_ASAP7_75t_R g1065 ( 
.A(n_830),
.B(n_780),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_864),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_888),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_822),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_824),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_824),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_901),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_834),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_R g1073 ( 
.A(n_902),
.B(n_782),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_822),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_923),
.B(n_797),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_R g1076 ( 
.A(n_902),
.B(n_782),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_840),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_822),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_826),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_906),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_826),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_826),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_906),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_R g1084 ( 
.A(n_808),
.B(n_786),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_914),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_923),
.B(n_798),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_840),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_901),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_840),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_914),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_904),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_914),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_857),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_914),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_R g1095 ( 
.A(n_808),
.B(n_786),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_914),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_825),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_904),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_917),
.Y(n_1099)
);

CKINVDCx16_ASAP7_75t_R g1100 ( 
.A(n_830),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_SL g1101 ( 
.A(n_835),
.B(n_505),
.Y(n_1101)
);

OR2x2_ASAP7_75t_L g1102 ( 
.A(n_830),
.B(n_723),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_827),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_951),
.Y(n_1104)
);

OR2x2_ASAP7_75t_L g1105 ( 
.A(n_953),
.B(n_835),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_992),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_948),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_1040),
.B(n_729),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_938),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_1013),
.Y(n_1110)
);

INVx4_ASAP7_75t_SL g1111 ( 
.A(n_1013),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1052),
.B(n_923),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_944),
.Y(n_1113)
);

AND2x6_ASAP7_75t_L g1114 ( 
.A(n_936),
.B(n_877),
.Y(n_1114)
);

AND2x6_ASAP7_75t_L g1115 ( 
.A(n_936),
.B(n_877),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_951),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_948),
.Y(n_1117)
);

INVx4_ASAP7_75t_L g1118 ( 
.A(n_1013),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_950),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1044),
.B(n_1045),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1075),
.B(n_827),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1075),
.B(n_1086),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_1086),
.B(n_827),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_997),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_1013),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1050),
.B(n_808),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_955),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1003),
.Y(n_1128)
);

INVx4_ASAP7_75t_SL g1129 ( 
.A(n_1013),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_1080),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_1025),
.B(n_745),
.Y(n_1131)
);

INVx5_ASAP7_75t_L g1132 ( 
.A(n_1006),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_950),
.Y(n_1133)
);

NAND2xp33_ASAP7_75t_L g1134 ( 
.A(n_981),
.B(n_917),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1025),
.A2(n_459),
.B1(n_869),
.B2(n_847),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1055),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_960),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_960),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_974),
.B(n_787),
.Y(n_1139)
);

AO21x2_ASAP7_75t_L g1140 ( 
.A1(n_1002),
.A2(n_542),
.B(n_531),
.Y(n_1140)
);

INVx5_ASAP7_75t_L g1141 ( 
.A(n_1006),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1017),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1004),
.Y(n_1143)
);

AND2x6_ASAP7_75t_L g1144 ( 
.A(n_1006),
.B(n_877),
.Y(n_1144)
);

INVx4_ASAP7_75t_L g1145 ( 
.A(n_1017),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_1017),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_1017),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1015),
.B(n_787),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1074),
.B(n_847),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1010),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1074),
.B(n_847),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_989),
.B(n_869),
.Y(n_1152)
);

AO22x2_ASAP7_75t_L g1153 ( 
.A1(n_1101),
.A2(n_869),
.B1(n_505),
.B2(n_803),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_1017),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_982),
.B(n_917),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_1077),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_964),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_964),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_949),
.B(n_792),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_973),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_973),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1020),
.B(n_792),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_939),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1016),
.Y(n_1164)
);

AND2x6_ASAP7_75t_L g1165 ( 
.A(n_1002),
.B(n_879),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_986),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1041),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1078),
.B(n_907),
.Y(n_1168)
);

NAND3x1_ASAP7_75t_L g1169 ( 
.A(n_975),
.B(n_411),
.C(n_408),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1058),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1069),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_1077),
.Y(n_1172)
);

INVx5_ASAP7_75t_L g1173 ( 
.A(n_1077),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_986),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1094),
.B(n_879),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1071),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1070),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1077),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_984),
.B(n_985),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_943),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1077),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1088),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_934),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1091),
.Y(n_1184)
);

AND2x6_ASAP7_75t_L g1185 ( 
.A(n_1018),
.B(n_1027),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1098),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1099),
.B(n_879),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_1000),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1018),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_935),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_SL g1191 ( 
.A(n_933),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_1087),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_1005),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1027),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_1087),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_1009),
.Y(n_1196)
);

BUFx10_ASAP7_75t_L g1197 ( 
.A(n_965),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_942),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1078),
.B(n_907),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_962),
.Y(n_1200)
);

INVx5_ASAP7_75t_L g1201 ( 
.A(n_1087),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1087),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_957),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1007),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_1014),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1079),
.B(n_915),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1026),
.B(n_800),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_958),
.Y(n_1208)
);

INVx5_ASAP7_75t_L g1209 ( 
.A(n_1087),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_968),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1011),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1035),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_991),
.B(n_800),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1089),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_969),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_970),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1089),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_972),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_993),
.B(n_801),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1089),
.Y(n_1220)
);

NOR3xp33_ASAP7_75t_L g1221 ( 
.A(n_967),
.B(n_946),
.C(n_945),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_947),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1035),
.Y(n_1223)
);

AND3x1_ASAP7_75t_L g1224 ( 
.A(n_961),
.B(n_415),
.C(n_411),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_977),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_983),
.Y(n_1226)
);

INVxp67_ASAP7_75t_SL g1227 ( 
.A(n_1008),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_945),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_947),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_987),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1042),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1089),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_994),
.B(n_917),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1042),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1089),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1001),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_963),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1001),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1001),
.Y(n_1239)
);

INVx4_ASAP7_75t_L g1240 ( 
.A(n_1093),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1056),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1056),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_998),
.B(n_917),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1032),
.A2(n_837),
.B1(n_910),
.B2(n_878),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1043),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1061),
.Y(n_1246)
);

AND2x6_ASAP7_75t_L g1247 ( 
.A(n_1061),
.B(n_453),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1083),
.Y(n_1248)
);

NAND2xp33_ASAP7_75t_L g1249 ( 
.A(n_966),
.B(n_878),
.Y(n_1249)
);

INVx4_ASAP7_75t_L g1250 ( 
.A(n_1093),
.Y(n_1250)
);

AND2x6_ASAP7_75t_L g1251 ( 
.A(n_1083),
.B(n_1085),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1026),
.B(n_801),
.Y(n_1252)
);

INVx2_ASAP7_75t_SL g1253 ( 
.A(n_1079),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_1081),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1073),
.B(n_915),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1085),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_1093),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1081),
.B(n_924),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1090),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_SL g1260 ( 
.A(n_933),
.B(n_789),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1093),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1082),
.B(n_924),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_946),
.Y(n_1263)
);

INVx4_ASAP7_75t_L g1264 ( 
.A(n_1093),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1031),
.B(n_683),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1090),
.Y(n_1266)
);

INVx4_ASAP7_75t_L g1267 ( 
.A(n_1008),
.Y(n_1267)
);

INVx5_ASAP7_75t_L g1268 ( 
.A(n_1008),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1092),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1092),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_976),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1096),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1096),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_952),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1076),
.B(n_1084),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1082),
.B(n_844),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1103),
.B(n_798),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1028),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1028),
.Y(n_1279)
);

INVx4_ASAP7_75t_L g1280 ( 
.A(n_1028),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1095),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1103),
.B(n_805),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1100),
.B(n_1102),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1059),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1064),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1062),
.B(n_988),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1047),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1060),
.B(n_806),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1063),
.B(n_844),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1064),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1068),
.B(n_971),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1032),
.A2(n_1036),
.B1(n_1053),
.B2(n_1012),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1036),
.B(n_790),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_999),
.A2(n_837),
.B1(n_910),
.B2(n_878),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1064),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1097),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1097),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1030),
.B(n_794),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1030),
.B(n_799),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1130),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1106),
.Y(n_1301)
);

NOR3xp33_ASAP7_75t_L g1302 ( 
.A(n_1131),
.B(n_1024),
.C(n_1023),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1168),
.B(n_1048),
.Y(n_1303)
);

OR2x2_ASAP7_75t_SL g1304 ( 
.A(n_1120),
.B(n_978),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1107),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1107),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1117),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_SL g1308 ( 
.A(n_1222),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1291),
.B(n_1023),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1290),
.B(n_996),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1109),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1168),
.B(n_1049),
.Y(n_1312)
);

BUFx8_ASAP7_75t_L g1313 ( 
.A(n_1191),
.Y(n_1313)
);

CKINVDCx11_ASAP7_75t_R g1314 ( 
.A(n_1180),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1298),
.B(n_1029),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1199),
.B(n_1051),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1106),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1109),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1199),
.B(n_1033),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1299),
.B(n_1024),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1159),
.A2(n_1038),
.B(n_995),
.C(n_1097),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1112),
.B(n_1022),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1207),
.A2(n_1034),
.B1(n_1065),
.B2(n_990),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1124),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1124),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1128),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1117),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1128),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1290),
.B(n_1267),
.Y(n_1329)
);

NOR3xp33_ASAP7_75t_L g1330 ( 
.A(n_1108),
.B(n_940),
.C(n_937),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1143),
.A2(n_980),
.B(n_806),
.C(n_1037),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1206),
.B(n_1037),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1143),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1150),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1253),
.B(n_1254),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1122),
.B(n_954),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_SL g1337 ( 
.A1(n_1200),
.A2(n_979),
.B1(n_1021),
.B2(n_1019),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1206),
.B(n_1039),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1150),
.A2(n_1039),
.B1(n_1046),
.B2(n_1072),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1170),
.A2(n_501),
.B1(n_502),
.B2(n_498),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1119),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1277),
.B(n_954),
.Y(n_1342)
);

INVxp67_ASAP7_75t_L g1343 ( 
.A(n_1113),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1282),
.B(n_956),
.Y(n_1344)
);

NOR2xp67_ASAP7_75t_L g1345 ( 
.A(n_1139),
.B(n_937),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1126),
.B(n_1123),
.Y(n_1346)
);

OAI22xp33_ASAP7_75t_SL g1347 ( 
.A1(n_1252),
.A2(n_1057),
.B1(n_1054),
.B2(n_956),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1170),
.A2(n_508),
.B1(n_510),
.B2(n_504),
.Y(n_1348)
);

OR2x6_ASAP7_75t_L g1349 ( 
.A(n_1130),
.B(n_952),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1126),
.B(n_959),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1253),
.A2(n_1066),
.B1(n_1067),
.B2(n_959),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1254),
.B(n_802),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1149),
.B(n_940),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1123),
.B(n_941),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1123),
.B(n_868),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1149),
.B(n_941),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1119),
.Y(n_1357)
);

NOR3xp33_ASAP7_75t_L g1358 ( 
.A(n_1162),
.B(n_419),
.C(n_415),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1276),
.B(n_868),
.Y(n_1359)
);

OAI221xp5_ASAP7_75t_L g1360 ( 
.A1(n_1224),
.A2(n_744),
.B1(n_772),
.B2(n_741),
.C(n_730),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_1113),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1198),
.A2(n_515),
.B1(n_516),
.B2(n_511),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1281),
.B(n_857),
.Y(n_1363)
);

NAND2xp33_ASAP7_75t_L g1364 ( 
.A(n_1290),
.B(n_878),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1151),
.B(n_793),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1198),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1114),
.A2(n_650),
.B1(n_507),
.B2(n_551),
.Y(n_1367)
);

CKINVDCx11_ASAP7_75t_R g1368 ( 
.A(n_1180),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1203),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1151),
.B(n_517),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1258),
.B(n_1262),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1290),
.B(n_825),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1276),
.B(n_871),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1203),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1121),
.B(n_519),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1208),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1288),
.B(n_871),
.Y(n_1377)
);

AOI221xp5_ASAP7_75t_L g1378 ( 
.A1(n_1148),
.A2(n_436),
.B1(n_437),
.B2(n_430),
.C(n_419),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1208),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1275),
.A2(n_436),
.B(n_437),
.C(n_430),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1215),
.Y(n_1381)
);

NAND3xp33_ASAP7_75t_L g1382 ( 
.A(n_1228),
.B(n_525),
.C(n_522),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1293),
.B(n_527),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1289),
.B(n_881),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1188),
.B(n_857),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1215),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1216),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1188),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1289),
.B(n_1114),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1271),
.B(n_685),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1114),
.B(n_881),
.Y(n_1391)
);

O2A1O1Ixp5_ASAP7_75t_L g1392 ( 
.A1(n_1155),
.A2(n_831),
.B(n_825),
.C(n_883),
.Y(n_1392)
);

AND2x6_ASAP7_75t_L g1393 ( 
.A(n_1290),
.B(n_495),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1135),
.B(n_529),
.Y(n_1394)
);

BUFx8_ASAP7_75t_L g1395 ( 
.A(n_1191),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1193),
.B(n_857),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1114),
.B(n_883),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1133),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1114),
.B(n_890),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1133),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1137),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1114),
.B(n_890),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1153),
.A2(n_878),
.B1(n_910),
.B2(n_882),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1115),
.B(n_891),
.Y(n_1404)
);

AOI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1115),
.A2(n_507),
.B1(n_551),
.B2(n_441),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1153),
.A2(n_878),
.B1(n_910),
.B2(n_882),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1284),
.B(n_534),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1193),
.B(n_857),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1284),
.B(n_536),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1283),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1115),
.B(n_891),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1196),
.B(n_861),
.Y(n_1412)
);

BUFx8_ASAP7_75t_L g1413 ( 
.A(n_1191),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1115),
.B(n_894),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1137),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1196),
.B(n_861),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1115),
.B(n_894),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1211),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1115),
.B(n_895),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1216),
.Y(n_1420)
);

OR2x6_ASAP7_75t_L g1421 ( 
.A(n_1222),
.B(n_895),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1236),
.A2(n_882),
.B(n_870),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1175),
.B(n_539),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1267),
.B(n_1280),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1271),
.B(n_686),
.Y(n_1425)
);

NOR2x1_ASAP7_75t_L g1426 ( 
.A(n_1211),
.B(n_897),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1218),
.B(n_897),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1218),
.B(n_861),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1138),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1153),
.A2(n_910),
.B1(n_882),
.B2(n_896),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_SL g1431 ( 
.A(n_1228),
.B(n_1019),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1225),
.Y(n_1432)
);

NOR2xp67_ASAP7_75t_L g1433 ( 
.A(n_1263),
.B(n_1021),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1153),
.A2(n_910),
.B1(n_896),
.B2(n_870),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1225),
.A2(n_544),
.B1(n_546),
.B2(n_541),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1138),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1226),
.B(n_861),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1226),
.B(n_861),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1152),
.B(n_863),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1175),
.B(n_550),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1164),
.B(n_863),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1167),
.Y(n_1442)
);

AND2x4_ASAP7_75t_SL g1443 ( 
.A(n_1197),
.B(n_588),
.Y(n_1443)
);

INVxp67_ASAP7_75t_L g1444 ( 
.A(n_1127),
.Y(n_1444)
);

NOR2xp67_ASAP7_75t_L g1445 ( 
.A(n_1263),
.B(n_687),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1171),
.A2(n_896),
.B1(n_870),
.B2(n_863),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1157),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1177),
.B(n_863),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1283),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1127),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1183),
.B(n_863),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1320),
.B(n_1287),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1424),
.A2(n_1141),
.B(n_1132),
.Y(n_1453)
);

NAND2xp33_ASAP7_75t_L g1454 ( 
.A(n_1321),
.B(n_1144),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1388),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1311),
.Y(n_1456)
);

BUFx8_ASAP7_75t_L g1457 ( 
.A(n_1308),
.Y(n_1457)
);

INVx5_ASAP7_75t_L g1458 ( 
.A(n_1393),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1371),
.B(n_1175),
.Y(n_1459)
);

NAND3xp33_ASAP7_75t_L g1460 ( 
.A(n_1320),
.B(n_1221),
.C(n_1260),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1322),
.B(n_1200),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1305),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1311),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1424),
.A2(n_1141),
.B(n_1132),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1371),
.A2(n_1141),
.B(n_1132),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1310),
.A2(n_1141),
.B(n_1132),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1310),
.A2(n_1141),
.B(n_1132),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1422),
.A2(n_1239),
.B(n_1238),
.Y(n_1468)
);

O2A1O1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1358),
.A2(n_1213),
.B(n_1219),
.C(n_1286),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1446),
.A2(n_1210),
.B(n_1190),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1301),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1306),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1329),
.A2(n_1134),
.B(n_1233),
.Y(n_1473)
);

OAI321xp33_ASAP7_75t_L g1474 ( 
.A1(n_1378),
.A2(n_460),
.A3(n_442),
.B1(n_478),
.B2(n_471),
.C(n_445),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1388),
.Y(n_1475)
);

O2A1O1Ixp5_ASAP7_75t_L g1476 ( 
.A1(n_1309),
.A2(n_1243),
.B(n_1179),
.C(n_1255),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1322),
.B(n_1105),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1329),
.A2(n_1134),
.B(n_1227),
.Y(n_1478)
);

OAI21xp33_ASAP7_75t_L g1479 ( 
.A1(n_1365),
.A2(n_1136),
.B(n_1230),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1331),
.A2(n_1249),
.B(n_1267),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1315),
.B(n_1105),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1343),
.B(n_1237),
.Y(n_1482)
);

INVx11_ASAP7_75t_L g1483 ( 
.A(n_1313),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1307),
.Y(n_1484)
);

INVx5_ASAP7_75t_L g1485 ( 
.A(n_1393),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1317),
.A2(n_1169),
.B1(n_1294),
.B2(n_1280),
.Y(n_1486)
);

O2A1O1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1342),
.A2(n_1152),
.B(n_1163),
.C(n_1204),
.Y(n_1487)
);

AND2x2_ASAP7_75t_SL g1488 ( 
.A(n_1302),
.B(n_1245),
.Y(n_1488)
);

OR2x6_ASAP7_75t_L g1489 ( 
.A(n_1349),
.B(n_1229),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1300),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1324),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1393),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1325),
.A2(n_1169),
.B1(n_1280),
.B2(n_1244),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1303),
.B(n_1274),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1312),
.B(n_1274),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1372),
.A2(n_1249),
.B(n_1268),
.Y(n_1496)
);

O2A1O1Ixp33_ASAP7_75t_L g1497 ( 
.A1(n_1344),
.A2(n_1152),
.B(n_1205),
.C(n_1245),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1316),
.B(n_1187),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1372),
.A2(n_1268),
.B(n_1125),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1428),
.A2(n_1268),
.B(n_1125),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1346),
.A2(n_1338),
.B1(n_1332),
.B2(n_1326),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1327),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1328),
.A2(n_1278),
.B1(n_1268),
.B2(n_1279),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1365),
.B(n_1187),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1437),
.A2(n_1268),
.B(n_1125),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1438),
.A2(n_1142),
.B(n_1110),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1393),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1319),
.B(n_1187),
.Y(n_1508)
);

AO21x2_ASAP7_75t_L g1509 ( 
.A1(n_1427),
.A2(n_1140),
.B(n_1441),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1333),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1341),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1375),
.B(n_1292),
.Y(n_1512)
);

O2A1O1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1394),
.A2(n_1237),
.B(n_442),
.C(n_460),
.Y(n_1513)
);

O2A1O1Ixp5_ASAP7_75t_L g1514 ( 
.A1(n_1385),
.A2(n_1118),
.B(n_1146),
.C(n_1145),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1364),
.A2(n_1142),
.B(n_1110),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1334),
.A2(n_1278),
.B1(n_1285),
.B2(n_1279),
.Y(n_1516)
);

OAI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1446),
.A2(n_1285),
.B(n_1295),
.Y(n_1517)
);

BUFx4f_ASAP7_75t_L g1518 ( 
.A(n_1354),
.Y(n_1518)
);

NAND3xp33_ASAP7_75t_L g1519 ( 
.A(n_1394),
.B(n_1229),
.C(n_1182),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1357),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1392),
.A2(n_1142),
.B(n_1110),
.Y(n_1521)
);

O2A1O1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1352),
.A2(n_445),
.B(n_478),
.C(n_471),
.Y(n_1522)
);

OAI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1448),
.A2(n_1297),
.B(n_1296),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1336),
.B(n_1197),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1361),
.B(n_1197),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1410),
.B(n_1265),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1451),
.A2(n_1156),
.B(n_1147),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1396),
.A2(n_1156),
.B(n_1147),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1410),
.B(n_1449),
.Y(n_1529)
);

A2O1A1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1375),
.A2(n_1336),
.B(n_1352),
.C(n_1380),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_1353),
.B(n_1104),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1353),
.B(n_1104),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1408),
.A2(n_1156),
.B(n_1147),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1370),
.B(n_1384),
.Y(n_1534)
);

OAI21xp33_ASAP7_75t_L g1535 ( 
.A1(n_1370),
.A2(n_561),
.B(n_558),
.Y(n_1535)
);

OAI21xp33_ASAP7_75t_L g1536 ( 
.A1(n_1407),
.A2(n_563),
.B(n_562),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1393),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1318),
.B(n_1265),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1412),
.A2(n_1178),
.B(n_1172),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1452),
.B(n_1356),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1518),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_1463),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1483),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1481),
.B(n_1323),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1471),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1491),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1456),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1518),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1465),
.A2(n_1369),
.B(n_1366),
.Y(n_1549)
);

INVx5_ASAP7_75t_L g1550 ( 
.A(n_1458),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1512),
.B(n_1356),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1504),
.A2(n_1403),
.B1(n_1406),
.B2(n_1383),
.Y(n_1552)
);

OAI22x1_ASAP7_75t_L g1553 ( 
.A1(n_1460),
.A2(n_1351),
.B1(n_1405),
.B2(n_1383),
.Y(n_1553)
);

BUFx12f_ASAP7_75t_L g1554 ( 
.A(n_1457),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1530),
.A2(n_1350),
.B1(n_1318),
.B2(n_1345),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1454),
.A2(n_1376),
.B(n_1374),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_R g1557 ( 
.A(n_1457),
.B(n_1314),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1490),
.Y(n_1558)
);

A2O1A1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1534),
.A2(n_1513),
.B(n_1479),
.C(n_1522),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1529),
.B(n_1449),
.Y(n_1560)
);

INVx6_ASAP7_75t_L g1561 ( 
.A(n_1490),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1480),
.A2(n_1496),
.B(n_1468),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_SL g1563 ( 
.A(n_1459),
.B(n_1339),
.Y(n_1563)
);

NOR3xp33_ASAP7_75t_SL g1564 ( 
.A(n_1524),
.B(n_1382),
.C(n_1335),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1510),
.Y(n_1565)
);

O2A1O1Ixp33_ASAP7_75t_L g1566 ( 
.A1(n_1536),
.A2(n_1330),
.B(n_1409),
.C(n_1407),
.Y(n_1566)
);

NOR3xp33_ASAP7_75t_L g1567 ( 
.A(n_1501),
.B(n_1409),
.C(n_1444),
.Y(n_1567)
);

O2A1O1Ixp33_ASAP7_75t_L g1568 ( 
.A1(n_1535),
.A2(n_1450),
.B(n_1360),
.C(n_1348),
.Y(n_1568)
);

NOR2x1_ASAP7_75t_L g1569 ( 
.A(n_1519),
.B(n_1349),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1489),
.Y(n_1570)
);

OAI21xp33_ASAP7_75t_L g1571 ( 
.A1(n_1461),
.A2(n_1367),
.B(n_1362),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1477),
.B(n_1389),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1468),
.A2(n_1381),
.B(n_1379),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1515),
.A2(n_1387),
.B(n_1386),
.Y(n_1574)
);

A2O1A1Ixp33_ASAP7_75t_L g1575 ( 
.A1(n_1469),
.A2(n_1445),
.B(n_1377),
.C(n_1432),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_R g1576 ( 
.A(n_1490),
.B(n_1368),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1482),
.B(n_1431),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1525),
.A2(n_1420),
.B1(n_1418),
.B2(n_1442),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1497),
.B(n_1354),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1526),
.B(n_1390),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1498),
.A2(n_1406),
.B1(n_1403),
.B2(n_1423),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1462),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_SL g1583 ( 
.A(n_1508),
.B(n_1300),
.Y(n_1583)
);

INVx4_ASAP7_75t_L g1584 ( 
.A(n_1455),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1538),
.B(n_1425),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1455),
.B(n_1421),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_1455),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1487),
.B(n_1104),
.Y(n_1588)
);

A2O1A1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1476),
.A2(n_1359),
.B(n_1373),
.C(n_1423),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1488),
.B(n_1440),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1473),
.A2(n_1232),
.B(n_1202),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_1458),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1542),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1592),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1556),
.A2(n_1503),
.B(n_1464),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1562),
.A2(n_1503),
.B(n_1453),
.Y(n_1596)
);

AOI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1591),
.A2(n_1521),
.B(n_1467),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1540),
.B(n_1475),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1567),
.B(n_1458),
.Y(n_1599)
);

OAI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1551),
.A2(n_1559),
.B(n_1567),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1560),
.B(n_1475),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1571),
.A2(n_1474),
.B1(n_1435),
.B2(n_1340),
.C(n_1440),
.Y(n_1602)
);

OAI21x1_ASAP7_75t_L g1603 ( 
.A1(n_1549),
.A2(n_1466),
.B(n_1506),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1585),
.B(n_1475),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1587),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1561),
.Y(n_1606)
);

AOI211x1_ASAP7_75t_L g1607 ( 
.A1(n_1563),
.A2(n_1495),
.B(n_1494),
.C(n_1578),
.Y(n_1607)
);

AOI21xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1566),
.A2(n_1493),
.B(n_1486),
.Y(n_1608)
);

NAND3x1_ASAP7_75t_L g1609 ( 
.A(n_1569),
.B(n_1590),
.C(n_1577),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1574),
.A2(n_1527),
.B(n_1505),
.Y(n_1610)
);

HAxp5_ASAP7_75t_L g1611 ( 
.A(n_1553),
.B(n_564),
.CON(n_1611),
.SN(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1547),
.B(n_1489),
.Y(n_1612)
);

NAND2x1p5_ASAP7_75t_L g1613 ( 
.A(n_1550),
.B(n_1458),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1582),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1575),
.A2(n_1474),
.B(n_1493),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_SL g1616 ( 
.A(n_1568),
.B(n_571),
.C(n_569),
.Y(n_1616)
);

AOI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1588),
.A2(n_1532),
.B(n_1531),
.Y(n_1617)
);

OAI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1573),
.A2(n_1500),
.B(n_1517),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1580),
.B(n_1489),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1550),
.A2(n_1478),
.B(n_1470),
.Y(n_1620)
);

AO31x2_ASAP7_75t_L g1621 ( 
.A1(n_1589),
.A2(n_1486),
.A3(n_1516),
.B(n_1499),
.Y(n_1621)
);

OAI22x1_ASAP7_75t_L g1622 ( 
.A1(n_1579),
.A2(n_1426),
.B1(n_1265),
.B2(n_1485),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1572),
.B(n_1304),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1541),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1544),
.B(n_1421),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1547),
.B(n_1349),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1545),
.A2(n_1517),
.B(n_1523),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1550),
.A2(n_1470),
.B(n_1516),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1550),
.A2(n_1485),
.B(n_1523),
.Y(n_1629)
);

CKINVDCx20_ASAP7_75t_R g1630 ( 
.A(n_1557),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1543),
.Y(n_1631)
);

AOI21x1_ASAP7_75t_SL g1632 ( 
.A1(n_1586),
.A2(n_1397),
.B(n_1391),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1546),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1565),
.Y(n_1634)
);

AND2x2_ASAP7_75t_SL g1635 ( 
.A(n_1552),
.B(n_1592),
.Y(n_1635)
);

NAND3xp33_ASAP7_75t_L g1636 ( 
.A(n_1555),
.B(n_1395),
.C(n_1313),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1541),
.B(n_1421),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1570),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1586),
.B(n_1485),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1564),
.A2(n_1514),
.B(n_1528),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1542),
.A2(n_1564),
.B1(n_1581),
.B2(n_1541),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1541),
.B(n_1308),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1633),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1612),
.B(n_1583),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1593),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1634),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1608),
.A2(n_1628),
.B(n_1595),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1614),
.Y(n_1648)
);

NAND2x1p5_ASAP7_75t_L g1649 ( 
.A(n_1599),
.B(n_1485),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1597),
.A2(n_1539),
.B(n_1533),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1614),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1638),
.Y(n_1652)
);

INVx2_ASAP7_75t_SL g1653 ( 
.A(n_1606),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1606),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1627),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1600),
.B(n_1509),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1627),
.Y(n_1657)
);

O2A1O1Ixp33_ASAP7_75t_L g1658 ( 
.A1(n_1611),
.A2(n_480),
.B(n_489),
.C(n_481),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1626),
.B(n_542),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1610),
.A2(n_1507),
.B(n_1492),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1605),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1636),
.B(n_1548),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1618),
.Y(n_1663)
);

BUFx2_ASAP7_75t_L g1664 ( 
.A(n_1618),
.Y(n_1664)
);

AO21x2_ASAP7_75t_L g1665 ( 
.A1(n_1615),
.A2(n_1509),
.B(n_1140),
.Y(n_1665)
);

OAI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1602),
.A2(n_1548),
.B1(n_1554),
.B2(n_1492),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1619),
.Y(n_1667)
);

OAI21x1_ASAP7_75t_L g1668 ( 
.A1(n_1610),
.A2(n_1537),
.B(n_1507),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1601),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1616),
.A2(n_1599),
.B(n_1641),
.Y(n_1670)
);

INVx2_ASAP7_75t_SL g1671 ( 
.A(n_1594),
.Y(n_1671)
);

BUFx12f_ASAP7_75t_L g1672 ( 
.A(n_1631),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1598),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1621),
.Y(n_1674)
);

AOI21x1_ASAP7_75t_L g1675 ( 
.A1(n_1596),
.A2(n_1363),
.B(n_1416),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1607),
.A2(n_1548),
.B1(n_1433),
.B2(n_1434),
.Y(n_1676)
);

OAI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1640),
.A2(n_1439),
.B(n_506),
.Y(n_1677)
);

CKINVDCx16_ASAP7_75t_R g1678 ( 
.A(n_1630),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1604),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1623),
.Y(n_1680)
);

OAI21x1_ASAP7_75t_L g1681 ( 
.A1(n_1603),
.A2(n_1537),
.B(n_1182),
.Y(n_1681)
);

OAI21x1_ASAP7_75t_L g1682 ( 
.A1(n_1603),
.A2(n_1620),
.B(n_1629),
.Y(n_1682)
);

OAI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1617),
.A2(n_1184),
.B(n_1176),
.Y(n_1683)
);

OAI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1623),
.A2(n_481),
.B(n_480),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1625),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1632),
.A2(n_1184),
.B(n_1176),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1609),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1635),
.A2(n_1434),
.B1(n_1430),
.B2(n_1347),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1621),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1635),
.A2(n_1592),
.B(n_1232),
.Y(n_1690)
);

OAI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1609),
.A2(n_494),
.B(n_489),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_SL g1692 ( 
.A1(n_1611),
.A2(n_1337),
.B1(n_1443),
.B2(n_1413),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1621),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1631),
.Y(n_1694)
);

OAI21x1_ASAP7_75t_L g1695 ( 
.A1(n_1613),
.A2(n_1186),
.B(n_1178),
.Y(n_1695)
);

BUFx2_ASAP7_75t_L g1696 ( 
.A(n_1621),
.Y(n_1696)
);

OAI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1613),
.A2(n_1186),
.B(n_1178),
.Y(n_1697)
);

AOI22x1_ASAP7_75t_L g1698 ( 
.A1(n_1622),
.A2(n_514),
.B1(n_518),
.B2(n_494),
.Y(n_1698)
);

OAI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1594),
.A2(n_1181),
.B(n_1172),
.Y(n_1699)
);

OAI21x1_ASAP7_75t_L g1700 ( 
.A1(n_1594),
.A2(n_1181),
.B(n_1172),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1637),
.Y(n_1701)
);

BUFx2_ASAP7_75t_L g1702 ( 
.A(n_1605),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1637),
.B(n_1558),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1630),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1624),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1639),
.A2(n_1592),
.B(n_1232),
.Y(n_1706)
);

OA21x2_ASAP7_75t_L g1707 ( 
.A1(n_1639),
.A2(n_1430),
.B(n_570),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1624),
.Y(n_1708)
);

OAI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1624),
.A2(n_1548),
.B1(n_1584),
.B2(n_1561),
.Y(n_1709)
);

OAI21x1_ASAP7_75t_SL g1710 ( 
.A1(n_1642),
.A2(n_1584),
.B(n_1402),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1639),
.A2(n_1484),
.B1(n_1502),
.B2(n_1472),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1624),
.Y(n_1712)
);

OAI21x1_ASAP7_75t_SL g1713 ( 
.A1(n_1642),
.A2(n_1404),
.B(n_1399),
.Y(n_1713)
);

OAI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1600),
.A2(n_518),
.B(n_514),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1594),
.B(n_1111),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1639),
.Y(n_1716)
);

OAI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1600),
.A2(n_524),
.B(n_520),
.Y(n_1717)
);

AO21x2_ASAP7_75t_L g1718 ( 
.A1(n_1615),
.A2(n_1140),
.B(n_1411),
.Y(n_1718)
);

OAI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1597),
.A2(n_1192),
.B(n_1181),
.Y(n_1719)
);

BUFx8_ASAP7_75t_SL g1720 ( 
.A(n_1630),
.Y(n_1720)
);

OAI21x1_ASAP7_75t_SL g1721 ( 
.A1(n_1600),
.A2(n_1417),
.B(n_1414),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1633),
.Y(n_1722)
);

OAI21x1_ASAP7_75t_L g1723 ( 
.A1(n_1597),
.A2(n_1214),
.B(n_1192),
.Y(n_1723)
);

OAI21x1_ASAP7_75t_L g1724 ( 
.A1(n_1597),
.A2(n_1214),
.B(n_1192),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1600),
.A2(n_524),
.B(n_520),
.Y(n_1725)
);

OAI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1600),
.A2(n_1561),
.B1(n_530),
.B2(n_532),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1600),
.A2(n_532),
.B1(n_543),
.B2(n_530),
.C(n_526),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1633),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1670),
.B(n_1576),
.Y(n_1729)
);

OAI21x1_ASAP7_75t_L g1730 ( 
.A1(n_1719),
.A2(n_1217),
.B(n_1214),
.Y(n_1730)
);

OAI21x1_ASAP7_75t_L g1731 ( 
.A1(n_1719),
.A2(n_1220),
.B(n_1217),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1643),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1656),
.B(n_526),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1656),
.B(n_543),
.Y(n_1734)
);

OAI21x1_ASAP7_75t_L g1735 ( 
.A1(n_1723),
.A2(n_1220),
.B(n_1217),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1645),
.B(n_401),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1648),
.Y(n_1737)
);

INVx6_ASAP7_75t_L g1738 ( 
.A(n_1716),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1643),
.B(n_1728),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1647),
.A2(n_1232),
.B(n_1202),
.Y(n_1740)
);

AO31x2_ASAP7_75t_L g1741 ( 
.A1(n_1696),
.A2(n_1520),
.A3(n_1511),
.B(n_1398),
.Y(n_1741)
);

INVx3_ASAP7_75t_L g1742 ( 
.A(n_1654),
.Y(n_1742)
);

AOI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1682),
.A2(n_1232),
.B(n_1202),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1653),
.B(n_1709),
.Y(n_1744)
);

OAI21x1_ASAP7_75t_SL g1745 ( 
.A1(n_1714),
.A2(n_560),
.B(n_547),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1728),
.Y(n_1746)
);

CKINVDCx6p67_ASAP7_75t_R g1747 ( 
.A(n_1678),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1646),
.B(n_547),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1722),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1651),
.Y(n_1750)
);

A2O1A1Ixp33_ASAP7_75t_L g1751 ( 
.A1(n_1717),
.A2(n_554),
.B(n_589),
.C(n_570),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1685),
.B(n_560),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1652),
.Y(n_1753)
);

OR2x6_ASAP7_75t_L g1754 ( 
.A(n_1687),
.B(n_1447),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1673),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1696),
.B(n_576),
.Y(n_1756)
);

A2O1A1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1725),
.A2(n_554),
.B(n_617),
.C(n_589),
.Y(n_1757)
);

OA21x2_ASAP7_75t_L g1758 ( 
.A1(n_1682),
.A2(n_581),
.B(n_576),
.Y(n_1758)
);

OAI21x1_ASAP7_75t_L g1759 ( 
.A1(n_1723),
.A2(n_1235),
.B(n_1220),
.Y(n_1759)
);

BUFx12f_ASAP7_75t_L g1760 ( 
.A(n_1694),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1667),
.Y(n_1761)
);

AOI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1664),
.A2(n_1202),
.B(n_1201),
.Y(n_1762)
);

AOI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1664),
.A2(n_1202),
.B(n_1201),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1693),
.B(n_581),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1702),
.B(n_401),
.Y(n_1765)
);

INVxp67_ASAP7_75t_SL g1766 ( 
.A(n_1674),
.Y(n_1766)
);

CKINVDCx20_ASAP7_75t_R g1767 ( 
.A(n_1720),
.Y(n_1767)
);

OAI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1684),
.A2(n_1691),
.B(n_1677),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1669),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1679),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1726),
.A2(n_590),
.B(n_587),
.Y(n_1771)
);

OAI21x1_ASAP7_75t_SL g1772 ( 
.A1(n_1710),
.A2(n_590),
.B(n_587),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1674),
.B(n_592),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1644),
.Y(n_1774)
);

AOI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1690),
.A2(n_1201),
.B(n_1173),
.Y(n_1775)
);

OA21x2_ASAP7_75t_L g1776 ( 
.A1(n_1663),
.A2(n_596),
.B(n_592),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1644),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1701),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1704),
.B(n_1395),
.Y(n_1779)
);

INVx2_ASAP7_75t_SL g1780 ( 
.A(n_1661),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1663),
.A2(n_1201),
.B(n_1173),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1705),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1720),
.B(n_1413),
.Y(n_1783)
);

INVx3_ASAP7_75t_L g1784 ( 
.A(n_1654),
.Y(n_1784)
);

OA21x2_ASAP7_75t_L g1785 ( 
.A1(n_1724),
.A2(n_598),
.B(n_596),
.Y(n_1785)
);

OAI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1727),
.A2(n_602),
.B(n_598),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1649),
.A2(n_1201),
.B(n_1173),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1689),
.B(n_602),
.Y(n_1788)
);

OAI21x1_ASAP7_75t_SL g1789 ( 
.A1(n_1710),
.A2(n_605),
.B(n_603),
.Y(n_1789)
);

CKINVDCx20_ASAP7_75t_R g1790 ( 
.A(n_1694),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1689),
.B(n_603),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1702),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1672),
.Y(n_1793)
);

OAI21x1_ASAP7_75t_L g1794 ( 
.A1(n_1724),
.A2(n_1261),
.B(n_1235),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1655),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1659),
.B(n_605),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1659),
.B(n_629),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1657),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1708),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1680),
.A2(n_645),
.B1(n_658),
.B2(n_629),
.Y(n_1800)
);

AOI21x1_ASAP7_75t_L g1801 ( 
.A1(n_1662),
.A2(n_658),
.B(n_645),
.Y(n_1801)
);

BUFx3_ASAP7_75t_L g1802 ( 
.A(n_1661),
.Y(n_1802)
);

CKINVDCx11_ASAP7_75t_R g1803 ( 
.A(n_1672),
.Y(n_1803)
);

OA21x2_ASAP7_75t_L g1804 ( 
.A1(n_1650),
.A2(n_665),
.B(n_659),
.Y(n_1804)
);

OAI21x1_ASAP7_75t_L g1805 ( 
.A1(n_1650),
.A2(n_1681),
.B(n_1668),
.Y(n_1805)
);

BUFx3_ASAP7_75t_L g1806 ( 
.A(n_1653),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1712),
.Y(n_1807)
);

OA21x2_ASAP7_75t_L g1808 ( 
.A1(n_1681),
.A2(n_665),
.B(n_659),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1671),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1692),
.B(n_0),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1703),
.Y(n_1811)
);

OA21x2_ASAP7_75t_L g1812 ( 
.A1(n_1660),
.A2(n_1668),
.B(n_1683),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1671),
.B(n_463),
.Y(n_1813)
);

AOI21x1_ASAP7_75t_L g1814 ( 
.A1(n_1675),
.A2(n_617),
.B(n_688),
.Y(n_1814)
);

A2O1A1Ixp33_ASAP7_75t_L g1815 ( 
.A1(n_1658),
.A2(n_403),
.B(n_521),
.C(n_450),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1665),
.Y(n_1816)
);

AO31x2_ASAP7_75t_L g1817 ( 
.A1(n_1676),
.A2(n_1400),
.A3(n_1415),
.B(n_1401),
.Y(n_1817)
);

AND2x4_ASAP7_75t_SL g1818 ( 
.A(n_1716),
.B(n_1272),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1665),
.Y(n_1819)
);

A2O1A1Ixp33_ASAP7_75t_L g1820 ( 
.A1(n_1688),
.A2(n_403),
.B(n_521),
.C(n_450),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1665),
.Y(n_1821)
);

INVx2_ASAP7_75t_SL g1822 ( 
.A(n_1716),
.Y(n_1822)
);

INVx2_ASAP7_75t_SL g1823 ( 
.A(n_1716),
.Y(n_1823)
);

AO31x2_ASAP7_75t_L g1824 ( 
.A1(n_1706),
.A2(n_1429),
.A3(n_1436),
.B(n_1273),
.Y(n_1824)
);

INVx6_ASAP7_75t_L g1825 ( 
.A(n_1716),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1718),
.B(n_463),
.Y(n_1826)
);

O2A1O1Ixp33_ASAP7_75t_L g1827 ( 
.A1(n_1666),
.A2(n_537),
.B(n_549),
.C(n_495),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1698),
.A2(n_503),
.B1(n_512),
.B2(n_463),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1718),
.B(n_463),
.Y(n_1829)
);

AOI21x1_ASAP7_75t_L g1830 ( 
.A1(n_1675),
.A2(n_690),
.B(n_689),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1715),
.B(n_0),
.Y(n_1831)
);

OA21x2_ASAP7_75t_L g1832 ( 
.A1(n_1660),
.A2(n_537),
.B(n_495),
.Y(n_1832)
);

BUFx2_ASAP7_75t_SL g1833 ( 
.A(n_1715),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1683),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_1721),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1707),
.A2(n_889),
.B1(n_866),
.B2(n_1157),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1718),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1649),
.A2(n_1209),
.B(n_1173),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1649),
.A2(n_1209),
.B(n_1173),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1713),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1713),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1715),
.B(n_1),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1699),
.B(n_3),
.Y(n_1843)
);

OA21x2_ASAP7_75t_L g1844 ( 
.A1(n_1699),
.A2(n_549),
.B(n_537),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1707),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1686),
.Y(n_1846)
);

INVx3_ASAP7_75t_L g1847 ( 
.A(n_1695),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_SL g1848 ( 
.A(n_1721),
.B(n_866),
.Y(n_1848)
);

OAI21x1_ASAP7_75t_L g1849 ( 
.A1(n_1695),
.A2(n_1261),
.B(n_1235),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1700),
.B(n_6),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1707),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1686),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_SL g1853 ( 
.A1(n_1698),
.A2(n_549),
.B(n_521),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1700),
.B(n_463),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1697),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1697),
.Y(n_1856)
);

OAI21x1_ASAP7_75t_SL g1857 ( 
.A1(n_1711),
.A2(n_726),
.B(n_724),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1643),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1645),
.Y(n_1859)
);

OA21x2_ASAP7_75t_L g1860 ( 
.A1(n_1682),
.A2(n_731),
.B(n_727),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1647),
.A2(n_1209),
.B(n_1145),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1647),
.A2(n_1209),
.B(n_1145),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1656),
.B(n_463),
.Y(n_1863)
);

OAI21x1_ASAP7_75t_L g1864 ( 
.A1(n_1719),
.A2(n_1261),
.B(n_1419),
.Y(n_1864)
);

INVx2_ASAP7_75t_SL g1865 ( 
.A(n_1661),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1656),
.B(n_503),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1643),
.Y(n_1867)
);

OA21x2_ASAP7_75t_L g1868 ( 
.A1(n_1682),
.A2(n_737),
.B(n_732),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1648),
.Y(n_1869)
);

OA21x2_ASAP7_75t_L g1870 ( 
.A1(n_1682),
.A2(n_747),
.B(n_739),
.Y(n_1870)
);

AOI221xp5_ASAP7_75t_L g1871 ( 
.A1(n_1714),
.A2(n_577),
.B1(n_579),
.B2(n_575),
.C(n_573),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1648),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1656),
.B(n_503),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1688),
.A2(n_889),
.B1(n_866),
.B2(n_1158),
.Y(n_1874)
);

AOI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1647),
.A2(n_1209),
.B(n_1146),
.Y(n_1875)
);

OA21x2_ASAP7_75t_L g1876 ( 
.A1(n_1682),
.A2(n_750),
.B(n_748),
.Y(n_1876)
);

OAI21x1_ASAP7_75t_L g1877 ( 
.A1(n_1719),
.A2(n_1355),
.B(n_1273),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1648),
.Y(n_1878)
);

CKINVDCx14_ASAP7_75t_R g1879 ( 
.A(n_1694),
.Y(n_1879)
);

OR2x6_ASAP7_75t_L g1880 ( 
.A(n_1647),
.B(n_1272),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1732),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1859),
.B(n_503),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1737),
.Y(n_1883)
);

CKINVDCx20_ASAP7_75t_R g1884 ( 
.A(n_1767),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1869),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1739),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1792),
.B(n_503),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1739),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1778),
.B(n_503),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1753),
.B(n_512),
.Y(n_1890)
);

INVx3_ASAP7_75t_L g1891 ( 
.A(n_1738),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1746),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1872),
.Y(n_1893)
);

OA21x2_ASAP7_75t_L g1894 ( 
.A1(n_1837),
.A2(n_755),
.B(n_752),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1878),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1750),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1809),
.B(n_512),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1858),
.Y(n_1898)
);

AO31x2_ASAP7_75t_L g1899 ( 
.A1(n_1819),
.A2(n_1242),
.A3(n_1256),
.B(n_1241),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1867),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1755),
.B(n_512),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1795),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1749),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1768),
.A2(n_889),
.B1(n_866),
.B2(n_566),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1798),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1811),
.B(n_512),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1733),
.B(n_512),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1777),
.Y(n_1908)
);

AO21x2_ASAP7_75t_L g1909 ( 
.A1(n_1826),
.A2(n_757),
.B(n_756),
.Y(n_1909)
);

OAI21x1_ASAP7_75t_L g1910 ( 
.A1(n_1740),
.A2(n_1266),
.B(n_1259),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1761),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1769),
.Y(n_1912)
);

BUFx2_ASAP7_75t_L g1913 ( 
.A(n_1742),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1770),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1782),
.Y(n_1915)
);

INVx3_ASAP7_75t_L g1916 ( 
.A(n_1738),
.Y(n_1916)
);

INVxp67_ASAP7_75t_L g1917 ( 
.A(n_1780),
.Y(n_1917)
);

AO21x2_ASAP7_75t_L g1918 ( 
.A1(n_1826),
.A2(n_1270),
.B(n_1194),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1756),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1741),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1799),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1742),
.B(n_8),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1756),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1741),
.Y(n_1924)
);

BUFx4f_ASAP7_75t_L g1925 ( 
.A(n_1747),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1741),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1733),
.B(n_580),
.Y(n_1927)
);

BUFx3_ASAP7_75t_L g1928 ( 
.A(n_1802),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1773),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1773),
.Y(n_1930)
);

BUFx6f_ASAP7_75t_L g1931 ( 
.A(n_1754),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1807),
.Y(n_1932)
);

BUFx3_ASAP7_75t_L g1933 ( 
.A(n_1803),
.Y(n_1933)
);

HB1xp67_ASAP7_75t_L g1934 ( 
.A(n_1806),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1788),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1788),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1774),
.B(n_8),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1791),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1784),
.B(n_9),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1791),
.Y(n_1940)
);

OAI21x1_ASAP7_75t_L g1941 ( 
.A1(n_1743),
.A2(n_1212),
.B(n_1189),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1784),
.B(n_9),
.Y(n_1942)
);

OR2x6_ASAP7_75t_L g1943 ( 
.A(n_1880),
.B(n_1272),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1734),
.B(n_582),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1764),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1865),
.B(n_10),
.Y(n_1946)
);

INVx2_ASAP7_75t_SL g1947 ( 
.A(n_1738),
.Y(n_1947)
);

AO21x1_ASAP7_75t_SL g1948 ( 
.A1(n_1835),
.A2(n_1841),
.B(n_1840),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1822),
.B(n_10),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1760),
.Y(n_1950)
);

INVx2_ASAP7_75t_SL g1951 ( 
.A(n_1825),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1823),
.B(n_11),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1855),
.B(n_13),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1764),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1734),
.Y(n_1955)
);

AO21x1_ASAP7_75t_SL g1956 ( 
.A1(n_1854),
.A2(n_1846),
.B(n_1856),
.Y(n_1956)
);

AOI22xp33_ASAP7_75t_SL g1957 ( 
.A1(n_1776),
.A2(n_1810),
.B1(n_1829),
.B2(n_1789),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1825),
.B(n_13),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1863),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1863),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1866),
.B(n_15),
.Y(n_1961)
);

OAI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1800),
.A2(n_585),
.B(n_583),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1866),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1873),
.Y(n_1964)
);

AO21x2_ASAP7_75t_L g1965 ( 
.A1(n_1829),
.A2(n_1223),
.B(n_1212),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1873),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1845),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1729),
.A2(n_595),
.B1(n_597),
.B2(n_594),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1825),
.B(n_1846),
.Y(n_1969)
);

HB1xp67_ASAP7_75t_L g1970 ( 
.A(n_1736),
.Y(n_1970)
);

INVx2_ASAP7_75t_SL g1971 ( 
.A(n_1736),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1754),
.B(n_15),
.Y(n_1972)
);

BUFx5_ASAP7_75t_L g1973 ( 
.A(n_1813),
.Y(n_1973)
);

HB1xp67_ASAP7_75t_L g1974 ( 
.A(n_1765),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1847),
.B(n_16),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1847),
.B(n_18),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1748),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1880),
.B(n_18),
.Y(n_1978)
);

OAI21x1_ASAP7_75t_L g1979 ( 
.A1(n_1743),
.A2(n_1231),
.B(n_1223),
.Y(n_1979)
);

OA21x2_ASAP7_75t_L g1980 ( 
.A1(n_1805),
.A2(n_839),
.B(n_838),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1748),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1880),
.B(n_19),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1796),
.B(n_20),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1776),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1854),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1824),
.Y(n_1986)
);

AND2x4_ASAP7_75t_L g1987 ( 
.A(n_1754),
.B(n_21),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1851),
.Y(n_1988)
);

INVx3_ASAP7_75t_L g1989 ( 
.A(n_1812),
.Y(n_1989)
);

HB1xp67_ASAP7_75t_L g1990 ( 
.A(n_1765),
.Y(n_1990)
);

HB1xp67_ASAP7_75t_L g1991 ( 
.A(n_1758),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1816),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1796),
.B(n_21),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1752),
.Y(n_1994)
);

INVx2_ASAP7_75t_SL g1995 ( 
.A(n_1744),
.Y(n_1995)
);

OA21x2_ASAP7_75t_L g1996 ( 
.A1(n_1821),
.A2(n_839),
.B(n_838),
.Y(n_1996)
);

INVx3_ASAP7_75t_L g1997 ( 
.A(n_1812),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1752),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1834),
.B(n_22),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1766),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1797),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1801),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1797),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1824),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1824),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_1793),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1766),
.Y(n_2007)
);

AO21x2_ASAP7_75t_L g2008 ( 
.A1(n_1781),
.A2(n_1234),
.B(n_1231),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1852),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1758),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1804),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1804),
.Y(n_2012)
);

INVx3_ASAP7_75t_L g2013 ( 
.A(n_1860),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1817),
.Y(n_2014)
);

INVx2_ASAP7_75t_SL g2015 ( 
.A(n_1848),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1833),
.B(n_24),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1817),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1817),
.Y(n_2018)
);

BUFx3_ASAP7_75t_L g2019 ( 
.A(n_1790),
.Y(n_2019)
);

OAI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1800),
.A2(n_1815),
.B(n_1757),
.Y(n_2020)
);

HB1xp67_ASAP7_75t_L g2021 ( 
.A(n_1785),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1843),
.B(n_601),
.Y(n_2022)
);

BUFx6f_ASAP7_75t_L g2023 ( 
.A(n_1785),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_1850),
.Y(n_2024)
);

HB1xp67_ASAP7_75t_L g2025 ( 
.A(n_1808),
.Y(n_2025)
);

HB1xp67_ASAP7_75t_L g2026 ( 
.A(n_1808),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1860),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1868),
.Y(n_2028)
);

NAND3xp33_ASAP7_75t_L g2029 ( 
.A(n_1901),
.B(n_1820),
.C(n_1771),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_2024),
.A2(n_1871),
.B1(n_1772),
.B2(n_1874),
.Y(n_2030)
);

OAI21x1_ASAP7_75t_L g2031 ( 
.A1(n_1989),
.A2(n_1997),
.B(n_1882),
.Y(n_2031)
);

AOI211xp5_ASAP7_75t_L g2032 ( 
.A1(n_2022),
.A2(n_1871),
.B(n_1827),
.C(n_1842),
.Y(n_2032)
);

AO21x2_ASAP7_75t_L g2033 ( 
.A1(n_1889),
.A2(n_1781),
.B(n_1763),
.Y(n_2033)
);

OA21x2_ASAP7_75t_L g2034 ( 
.A1(n_2000),
.A2(n_2007),
.B(n_1992),
.Y(n_2034)
);

OAI211xp5_ASAP7_75t_L g2035 ( 
.A1(n_2020),
.A2(n_1786),
.B(n_1831),
.C(n_1751),
.Y(n_2035)
);

AOI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_1995),
.A2(n_1828),
.B1(n_1779),
.B2(n_1783),
.Y(n_2036)
);

OAI211xp5_ASAP7_75t_SL g2037 ( 
.A1(n_1983),
.A2(n_1879),
.B(n_1827),
.C(n_1853),
.Y(n_2037)
);

INVx2_ASAP7_75t_SL g2038 ( 
.A(n_1933),
.Y(n_2038)
);

OR2x2_ASAP7_75t_L g2039 ( 
.A(n_1921),
.B(n_1762),
.Y(n_2039)
);

AOI22xp33_ASAP7_75t_L g2040 ( 
.A1(n_1957),
.A2(n_1857),
.B1(n_1745),
.B2(n_1828),
.Y(n_2040)
);

AOI22xp33_ASAP7_75t_L g2041 ( 
.A1(n_2002),
.A2(n_1836),
.B1(n_1844),
.B2(n_1832),
.Y(n_2041)
);

INVx3_ASAP7_75t_L g2042 ( 
.A(n_1928),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1913),
.B(n_1762),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_1887),
.Y(n_2044)
);

OAI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_1995),
.A2(n_1861),
.B1(n_1875),
.B2(n_1862),
.Y(n_2045)
);

AOI221xp5_ASAP7_75t_L g2046 ( 
.A1(n_1927),
.A2(n_1944),
.B1(n_1962),
.B2(n_1981),
.C(n_1983),
.Y(n_2046)
);

INVx3_ASAP7_75t_L g2047 ( 
.A(n_1928),
.Y(n_2047)
);

AOI221xp5_ASAP7_75t_L g2048 ( 
.A1(n_1981),
.A2(n_616),
.B1(n_619),
.B2(n_613),
.C(n_611),
.Y(n_2048)
);

NAND2x1p5_ASAP7_75t_L g2049 ( 
.A(n_1972),
.B(n_1832),
.Y(n_2049)
);

AOI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_2002),
.A2(n_1844),
.B1(n_1870),
.B2(n_1868),
.Y(n_2050)
);

OAI21x1_ASAP7_75t_L g2051 ( 
.A1(n_1989),
.A2(n_1763),
.B(n_1814),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1890),
.Y(n_2052)
);

AOI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_1972),
.A2(n_1876),
.B1(n_1870),
.B2(n_1818),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1898),
.Y(n_2054)
);

AOI22xp33_ASAP7_75t_L g2055 ( 
.A1(n_2002),
.A2(n_1876),
.B1(n_566),
.B2(n_606),
.Y(n_2055)
);

OAI22xp5_ASAP7_75t_L g2056 ( 
.A1(n_1978),
.A2(n_1861),
.B1(n_1875),
.B2(n_1862),
.Y(n_2056)
);

AOI22xp33_ASAP7_75t_L g2057 ( 
.A1(n_2002),
.A2(n_566),
.B1(n_606),
.B2(n_450),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_L g2058 ( 
.A(n_1933),
.B(n_24),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1898),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_1919),
.B(n_1877),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1881),
.Y(n_2061)
);

AOI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_1972),
.A2(n_1775),
.B1(n_623),
.B2(n_588),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1881),
.Y(n_2063)
);

OAI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_1978),
.A2(n_1775),
.B(n_1787),
.Y(n_2064)
);

OAI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_1982),
.A2(n_1838),
.B1(n_1839),
.B2(n_1787),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_SL g2066 ( 
.A1(n_1987),
.A2(n_623),
.B1(n_588),
.B2(n_621),
.Y(n_2066)
);

OAI31xp33_ASAP7_75t_L g2067 ( 
.A1(n_1987),
.A2(n_655),
.A3(n_606),
.B(n_441),
.Y(n_2067)
);

AOI222xp33_ASAP7_75t_L g2068 ( 
.A1(n_1955),
.A2(n_623),
.B1(n_588),
.B2(n_655),
.C1(n_626),
.C2(n_622),
.Y(n_2068)
);

OAI21x1_ASAP7_75t_L g2069 ( 
.A1(n_1989),
.A2(n_1830),
.B(n_1731),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_2002),
.A2(n_655),
.B1(n_889),
.B2(n_866),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1890),
.Y(n_2071)
);

AO21x2_ASAP7_75t_L g2072 ( 
.A1(n_1906),
.A2(n_1864),
.B(n_1735),
.Y(n_2072)
);

AOI22xp33_ASAP7_75t_L g2073 ( 
.A1(n_1935),
.A2(n_889),
.B1(n_623),
.B2(n_1247),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1915),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1892),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_1884),
.B(n_25),
.Y(n_2076)
);

OAI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_1982),
.A2(n_1839),
.B1(n_1838),
.B2(n_632),
.Y(n_2077)
);

AOI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_1935),
.A2(n_1247),
.B1(n_1246),
.B2(n_1234),
.Y(n_2078)
);

AOI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_1936),
.A2(n_1247),
.B1(n_1248),
.B2(n_1246),
.Y(n_2079)
);

AOI22xp33_ASAP7_75t_L g2080 ( 
.A1(n_1936),
.A2(n_1247),
.B1(n_1269),
.B2(n_1248),
.Y(n_2080)
);

AND2x4_ASAP7_75t_L g2081 ( 
.A(n_1934),
.B(n_1913),
.Y(n_2081)
);

OAI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_1961),
.A2(n_635),
.B1(n_639),
.B2(n_620),
.Y(n_2082)
);

AOI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_1987),
.A2(n_1247),
.B1(n_559),
.B2(n_642),
.Y(n_2083)
);

OAI22xp5_ASAP7_75t_L g2084 ( 
.A1(n_1993),
.A2(n_644),
.B1(n_646),
.B2(n_641),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1892),
.Y(n_2085)
);

AOI222xp33_ASAP7_75t_L g2086 ( 
.A1(n_2001),
.A2(n_653),
.B1(n_649),
.B2(n_654),
.C1(n_652),
.C2(n_648),
.Y(n_2086)
);

AOI21xp5_ASAP7_75t_L g2087 ( 
.A1(n_1943),
.A2(n_1849),
.B(n_1759),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1947),
.B(n_1730),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1900),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1915),
.Y(n_2090)
);

AOI21xp33_ASAP7_75t_L g2091 ( 
.A1(n_1964),
.A2(n_657),
.B(n_656),
.Y(n_2091)
);

INVx1_ASAP7_75t_SL g2092 ( 
.A(n_1884),
.Y(n_2092)
);

OAI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_1993),
.A2(n_663),
.B1(n_664),
.B2(n_662),
.Y(n_2093)
);

OAI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_1961),
.A2(n_559),
.B1(n_553),
.B2(n_461),
.Y(n_2094)
);

OAI222xp33_ASAP7_75t_L g2095 ( 
.A1(n_1937),
.A2(n_369),
.B1(n_366),
.B2(n_363),
.C1(n_365),
.C2(n_360),
.Y(n_2095)
);

OAI221xp5_ASAP7_75t_L g2096 ( 
.A1(n_1904),
.A2(n_553),
.B1(n_875),
.B2(n_850),
.C(n_400),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1902),
.Y(n_2097)
);

OAI211xp5_ASAP7_75t_L g2098 ( 
.A1(n_1999),
.A2(n_32),
.B(n_25),
.C(n_28),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1902),
.Y(n_2099)
);

NOR2x1_ASAP7_75t_SL g2100 ( 
.A(n_1948),
.B(n_553),
.Y(n_2100)
);

AOI22xp33_ASAP7_75t_L g2101 ( 
.A1(n_2003),
.A2(n_1247),
.B1(n_1269),
.B2(n_1158),
.Y(n_2101)
);

BUFx2_ASAP7_75t_L g2102 ( 
.A(n_1891),
.Y(n_2102)
);

OAI221xp5_ASAP7_75t_L g2103 ( 
.A1(n_1968),
.A2(n_553),
.B1(n_875),
.B2(n_850),
.C(n_404),
.Y(n_2103)
);

OAI22xp33_ASAP7_75t_SL g2104 ( 
.A1(n_1937),
.A2(n_1998),
.B1(n_1994),
.B2(n_1919),
.Y(n_2104)
);

AOI22xp33_ASAP7_75t_L g2105 ( 
.A1(n_1923),
.A2(n_1161),
.B1(n_1166),
.B2(n_1160),
.Y(n_2105)
);

AOI222xp33_ASAP7_75t_L g2106 ( 
.A1(n_1923),
.A2(n_371),
.B1(n_373),
.B2(n_407),
.C1(n_416),
.C2(n_417),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_1897),
.B(n_1794),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1905),
.Y(n_2108)
);

AOI21xp5_ASAP7_75t_L g2109 ( 
.A1(n_1943),
.A2(n_2008),
.B(n_1991),
.Y(n_2109)
);

OA21x2_ASAP7_75t_L g2110 ( 
.A1(n_2000),
.A2(n_1161),
.B(n_1160),
.Y(n_2110)
);

BUFx3_ASAP7_75t_L g2111 ( 
.A(n_2019),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1900),
.Y(n_2112)
);

AO31x2_ASAP7_75t_L g2113 ( 
.A1(n_2014),
.A2(n_1174),
.A3(n_1166),
.B(n_1118),
.Y(n_2113)
);

AOI22xp33_ASAP7_75t_SL g2114 ( 
.A1(n_2023),
.A2(n_628),
.B1(n_896),
.B2(n_870),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1905),
.Y(n_2115)
);

NAND3xp33_ASAP7_75t_L g2116 ( 
.A(n_1964),
.B(n_837),
.C(n_1272),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1896),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1947),
.B(n_28),
.Y(n_2118)
);

CKINVDCx5p33_ASAP7_75t_R g2119 ( 
.A(n_2006),
.Y(n_2119)
);

AOI22xp33_ASAP7_75t_L g2120 ( 
.A1(n_1929),
.A2(n_1174),
.B1(n_837),
.B2(n_628),
.Y(n_2120)
);

AND2x6_ASAP7_75t_L g2121 ( 
.A(n_2016),
.B(n_1272),
.Y(n_2121)
);

OAI21x1_ASAP7_75t_SL g2122 ( 
.A1(n_1903),
.A2(n_33),
.B(n_34),
.Y(n_2122)
);

AOI211xp5_ASAP7_75t_L g2123 ( 
.A1(n_1999),
.A2(n_37),
.B(n_33),
.C(n_35),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1896),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1886),
.Y(n_2125)
);

AOI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_1929),
.A2(n_628),
.B1(n_1116),
.B2(n_1104),
.Y(n_2126)
);

AOI22xp33_ASAP7_75t_L g2127 ( 
.A1(n_1930),
.A2(n_628),
.B1(n_1116),
.B2(n_1104),
.Y(n_2127)
);

OAI22xp33_ASAP7_75t_L g2128 ( 
.A1(n_2023),
.A2(n_424),
.B1(n_425),
.B2(n_418),
.Y(n_2128)
);

INVx3_ASAP7_75t_L g2129 ( 
.A(n_1891),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1887),
.Y(n_2130)
);

OAI221xp5_ASAP7_75t_L g2131 ( 
.A1(n_1977),
.A2(n_451),
.B1(n_468),
.B2(n_435),
.C(n_426),
.Y(n_2131)
);

AO21x2_ASAP7_75t_L g2132 ( 
.A1(n_1986),
.A2(n_2005),
.B(n_2004),
.Y(n_2132)
);

OA21x2_ASAP7_75t_L g2133 ( 
.A1(n_2007),
.A2(n_475),
.B(n_472),
.Y(n_2133)
);

OAI21x1_ASAP7_75t_L g2134 ( 
.A1(n_1997),
.A2(n_35),
.B(n_39),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1888),
.B(n_39),
.Y(n_2135)
);

AOI221xp5_ASAP7_75t_SL g2136 ( 
.A1(n_1917),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.C(n_46),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_1951),
.B(n_40),
.Y(n_2137)
);

OAI22xp33_ASAP7_75t_L g2138 ( 
.A1(n_2023),
.A2(n_1971),
.B1(n_1990),
.B2(n_1974),
.Y(n_2138)
);

HB1xp67_ASAP7_75t_L g2139 ( 
.A(n_1932),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1883),
.Y(n_2140)
);

OAI22xp33_ASAP7_75t_L g2141 ( 
.A1(n_2023),
.A2(n_492),
.B1(n_497),
.B2(n_479),
.Y(n_2141)
);

OAI22xp33_ASAP7_75t_L g2142 ( 
.A1(n_2023),
.A2(n_500),
.B1(n_523),
.B2(n_499),
.Y(n_2142)
);

AOI22xp33_ASAP7_75t_L g2143 ( 
.A1(n_1930),
.A2(n_628),
.B1(n_1116),
.B2(n_1185),
.Y(n_2143)
);

AOI21xp33_ASAP7_75t_L g2144 ( 
.A1(n_1966),
.A2(n_41),
.B(n_42),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1883),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1911),
.Y(n_2146)
);

HB1xp67_ASAP7_75t_L g2147 ( 
.A(n_1997),
.Y(n_2147)
);

OA21x2_ASAP7_75t_L g2148 ( 
.A1(n_1992),
.A2(n_538),
.B(n_535),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_1897),
.B(n_48),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1911),
.Y(n_2150)
);

INVx4_ASAP7_75t_L g2151 ( 
.A(n_1950),
.Y(n_2151)
);

AOI221xp5_ASAP7_75t_L g2152 ( 
.A1(n_1945),
.A2(n_555),
.B1(n_556),
.B2(n_545),
.C(n_540),
.Y(n_2152)
);

AOI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_1938),
.A2(n_628),
.B1(n_1251),
.B2(n_1185),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_1951),
.B(n_48),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1912),
.Y(n_2155)
);

OA21x2_ASAP7_75t_L g2156 ( 
.A1(n_2014),
.A2(n_584),
.B(n_574),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1912),
.Y(n_2157)
);

AOI22xp33_ASAP7_75t_SL g2158 ( 
.A1(n_2021),
.A2(n_628),
.B1(n_599),
.B2(n_600),
.Y(n_2158)
);

AOI22xp33_ASAP7_75t_L g2159 ( 
.A1(n_1938),
.A2(n_628),
.B1(n_1116),
.B2(n_1185),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_1891),
.B(n_50),
.Y(n_2160)
);

CKINVDCx5p33_ASAP7_75t_R g2161 ( 
.A(n_2006),
.Y(n_2161)
);

BUFx3_ASAP7_75t_L g2162 ( 
.A(n_2019),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1885),
.Y(n_2163)
);

AOI221xp5_ASAP7_75t_L g2164 ( 
.A1(n_1945),
.A2(n_608),
.B1(n_609),
.B2(n_607),
.C(n_593),
.Y(n_2164)
);

HB1xp67_ASAP7_75t_L g2165 ( 
.A(n_1914),
.Y(n_2165)
);

INVx3_ASAP7_75t_L g2166 ( 
.A(n_1916),
.Y(n_2166)
);

OAI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_1925),
.A2(n_614),
.B1(n_615),
.B2(n_610),
.Y(n_2167)
);

AOI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_1943),
.A2(n_1146),
.B(n_1118),
.Y(n_2168)
);

AOI221xp5_ASAP7_75t_L g2169 ( 
.A1(n_1954),
.A2(n_638),
.B1(n_637),
.B2(n_634),
.C(n_624),
.Y(n_2169)
);

BUFx3_ASAP7_75t_L g2170 ( 
.A(n_1950),
.Y(n_2170)
);

AOI22xp33_ASAP7_75t_L g2171 ( 
.A1(n_1940),
.A2(n_628),
.B1(n_1116),
.B2(n_1185),
.Y(n_2171)
);

AOI22xp33_ASAP7_75t_L g2172 ( 
.A1(n_1940),
.A2(n_1251),
.B1(n_1185),
.B2(n_1165),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_1916),
.B(n_50),
.Y(n_2173)
);

OAI211xp5_ASAP7_75t_L g2174 ( 
.A1(n_2016),
.A2(n_55),
.B(n_51),
.C(n_54),
.Y(n_2174)
);

OR2x2_ASAP7_75t_L g2175 ( 
.A(n_1908),
.B(n_51),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1914),
.Y(n_2176)
);

OAI22xp5_ASAP7_75t_L g2177 ( 
.A1(n_1925),
.A2(n_618),
.B1(n_1195),
.B2(n_1154),
.Y(n_2177)
);

NAND3xp33_ASAP7_75t_L g2178 ( 
.A(n_1966),
.B(n_1195),
.C(n_1154),
.Y(n_2178)
);

AOI22xp33_ASAP7_75t_SL g2179 ( 
.A1(n_2025),
.A2(n_1144),
.B1(n_56),
.B2(n_54),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1959),
.Y(n_2180)
);

AOI21x1_ASAP7_75t_L g2181 ( 
.A1(n_1907),
.A2(n_55),
.B(n_57),
.Y(n_2181)
);

OA21x2_ASAP7_75t_L g2182 ( 
.A1(n_2017),
.A2(n_59),
.B(n_60),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2081),
.B(n_1916),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2165),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2165),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2146),
.Y(n_2186)
);

OR2x2_ASAP7_75t_L g2187 ( 
.A(n_2044),
.B(n_1985),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2081),
.B(n_1969),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2102),
.B(n_1969),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2034),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2150),
.Y(n_2191)
);

INVxp67_ASAP7_75t_L g2192 ( 
.A(n_2044),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2129),
.B(n_1948),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2034),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2155),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2157),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2176),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2129),
.B(n_1956),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2166),
.B(n_1956),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2166),
.B(n_2042),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2061),
.Y(n_2201)
);

INVx3_ASAP7_75t_L g2202 ( 
.A(n_2043),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2042),
.B(n_1970),
.Y(n_2203)
);

AND2x4_ASAP7_75t_L g2204 ( 
.A(n_2031),
.B(n_1975),
.Y(n_2204)
);

OR2x2_ASAP7_75t_L g2205 ( 
.A(n_2139),
.B(n_2039),
.Y(n_2205)
);

OAI22xp5_ASAP7_75t_L g2206 ( 
.A1(n_2123),
.A2(n_1925),
.B1(n_2015),
.B2(n_1971),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2139),
.B(n_1953),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2063),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2132),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2180),
.B(n_1953),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2075),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_2151),
.B(n_1946),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2047),
.B(n_1973),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2047),
.B(n_1973),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2085),
.Y(n_2215)
);

OR2x2_ASAP7_75t_L g2216 ( 
.A(n_2125),
.B(n_1985),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2132),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2182),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_2182),
.Y(n_2219)
);

NOR2xp33_ASAP7_75t_L g2220 ( 
.A(n_2151),
.B(n_1946),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2060),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2089),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2112),
.Y(n_2223)
);

OAI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_2098),
.A2(n_2015),
.B1(n_1939),
.B2(n_1942),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2046),
.B(n_1975),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2046),
.B(n_2130),
.Y(n_2226)
);

INVx2_ASAP7_75t_SL g2227 ( 
.A(n_2111),
.Y(n_2227)
);

INVxp33_ASAP7_75t_L g2228 ( 
.A(n_2100),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2115),
.Y(n_2229)
);

AND2x4_ASAP7_75t_L g2230 ( 
.A(n_2064),
.B(n_1976),
.Y(n_2230)
);

AOI22xp33_ASAP7_75t_L g2231 ( 
.A1(n_2156),
.A2(n_1909),
.B1(n_1984),
.B2(n_1954),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2088),
.B(n_1973),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2104),
.B(n_1976),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2135),
.B(n_1960),
.Y(n_2234)
);

OR2x6_ASAP7_75t_L g2235 ( 
.A(n_2049),
.B(n_1943),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2147),
.Y(n_2236)
);

OR2x2_ASAP7_75t_L g2237 ( 
.A(n_2054),
.B(n_1963),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2117),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2147),
.Y(n_2239)
);

INVx2_ASAP7_75t_SL g2240 ( 
.A(n_2162),
.Y(n_2240)
);

NAND2x1p5_ASAP7_75t_SL g2241 ( 
.A(n_2038),
.B(n_2160),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2107),
.B(n_1973),
.Y(n_2242)
);

NOR2xp67_ASAP7_75t_L g2243 ( 
.A(n_2119),
.B(n_2026),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2124),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2059),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2107),
.B(n_1973),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2052),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2118),
.B(n_1973),
.Y(n_2248)
);

BUFx3_ASAP7_75t_L g2249 ( 
.A(n_2170),
.Y(n_2249)
);

HB1xp67_ASAP7_75t_L g2250 ( 
.A(n_2175),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2071),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2121),
.B(n_1922),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2097),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2137),
.B(n_1973),
.Y(n_2254)
);

AND2x4_ASAP7_75t_L g2255 ( 
.A(n_2121),
.B(n_1922),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_2099),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2154),
.B(n_1973),
.Y(n_2257)
);

OR2x2_ASAP7_75t_L g2258 ( 
.A(n_2108),
.B(n_2010),
.Y(n_2258)
);

BUFx6f_ASAP7_75t_L g2259 ( 
.A(n_2181),
.Y(n_2259)
);

AOI22xp33_ASAP7_75t_L g2260 ( 
.A1(n_2156),
.A2(n_2133),
.B1(n_2148),
.B2(n_2094),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2074),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2092),
.B(n_1939),
.Y(n_2262)
);

BUFx2_ASAP7_75t_L g2263 ( 
.A(n_2161),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2173),
.B(n_1942),
.Y(n_2264)
);

HB1xp67_ASAP7_75t_L g2265 ( 
.A(n_2133),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2090),
.Y(n_2266)
);

OR2x2_ASAP7_75t_L g2267 ( 
.A(n_2138),
.B(n_2010),
.Y(n_2267)
);

AND2x4_ASAP7_75t_L g2268 ( 
.A(n_2121),
.B(n_2109),
.Y(n_2268)
);

AND2x4_ASAP7_75t_L g2269 ( 
.A(n_2121),
.B(n_1958),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2140),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_2145),
.Y(n_2271)
);

AND2x4_ASAP7_75t_SL g2272 ( 
.A(n_2149),
.B(n_1958),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2058),
.B(n_2065),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2163),
.Y(n_2274)
);

AOI22xp33_ASAP7_75t_L g2275 ( 
.A1(n_2148),
.A2(n_1909),
.B1(n_1984),
.B2(n_2011),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2110),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2121),
.B(n_1949),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2069),
.B(n_1949),
.Y(n_2278)
);

OR2x2_ASAP7_75t_L g2279 ( 
.A(n_2138),
.B(n_1885),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2149),
.B(n_1952),
.Y(n_2280)
);

HB1xp67_ASAP7_75t_L g2281 ( 
.A(n_2134),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2036),
.B(n_1952),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2110),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2178),
.Y(n_2284)
);

OAI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_2098),
.A2(n_1931),
.B1(n_2013),
.B2(n_2009),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2056),
.B(n_1931),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2049),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2076),
.B(n_2033),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2113),
.Y(n_2289)
);

AOI22xp33_ASAP7_75t_L g2290 ( 
.A1(n_2094),
.A2(n_1909),
.B1(n_2012),
.B2(n_2011),
.Y(n_2290)
);

AND2x4_ASAP7_75t_L g2291 ( 
.A(n_2109),
.B(n_2013),
.Y(n_2291)
);

INVx4_ASAP7_75t_L g2292 ( 
.A(n_2136),
.Y(n_2292)
);

HB1xp67_ASAP7_75t_L g2293 ( 
.A(n_2072),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2033),
.B(n_1931),
.Y(n_2294)
);

AND2x4_ASAP7_75t_L g2295 ( 
.A(n_2072),
.B(n_2013),
.Y(n_2295)
);

AND2x4_ASAP7_75t_L g2296 ( 
.A(n_2051),
.B(n_1931),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2087),
.B(n_1931),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2082),
.B(n_2009),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_2087),
.B(n_1893),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2122),
.Y(n_2300)
);

NOR2x1_ASAP7_75t_R g2301 ( 
.A(n_2066),
.B(n_2174),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2045),
.B(n_1893),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2035),
.A2(n_2012),
.B1(n_1988),
.B2(n_1967),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2053),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2082),
.B(n_1895),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2113),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2113),
.Y(n_2307)
);

NAND2x1p5_ASAP7_75t_SL g2308 ( 
.A(n_2174),
.B(n_2028),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2202),
.B(n_2084),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2202),
.B(n_2188),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2202),
.B(n_2188),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_2200),
.B(n_2093),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2186),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2288),
.B(n_2086),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2191),
.Y(n_2315)
);

OA21x2_ASAP7_75t_L g2316 ( 
.A1(n_2218),
.A2(n_2018),
.B(n_2017),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2190),
.Y(n_2317)
);

AND2x4_ASAP7_75t_L g2318 ( 
.A(n_2235),
.B(n_2062),
.Y(n_2318)
);

INVx3_ASAP7_75t_L g2319 ( 
.A(n_2295),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2195),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2288),
.B(n_2032),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2196),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2200),
.B(n_2077),
.Y(n_2323)
);

OR2x2_ASAP7_75t_L g2324 ( 
.A(n_2187),
.B(n_1895),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2197),
.Y(n_2325)
);

AOI22xp33_ASAP7_75t_L g2326 ( 
.A1(n_2292),
.A2(n_2037),
.B1(n_2066),
.B2(n_2029),
.Y(n_2326)
);

NAND3xp33_ASAP7_75t_L g2327 ( 
.A(n_2292),
.B(n_2179),
.C(n_2068),
.Y(n_2327)
);

OR2x2_ASAP7_75t_L g2328 ( 
.A(n_2187),
.B(n_2205),
.Y(n_2328)
);

NOR2x1_ASAP7_75t_L g2329 ( 
.A(n_2249),
.B(n_2037),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2183),
.B(n_2179),
.Y(n_2330)
);

HB1xp67_ASAP7_75t_L g2331 ( 
.A(n_2281),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2201),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_2183),
.B(n_2030),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2208),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2190),
.Y(n_2335)
);

NOR2x1_ASAP7_75t_L g2336 ( 
.A(n_2249),
.B(n_2035),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2193),
.B(n_2158),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2194),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2194),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2211),
.Y(n_2340)
);

AND2x4_ASAP7_75t_L g2341 ( 
.A(n_2235),
.B(n_2027),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2215),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2209),
.Y(n_2343)
);

OAI211xp5_ASAP7_75t_SL g2344 ( 
.A1(n_2192),
.A2(n_2048),
.B(n_2091),
.C(n_2067),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2193),
.B(n_2158),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2198),
.B(n_2027),
.Y(n_2346)
);

AND2x4_ASAP7_75t_L g2347 ( 
.A(n_2235),
.B(n_1967),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2222),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2198),
.B(n_2144),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2199),
.B(n_2083),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2223),
.Y(n_2351)
);

HB1xp67_ASAP7_75t_L g2352 ( 
.A(n_2205),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2209),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2199),
.B(n_2040),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2250),
.Y(n_2355)
);

NAND2x1p5_ASAP7_75t_L g2356 ( 
.A(n_2255),
.B(n_1894),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2218),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2217),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2278),
.B(n_1988),
.Y(n_2359)
);

OR2x2_ASAP7_75t_L g2360 ( 
.A(n_2241),
.B(n_2028),
.Y(n_2360)
);

AOI22xp33_ASAP7_75t_L g2361 ( 
.A1(n_2292),
.A2(n_2048),
.B1(n_2004),
.B2(n_2005),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_2278),
.B(n_1910),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2217),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2219),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2219),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2207),
.Y(n_2366)
);

INVxp67_ASAP7_75t_L g2367 ( 
.A(n_2301),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2210),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2234),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2216),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2265),
.B(n_2106),
.Y(n_2371)
);

HB1xp67_ASAP7_75t_L g2372 ( 
.A(n_2284),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2216),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2273),
.B(n_1910),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_2243),
.B(n_2128),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2184),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2185),
.Y(n_2377)
);

OR2x2_ASAP7_75t_L g2378 ( 
.A(n_2241),
.B(n_1986),
.Y(n_2378)
);

HB1xp67_ASAP7_75t_L g2379 ( 
.A(n_2259),
.Y(n_2379)
);

INVx3_ASAP7_75t_L g2380 ( 
.A(n_2295),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2225),
.B(n_2152),
.Y(n_2381)
);

OR2x2_ASAP7_75t_L g2382 ( 
.A(n_2226),
.B(n_1918),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2273),
.B(n_2152),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2279),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2237),
.Y(n_2385)
);

HB1xp67_ASAP7_75t_L g2386 ( 
.A(n_2259),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2237),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2189),
.B(n_1918),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2305),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_2189),
.B(n_1918),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2229),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2279),
.Y(n_2392)
);

AND2x4_ASAP7_75t_L g2393 ( 
.A(n_2235),
.B(n_2168),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2308),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2308),
.Y(n_2395)
);

OAI22xp5_ASAP7_75t_L g2396 ( 
.A1(n_2230),
.A2(n_2057),
.B1(n_2141),
.B2(n_2128),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2230),
.B(n_2164),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2238),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2244),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2245),
.Y(n_2400)
);

BUFx3_ASAP7_75t_L g2401 ( 
.A(n_2263),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2230),
.B(n_2164),
.Y(n_2402)
);

OR2x2_ASAP7_75t_L g2403 ( 
.A(n_2221),
.B(n_1899),
.Y(n_2403)
);

AND2x4_ASAP7_75t_L g2404 ( 
.A(n_2255),
.B(n_2168),
.Y(n_2404)
);

AND2x4_ASAP7_75t_L g2405 ( 
.A(n_2255),
.B(n_1965),
.Y(n_2405)
);

AND2x4_ASAP7_75t_L g2406 ( 
.A(n_2204),
.B(n_1965),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2259),
.B(n_2169),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2259),
.B(n_2169),
.Y(n_2408)
);

NOR2xp33_ASAP7_75t_L g2409 ( 
.A(n_2300),
.B(n_2095),
.Y(n_2409)
);

HB1xp67_ASAP7_75t_L g2410 ( 
.A(n_2221),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2213),
.B(n_2055),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2276),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_2213),
.B(n_2050),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2214),
.B(n_2041),
.Y(n_2414)
);

HB1xp67_ASAP7_75t_L g2415 ( 
.A(n_2304),
.Y(n_2415)
);

NAND2x1_ASAP7_75t_SL g2416 ( 
.A(n_2268),
.B(n_2153),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2247),
.Y(n_2417)
);

OR2x2_ASAP7_75t_L g2418 ( 
.A(n_2233),
.B(n_2267),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2251),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2298),
.Y(n_2420)
);

OR2x2_ASAP7_75t_L g2421 ( 
.A(n_2267),
.B(n_1899),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2383),
.B(n_2282),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2314),
.B(n_2302),
.Y(n_2423)
);

AOI211xp5_ASAP7_75t_L g2424 ( 
.A1(n_2394),
.A2(n_2228),
.B(n_2285),
.C(n_2206),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_2310),
.B(n_2242),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2313),
.Y(n_2426)
);

OAI33xp33_ASAP7_75t_L g2427 ( 
.A1(n_2321),
.A2(n_2224),
.A3(n_2239),
.B1(n_2236),
.B2(n_2287),
.B3(n_2258),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2315),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2310),
.B(n_2242),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2311),
.B(n_2246),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2394),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2361),
.B(n_2302),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2395),
.Y(n_2433)
);

AOI22xp33_ASAP7_75t_L g2434 ( 
.A1(n_2395),
.A2(n_2260),
.B1(n_2231),
.B2(n_2290),
.Y(n_2434)
);

OR2x2_ASAP7_75t_L g2435 ( 
.A(n_2328),
.B(n_2236),
.Y(n_2435)
);

HB1xp67_ASAP7_75t_L g2436 ( 
.A(n_2372),
.Y(n_2436)
);

INVx3_ASAP7_75t_L g2437 ( 
.A(n_2401),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2356),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2356),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_2311),
.B(n_2337),
.Y(n_2440)
);

AND2x4_ASAP7_75t_L g2441 ( 
.A(n_2401),
.B(n_2227),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2356),
.Y(n_2442)
);

HB1xp67_ASAP7_75t_L g2443 ( 
.A(n_2352),
.Y(n_2443)
);

BUFx6f_ASAP7_75t_L g2444 ( 
.A(n_2407),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2320),
.Y(n_2445)
);

OAI211xp5_ASAP7_75t_L g2446 ( 
.A1(n_2336),
.A2(n_2212),
.B(n_2220),
.C(n_2227),
.Y(n_2446)
);

OAI31xp33_ASAP7_75t_L g2447 ( 
.A1(n_2418),
.A2(n_2268),
.A3(n_2297),
.B(n_2299),
.Y(n_2447)
);

OAI22xp5_ASAP7_75t_L g2448 ( 
.A1(n_2327),
.A2(n_2228),
.B1(n_2240),
.B2(n_2252),
.Y(n_2448)
);

AOI22xp33_ASAP7_75t_L g2449 ( 
.A1(n_2381),
.A2(n_2303),
.B1(n_2268),
.B2(n_2275),
.Y(n_2449)
);

AND2x2_ASAP7_75t_L g2450 ( 
.A(n_2337),
.B(n_2345),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2316),
.Y(n_2451)
);

AOI33xp33_ASAP7_75t_L g2452 ( 
.A1(n_2326),
.A2(n_2291),
.A3(n_2239),
.B1(n_2240),
.B2(n_2295),
.B3(n_2204),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2322),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2325),
.Y(n_2454)
);

INVx1_ASAP7_75t_SL g2455 ( 
.A(n_2309),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2332),
.Y(n_2456)
);

HB1xp67_ASAP7_75t_L g2457 ( 
.A(n_2331),
.Y(n_2457)
);

INVx5_ASAP7_75t_SL g2458 ( 
.A(n_2318),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2316),
.Y(n_2459)
);

NAND3xp33_ASAP7_75t_L g2460 ( 
.A(n_2367),
.B(n_2293),
.C(n_2291),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2316),
.Y(n_2461)
);

NOR3xp33_ASAP7_75t_L g2462 ( 
.A(n_2408),
.B(n_2095),
.C(n_2131),
.Y(n_2462)
);

AOI322xp5_ASAP7_75t_L g2463 ( 
.A1(n_2371),
.A2(n_2291),
.A3(n_2299),
.B1(n_2297),
.B2(n_2286),
.C1(n_2204),
.C2(n_2294),
.Y(n_2463)
);

INVx2_ASAP7_75t_SL g2464 ( 
.A(n_2329),
.Y(n_2464)
);

AOI221xp5_ASAP7_75t_L g2465 ( 
.A1(n_2420),
.A2(n_2131),
.B1(n_2294),
.B2(n_2286),
.C(n_2142),
.Y(n_2465)
);

HB1xp67_ASAP7_75t_L g2466 ( 
.A(n_2379),
.Y(n_2466)
);

INVx1_ASAP7_75t_SL g2467 ( 
.A(n_2309),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2345),
.B(n_2246),
.Y(n_2468)
);

OAI21xp33_ASAP7_75t_L g2469 ( 
.A1(n_2349),
.A2(n_2203),
.B(n_2232),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2334),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2359),
.Y(n_2471)
);

OR2x2_ASAP7_75t_L g2472 ( 
.A(n_2328),
.B(n_2258),
.Y(n_2472)
);

NAND3xp33_ASAP7_75t_SL g2473 ( 
.A(n_2375),
.B(n_2277),
.C(n_2280),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2354),
.B(n_2232),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2359),
.Y(n_2475)
);

OAI33xp33_ASAP7_75t_L g2476 ( 
.A1(n_2418),
.A2(n_2253),
.A3(n_2270),
.B1(n_2274),
.B2(n_2142),
.B3(n_2141),
.Y(n_2476)
);

NAND4xp25_ASAP7_75t_L g2477 ( 
.A(n_2355),
.B(n_2354),
.C(n_2312),
.D(n_2349),
.Y(n_2477)
);

BUFx3_ASAP7_75t_L g2478 ( 
.A(n_2312),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2364),
.Y(n_2479)
);

AND2x2_ASAP7_75t_L g2480 ( 
.A(n_2330),
.B(n_2248),
.Y(n_2480)
);

AND2x4_ASAP7_75t_L g2481 ( 
.A(n_2404),
.B(n_2280),
.Y(n_2481)
);

OAI33xp33_ASAP7_75t_L g2482 ( 
.A1(n_2389),
.A2(n_2167),
.A3(n_2256),
.B1(n_2271),
.B2(n_2261),
.B3(n_2266),
.Y(n_2482)
);

AND2x2_ASAP7_75t_L g2483 ( 
.A(n_2330),
.B(n_2248),
.Y(n_2483)
);

INVxp67_ASAP7_75t_SL g2484 ( 
.A(n_2375),
.Y(n_2484)
);

BUFx3_ASAP7_75t_L g2485 ( 
.A(n_2386),
.Y(n_2485)
);

OAI221xp5_ASAP7_75t_L g2486 ( 
.A1(n_2397),
.A2(n_2256),
.B1(n_2271),
.B2(n_2266),
.C(n_2261),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2364),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2340),
.Y(n_2488)
);

AOI221xp5_ASAP7_75t_L g2489 ( 
.A1(n_2402),
.A2(n_2365),
.B1(n_2357),
.B2(n_2409),
.C(n_2415),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2342),
.Y(n_2490)
);

OAI31xp33_ASAP7_75t_SL g2491 ( 
.A1(n_2350),
.A2(n_2318),
.A3(n_2323),
.B(n_2333),
.Y(n_2491)
);

BUFx12f_ASAP7_75t_L g2492 ( 
.A(n_2318),
.Y(n_2492)
);

AND2x4_ASAP7_75t_L g2493 ( 
.A(n_2404),
.B(n_2264),
.Y(n_2493)
);

AND3x2_ASAP7_75t_L g2494 ( 
.A(n_2409),
.B(n_2269),
.C(n_2264),
.Y(n_2494)
);

AND2x4_ASAP7_75t_L g2495 ( 
.A(n_2404),
.B(n_2262),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2350),
.B(n_2254),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2369),
.B(n_2262),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2348),
.Y(n_2498)
);

AOI22xp33_ASAP7_75t_L g2499 ( 
.A1(n_2384),
.A2(n_2392),
.B1(n_2333),
.B2(n_2335),
.Y(n_2499)
);

OAI22xp5_ASAP7_75t_L g2500 ( 
.A1(n_2360),
.A2(n_2269),
.B1(n_2257),
.B2(n_2254),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2368),
.B(n_2203),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2323),
.B(n_2413),
.Y(n_2502)
);

INVxp67_ASAP7_75t_SL g2503 ( 
.A(n_2319),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2317),
.Y(n_2504)
);

NAND3xp33_ASAP7_75t_L g2505 ( 
.A(n_2396),
.B(n_2296),
.C(n_2269),
.Y(n_2505)
);

AOI22xp5_ASAP7_75t_L g2506 ( 
.A1(n_2344),
.A2(n_2257),
.B1(n_2296),
.B2(n_2272),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_SL g2507 ( 
.A(n_2319),
.B(n_2380),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2413),
.B(n_2214),
.Y(n_2508)
);

NAND3xp33_ASAP7_75t_L g2509 ( 
.A(n_2376),
.B(n_2296),
.C(n_2289),
.Y(n_2509)
);

AND3x2_ASAP7_75t_L g2510 ( 
.A(n_2484),
.B(n_2410),
.C(n_2393),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2502),
.B(n_2366),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2440),
.B(n_2370),
.Y(n_2512)
);

AND2x2_ASAP7_75t_L g2513 ( 
.A(n_2440),
.B(n_2373),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2443),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2474),
.B(n_2346),
.Y(n_2515)
);

OR2x2_ASAP7_75t_L g2516 ( 
.A(n_2455),
.B(n_2385),
.Y(n_2516)
);

INVx1_ASAP7_75t_SL g2517 ( 
.A(n_2478),
.Y(n_2517)
);

OR2x2_ASAP7_75t_L g2518 ( 
.A(n_2467),
.B(n_2387),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2474),
.B(n_2346),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2480),
.B(n_2483),
.Y(n_2520)
);

OAI221xp5_ASAP7_75t_L g2521 ( 
.A1(n_2449),
.A2(n_2416),
.B1(n_2360),
.B2(n_2421),
.C(n_2384),
.Y(n_2521)
);

INVxp67_ASAP7_75t_SL g2522 ( 
.A(n_2478),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2480),
.B(n_2374),
.Y(n_2523)
);

OAI211xp5_ASAP7_75t_SL g2524 ( 
.A1(n_2452),
.A2(n_2380),
.B(n_2319),
.C(n_2377),
.Y(n_2524)
);

OR2x2_ASAP7_75t_L g2525 ( 
.A(n_2477),
.B(n_2351),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2483),
.B(n_2374),
.Y(n_2526)
);

AOI22xp33_ASAP7_75t_L g2527 ( 
.A1(n_2462),
.A2(n_2392),
.B1(n_2335),
.B2(n_2338),
.Y(n_2527)
);

OR2x6_ASAP7_75t_L g2528 ( 
.A(n_2464),
.B(n_2416),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2451),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2451),
.Y(n_2530)
);

NAND2xp33_ASAP7_75t_L g2531 ( 
.A(n_2464),
.B(n_2378),
.Y(n_2531)
);

OR2x2_ASAP7_75t_L g2532 ( 
.A(n_2472),
.B(n_2391),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2459),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2450),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2450),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2496),
.B(n_2362),
.Y(n_2536)
);

OR2x2_ASAP7_75t_L g2537 ( 
.A(n_2472),
.B(n_2398),
.Y(n_2537)
);

OR2x2_ASAP7_75t_L g2538 ( 
.A(n_2435),
.B(n_2399),
.Y(n_2538)
);

INVx1_ASAP7_75t_SL g2539 ( 
.A(n_2502),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2431),
.Y(n_2540)
);

INVxp67_ASAP7_75t_L g2541 ( 
.A(n_2441),
.Y(n_2541)
);

NOR3xp33_ASAP7_75t_L g2542 ( 
.A(n_2427),
.B(n_2380),
.C(n_2338),
.Y(n_2542)
);

AOI221xp5_ASAP7_75t_L g2543 ( 
.A1(n_2489),
.A2(n_2339),
.B1(n_2317),
.B2(n_2382),
.C(n_2421),
.Y(n_2543)
);

AND2x2_ASAP7_75t_L g2544 ( 
.A(n_2496),
.B(n_2362),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2437),
.B(n_2414),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2437),
.B(n_2414),
.Y(n_2546)
);

OR2x2_ASAP7_75t_L g2547 ( 
.A(n_2435),
.B(n_2400),
.Y(n_2547)
);

HB1xp67_ASAP7_75t_L g2548 ( 
.A(n_2485),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2437),
.B(n_2411),
.Y(n_2549)
);

AND2x4_ASAP7_75t_L g2550 ( 
.A(n_2441),
.B(n_2341),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2459),
.Y(n_2551)
);

INVxp67_ASAP7_75t_SL g2552 ( 
.A(n_2436),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2461),
.Y(n_2553)
);

AND2x2_ASAP7_75t_L g2554 ( 
.A(n_2493),
.B(n_2411),
.Y(n_2554)
);

OR2x2_ASAP7_75t_L g2555 ( 
.A(n_2431),
.B(n_2417),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_2461),
.Y(n_2556)
);

OAI322xp33_ASAP7_75t_L g2557 ( 
.A1(n_2448),
.A2(n_2423),
.A3(n_2433),
.B1(n_2432),
.B2(n_2422),
.C1(n_2460),
.C2(n_2505),
.Y(n_2557)
);

AND2x2_ASAP7_75t_L g2558 ( 
.A(n_2493),
.B(n_2341),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2466),
.B(n_2419),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2468),
.B(n_2378),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2458),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2493),
.B(n_2341),
.Y(n_2562)
);

NAND3xp33_ASAP7_75t_L g2563 ( 
.A(n_2465),
.B(n_2339),
.C(n_2382),
.Y(n_2563)
);

AOI21xp5_ASAP7_75t_L g2564 ( 
.A1(n_2473),
.A2(n_2393),
.B(n_2406),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2441),
.B(n_2388),
.Y(n_2565)
);

HB1xp67_ASAP7_75t_L g2566 ( 
.A(n_2485),
.Y(n_2566)
);

AOI22xp5_ASAP7_75t_L g2567 ( 
.A1(n_2476),
.A2(n_2393),
.B1(n_2347),
.B2(n_2412),
.Y(n_2567)
);

AND2x2_ASAP7_75t_L g2568 ( 
.A(n_2481),
.B(n_2495),
.Y(n_2568)
);

INVx1_ASAP7_75t_SL g2569 ( 
.A(n_2494),
.Y(n_2569)
);

OR2x2_ASAP7_75t_L g2570 ( 
.A(n_2433),
.B(n_2324),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2468),
.B(n_2388),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_SL g2572 ( 
.A(n_2452),
.B(n_2406),
.Y(n_2572)
);

AND2x2_ASAP7_75t_L g2573 ( 
.A(n_2481),
.B(n_2390),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2481),
.B(n_2390),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2495),
.B(n_2324),
.Y(n_2575)
);

INVx3_ASAP7_75t_L g2576 ( 
.A(n_2495),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2458),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2497),
.B(n_2272),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2426),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2428),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2445),
.Y(n_2581)
);

INVx1_ASAP7_75t_SL g2582 ( 
.A(n_2492),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_SL g2583 ( 
.A(n_2424),
.B(n_2406),
.Y(n_2583)
);

BUFx2_ASAP7_75t_SL g2584 ( 
.A(n_2503),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2508),
.B(n_2347),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2457),
.B(n_2412),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2458),
.Y(n_2587)
);

AND2x2_ASAP7_75t_L g2588 ( 
.A(n_2508),
.B(n_2347),
.Y(n_2588)
);

AND2x2_ASAP7_75t_L g2589 ( 
.A(n_2425),
.B(n_2405),
.Y(n_2589)
);

NAND3xp33_ASAP7_75t_L g2590 ( 
.A(n_2463),
.B(n_2353),
.C(n_2343),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2458),
.Y(n_2591)
);

AND2x2_ASAP7_75t_L g2592 ( 
.A(n_2520),
.B(n_2425),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2534),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2520),
.B(n_2429),
.Y(n_2594)
);

OR2x2_ASAP7_75t_L g2595 ( 
.A(n_2539),
.B(n_2501),
.Y(n_2595)
);

OR2x2_ASAP7_75t_L g2596 ( 
.A(n_2535),
.B(n_2453),
.Y(n_2596)
);

OAI21xp33_ASAP7_75t_L g2597 ( 
.A1(n_2524),
.A2(n_2469),
.B(n_2506),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2528),
.Y(n_2598)
);

INVx3_ASAP7_75t_L g2599 ( 
.A(n_2510),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2522),
.B(n_2454),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2529),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2545),
.B(n_2429),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2545),
.B(n_2546),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2529),
.Y(n_2604)
);

HB1xp67_ASAP7_75t_L g2605 ( 
.A(n_2548),
.Y(n_2605)
);

OR2x2_ASAP7_75t_L g2606 ( 
.A(n_2517),
.B(n_2456),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2530),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2549),
.B(n_2470),
.Y(n_2608)
);

OR2x6_ASAP7_75t_L g2609 ( 
.A(n_2528),
.B(n_2492),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2530),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2549),
.B(n_2488),
.Y(n_2611)
);

NOR2xp33_ASAP7_75t_L g2612 ( 
.A(n_2541),
.B(n_2446),
.Y(n_2612)
);

HB1xp67_ASAP7_75t_L g2613 ( 
.A(n_2566),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2546),
.B(n_2490),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2554),
.B(n_2430),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2533),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2554),
.B(n_2498),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2515),
.B(n_2430),
.Y(n_2618)
);

AND2x2_ASAP7_75t_L g2619 ( 
.A(n_2515),
.B(n_2507),
.Y(n_2619)
);

AND2x2_ASAP7_75t_L g2620 ( 
.A(n_2519),
.B(n_2507),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2568),
.B(n_2512),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_L g2622 ( 
.A(n_2582),
.B(n_2482),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2512),
.B(n_2491),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2533),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2551),
.Y(n_2625)
);

OR2x2_ASAP7_75t_L g2626 ( 
.A(n_2511),
.B(n_2471),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2528),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2513),
.B(n_2471),
.Y(n_2628)
);

HB1xp67_ASAP7_75t_L g2629 ( 
.A(n_2514),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2513),
.B(n_2475),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2568),
.B(n_2500),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2552),
.B(n_2475),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2551),
.Y(n_2633)
);

OR2x2_ASAP7_75t_L g2634 ( 
.A(n_2516),
.B(n_2499),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2576),
.B(n_2584),
.Y(n_2635)
);

AND2x4_ASAP7_75t_L g2636 ( 
.A(n_2576),
.B(n_2509),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2553),
.Y(n_2637)
);

OR2x2_ASAP7_75t_L g2638 ( 
.A(n_2516),
.B(n_2434),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2576),
.B(n_2444),
.Y(n_2639)
);

OR2x2_ASAP7_75t_L g2640 ( 
.A(n_2518),
.B(n_2438),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2519),
.B(n_2558),
.Y(n_2641)
);

INVx1_ASAP7_75t_SL g2642 ( 
.A(n_2569),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2558),
.B(n_2438),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2584),
.B(n_2444),
.Y(n_2644)
);

INVx2_ASAP7_75t_SL g2645 ( 
.A(n_2550),
.Y(n_2645)
);

NOR2xp33_ASAP7_75t_L g2646 ( 
.A(n_2557),
.B(n_2444),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2562),
.B(n_2439),
.Y(n_2647)
);

OR2x2_ASAP7_75t_L g2648 ( 
.A(n_2518),
.B(n_2439),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2553),
.Y(n_2649)
);

OR2x2_ASAP7_75t_L g2650 ( 
.A(n_2525),
.B(n_2442),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2556),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2575),
.B(n_2444),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2528),
.Y(n_2653)
);

INVxp67_ASAP7_75t_SL g2654 ( 
.A(n_2599),
.Y(n_2654)
);

HB1xp67_ASAP7_75t_L g2655 ( 
.A(n_2603),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2603),
.Y(n_2656)
);

AND2x2_ASAP7_75t_L g2657 ( 
.A(n_2592),
.B(n_2562),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2605),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2592),
.Y(n_2659)
);

INVxp67_ASAP7_75t_L g2660 ( 
.A(n_2646),
.Y(n_2660)
);

NAND2x1_ASAP7_75t_SL g2661 ( 
.A(n_2599),
.B(n_2550),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2605),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2613),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2613),
.Y(n_2664)
);

NOR2xp33_ASAP7_75t_SL g2665 ( 
.A(n_2646),
.B(n_2561),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2629),
.Y(n_2666)
);

NOR3xp33_ASAP7_75t_L g2667 ( 
.A(n_2599),
.B(n_2531),
.C(n_2542),
.Y(n_2667)
);

OAI21xp33_ASAP7_75t_L g2668 ( 
.A1(n_2597),
.A2(n_2560),
.B(n_2572),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2629),
.Y(n_2669)
);

AND2x4_ASAP7_75t_L g2670 ( 
.A(n_2645),
.B(n_2561),
.Y(n_2670)
);

OAI21xp5_ASAP7_75t_L g2671 ( 
.A1(n_2622),
.A2(n_2531),
.B(n_2590),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2594),
.B(n_2602),
.Y(n_2672)
);

AOI32xp33_ASAP7_75t_L g2673 ( 
.A1(n_2622),
.A2(n_2521),
.A3(n_2583),
.B1(n_2527),
.B2(n_2543),
.Y(n_2673)
);

AOI33xp33_ASAP7_75t_L g2674 ( 
.A1(n_2642),
.A2(n_2591),
.A3(n_2577),
.B1(n_2587),
.B2(n_2579),
.B3(n_2580),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2594),
.B(n_2550),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2602),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2628),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2630),
.Y(n_2678)
);

OAI22xp5_ASAP7_75t_L g2679 ( 
.A1(n_2623),
.A2(n_2525),
.B1(n_2586),
.B2(n_2537),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2632),
.Y(n_2680)
);

INVx2_ASAP7_75t_SL g2681 ( 
.A(n_2641),
.Y(n_2681)
);

OAI21xp5_ASAP7_75t_L g2682 ( 
.A1(n_2612),
.A2(n_2556),
.B(n_2540),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2601),
.B(n_2579),
.Y(n_2683)
);

AOI22xp5_ASAP7_75t_L g2684 ( 
.A1(n_2638),
.A2(n_2563),
.B1(n_2567),
.B2(n_2540),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2618),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2615),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2618),
.Y(n_2687)
);

OR2x6_ASAP7_75t_L g2688 ( 
.A(n_2609),
.B(n_2577),
.Y(n_2688)
);

NOR2xp33_ASAP7_75t_L g2689 ( 
.A(n_2609),
.B(n_2587),
.Y(n_2689)
);

AOI22xp5_ASAP7_75t_L g2690 ( 
.A1(n_2634),
.A2(n_2591),
.B1(n_2442),
.B2(n_2575),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2604),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2621),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2607),
.B(n_2580),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2641),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2619),
.B(n_2585),
.Y(n_2695)
);

AOI22xp5_ASAP7_75t_L g2696 ( 
.A1(n_2610),
.A2(n_2585),
.B1(n_2588),
.B2(n_2570),
.Y(n_2696)
);

NAND4xp25_ASAP7_75t_L g2697 ( 
.A(n_2612),
.B(n_2559),
.C(n_2564),
.D(n_2581),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2616),
.Y(n_2698)
);

AOI22xp5_ASAP7_75t_L g2699 ( 
.A1(n_2624),
.A2(n_2588),
.B1(n_2570),
.B2(n_2479),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2625),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2661),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2655),
.Y(n_2702)
);

O2A1O1Ixp33_ASAP7_75t_L g2703 ( 
.A1(n_2671),
.A2(n_2609),
.B(n_2644),
.C(n_2637),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2672),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2681),
.B(n_2619),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2671),
.B(n_2633),
.Y(n_2706)
);

AOI22xp33_ASAP7_75t_L g2707 ( 
.A1(n_2667),
.A2(n_2651),
.B1(n_2649),
.B2(n_2487),
.Y(n_2707)
);

AOI22xp5_ASAP7_75t_L g2708 ( 
.A1(n_2665),
.A2(n_2652),
.B1(n_2647),
.B2(n_2643),
.Y(n_2708)
);

OAI21xp33_ASAP7_75t_L g2709 ( 
.A1(n_2668),
.A2(n_2665),
.B(n_2695),
.Y(n_2709)
);

OAI32xp33_ASAP7_75t_L g2710 ( 
.A1(n_2667),
.A2(n_2650),
.A3(n_2620),
.B1(n_2639),
.B2(n_2608),
.Y(n_2710)
);

OR2x2_ASAP7_75t_L g2711 ( 
.A(n_2659),
.B(n_2611),
.Y(n_2711)
);

INVx1_ASAP7_75t_SL g2712 ( 
.A(n_2675),
.Y(n_2712)
);

INVx3_ASAP7_75t_L g2713 ( 
.A(n_2670),
.Y(n_2713)
);

AOI21xp5_ASAP7_75t_L g2714 ( 
.A1(n_2682),
.A2(n_2636),
.B(n_2635),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2694),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2656),
.Y(n_2716)
);

O2A1O1Ixp33_ASAP7_75t_SL g2717 ( 
.A1(n_2685),
.A2(n_2645),
.B(n_2617),
.C(n_2614),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2682),
.B(n_2581),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2687),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2676),
.Y(n_2720)
);

NOR3xp33_ASAP7_75t_L g2721 ( 
.A(n_2660),
.B(n_2627),
.C(n_2598),
.Y(n_2721)
);

AOI221x1_ASAP7_75t_L g2722 ( 
.A1(n_2658),
.A2(n_2653),
.B1(n_2627),
.B2(n_2598),
.C(n_2600),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2654),
.Y(n_2723)
);

A2O1A1Ixp33_ASAP7_75t_L g2724 ( 
.A1(n_2673),
.A2(n_2636),
.B(n_2447),
.C(n_2640),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2657),
.B(n_2620),
.Y(n_2725)
);

OAI22xp33_ASAP7_75t_L g2726 ( 
.A1(n_2684),
.A2(n_2648),
.B1(n_2555),
.B2(n_2653),
.Y(n_2726)
);

OAI22xp5_ASAP7_75t_L g2727 ( 
.A1(n_2660),
.A2(n_2636),
.B1(n_2595),
.B2(n_2626),
.Y(n_2727)
);

OAI22xp33_ASAP7_75t_L g2728 ( 
.A1(n_2690),
.A2(n_2555),
.B1(n_2486),
.B2(n_2547),
.Y(n_2728)
);

INVx1_ASAP7_75t_SL g2729 ( 
.A(n_2670),
.Y(n_2729)
);

O2A1O1Ixp33_ASAP7_75t_L g2730 ( 
.A1(n_2679),
.A2(n_2606),
.B(n_2593),
.C(n_2596),
.Y(n_2730)
);

NOR2xp33_ASAP7_75t_L g2731 ( 
.A(n_2688),
.B(n_2578),
.Y(n_2731)
);

O2A1O1Ixp33_ASAP7_75t_SL g2732 ( 
.A1(n_2679),
.A2(n_2537),
.B(n_2532),
.C(n_2538),
.Y(n_2732)
);

AOI22xp5_ASAP7_75t_L g2733 ( 
.A1(n_2697),
.A2(n_2643),
.B1(n_2647),
.B2(n_2631),
.Y(n_2733)
);

HB1xp67_ASAP7_75t_L g2734 ( 
.A(n_2692),
.Y(n_2734)
);

O2A1O1Ixp33_ASAP7_75t_L g2735 ( 
.A1(n_2666),
.A2(n_2538),
.B(n_2547),
.C(n_2532),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2686),
.B(n_2523),
.Y(n_2736)
);

OAI22xp33_ASAP7_75t_L g2737 ( 
.A1(n_2699),
.A2(n_2696),
.B1(n_2693),
.B2(n_2683),
.Y(n_2737)
);

AOI22xp5_ASAP7_75t_L g2738 ( 
.A1(n_2689),
.A2(n_2479),
.B1(n_2504),
.B2(n_2487),
.Y(n_2738)
);

AOI221xp5_ASAP7_75t_L g2739 ( 
.A1(n_2726),
.A2(n_2700),
.B1(n_2698),
.B2(n_2691),
.C(n_2683),
.Y(n_2739)
);

OAI21xp5_ASAP7_75t_L g2740 ( 
.A1(n_2706),
.A2(n_2669),
.B(n_2688),
.Y(n_2740)
);

HB1xp67_ASAP7_75t_L g2741 ( 
.A(n_2725),
.Y(n_2741)
);

OAI21xp33_ASAP7_75t_L g2742 ( 
.A1(n_2709),
.A2(n_2674),
.B(n_2688),
.Y(n_2742)
);

NOR2xp33_ASAP7_75t_L g2743 ( 
.A(n_2713),
.B(n_2680),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2713),
.B(n_2677),
.Y(n_2744)
);

INVxp67_ASAP7_75t_L g2745 ( 
.A(n_2701),
.Y(n_2745)
);

INVxp67_ASAP7_75t_L g2746 ( 
.A(n_2734),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2712),
.B(n_2678),
.Y(n_2747)
);

OAI221xp5_ASAP7_75t_L g2748 ( 
.A1(n_2706),
.A2(n_2693),
.B1(n_2663),
.B2(n_2664),
.C(n_2662),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2705),
.Y(n_2749)
);

NOR2xp33_ASAP7_75t_L g2750 ( 
.A(n_2729),
.B(n_2565),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2736),
.Y(n_2751)
);

NOR3xp33_ASAP7_75t_L g2752 ( 
.A(n_2727),
.B(n_2504),
.C(n_2571),
.Y(n_2752)
);

AOI322xp5_ASAP7_75t_L g2753 ( 
.A1(n_2718),
.A2(n_2523),
.A3(n_2526),
.B1(n_2544),
.B2(n_2536),
.C1(n_2565),
.C2(n_2573),
.Y(n_2753)
);

O2A1O1Ixp33_ASAP7_75t_L g2754 ( 
.A1(n_2732),
.A2(n_2103),
.B(n_2526),
.C(n_2353),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2733),
.B(n_2536),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2704),
.B(n_2544),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2711),
.Y(n_2757)
);

NOR2xp33_ASAP7_75t_L g2758 ( 
.A(n_2727),
.B(n_2708),
.Y(n_2758)
);

AOI21xp5_ASAP7_75t_L g2759 ( 
.A1(n_2718),
.A2(n_2358),
.B(n_2343),
.Y(n_2759)
);

AOI21xp33_ASAP7_75t_L g2760 ( 
.A1(n_2730),
.A2(n_2363),
.B(n_2358),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2723),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2702),
.Y(n_2762)
);

NAND3xp33_ASAP7_75t_L g2763 ( 
.A(n_2722),
.B(n_2714),
.C(n_2707),
.Y(n_2763)
);

AOI221xp5_ASAP7_75t_L g2764 ( 
.A1(n_2728),
.A2(n_2363),
.B1(n_2573),
.B2(n_2574),
.C(n_2589),
.Y(n_2764)
);

OAI21xp5_ASAP7_75t_SL g2765 ( 
.A1(n_2703),
.A2(n_2574),
.B(n_2589),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2724),
.B(n_2405),
.Y(n_2766)
);

OAI22xp33_ASAP7_75t_SL g2767 ( 
.A1(n_2738),
.A2(n_2403),
.B1(n_2405),
.B2(n_2289),
.Y(n_2767)
);

AOI22xp33_ASAP7_75t_SL g2768 ( 
.A1(n_2710),
.A2(n_2715),
.B1(n_2716),
.B2(n_2731),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2735),
.Y(n_2769)
);

OAI22xp33_ASAP7_75t_L g2770 ( 
.A1(n_2737),
.A2(n_2403),
.B1(n_2276),
.B2(n_2283),
.Y(n_2770)
);

NOR2xp33_ASAP7_75t_SL g2771 ( 
.A(n_2741),
.B(n_2719),
.Y(n_2771)
);

AOI211xp5_ASAP7_75t_SL g2772 ( 
.A1(n_2758),
.A2(n_2717),
.B(n_2720),
.C(n_2721),
.Y(n_2772)
);

INVxp67_ASAP7_75t_SL g2773 ( 
.A(n_2746),
.Y(n_2773)
);

AOI221xp5_ASAP7_75t_L g2774 ( 
.A1(n_2763),
.A2(n_2103),
.B1(n_2306),
.B2(n_2307),
.C(n_2283),
.Y(n_2774)
);

NAND3xp33_ASAP7_75t_SL g2775 ( 
.A(n_2768),
.B(n_2177),
.C(n_2096),
.Y(n_2775)
);

AOI221x1_ASAP7_75t_SL g2776 ( 
.A1(n_2742),
.A2(n_64),
.B1(n_60),
.B2(n_62),
.C(n_65),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2756),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2768),
.B(n_64),
.Y(n_2778)
);

AOI22xp33_ASAP7_75t_L g2779 ( 
.A1(n_2769),
.A2(n_2760),
.B1(n_2752),
.B2(n_2766),
.Y(n_2779)
);

NOR2xp33_ASAP7_75t_SL g2780 ( 
.A(n_2747),
.B(n_2096),
.Y(n_2780)
);

AOI221xp5_ASAP7_75t_L g2781 ( 
.A1(n_2754),
.A2(n_2307),
.B1(n_2306),
.B2(n_2127),
.C(n_2126),
.Y(n_2781)
);

OAI222xp33_ASAP7_75t_L g2782 ( 
.A1(n_2754),
.A2(n_2070),
.B1(n_2114),
.B2(n_2073),
.C1(n_2143),
.C2(n_2159),
.Y(n_2782)
);

NAND4xp75_ASAP7_75t_L g2783 ( 
.A(n_2740),
.B(n_1894),
.C(n_67),
.D(n_65),
.Y(n_2783)
);

NOR2xp67_ASAP7_75t_L g2784 ( 
.A(n_2751),
.B(n_2757),
.Y(n_2784)
);

AOI22xp33_ASAP7_75t_L g2785 ( 
.A1(n_2759),
.A2(n_1894),
.B1(n_2018),
.B2(n_1924),
.Y(n_2785)
);

AOI221xp5_ASAP7_75t_L g2786 ( 
.A1(n_2739),
.A2(n_2114),
.B1(n_2171),
.B2(n_2120),
.C(n_2116),
.Y(n_2786)
);

AOI221xp5_ASAP7_75t_L g2787 ( 
.A1(n_2748),
.A2(n_2759),
.B1(n_2770),
.B2(n_2745),
.C(n_2764),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2744),
.Y(n_2788)
);

OAI222xp33_ASAP7_75t_L g2789 ( 
.A1(n_2755),
.A2(n_2105),
.B1(n_2172),
.B2(n_2101),
.C1(n_2080),
.C2(n_2079),
.Y(n_2789)
);

AOI21xp5_ASAP7_75t_L g2790 ( 
.A1(n_2765),
.A2(n_66),
.B(n_68),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2750),
.B(n_66),
.Y(n_2791)
);

A2O1A1Ixp33_ASAP7_75t_L g2792 ( 
.A1(n_2743),
.A2(n_2761),
.B(n_2753),
.C(n_2762),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_SL g2793 ( 
.A(n_2749),
.B(n_2078),
.Y(n_2793)
);

AOI21xp5_ASAP7_75t_L g2794 ( 
.A1(n_2767),
.A2(n_68),
.B(n_69),
.Y(n_2794)
);

OAI21xp33_ASAP7_75t_SL g2795 ( 
.A1(n_2753),
.A2(n_71),
.B(n_72),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2791),
.Y(n_2796)
);

OAI31xp33_ASAP7_75t_L g2797 ( 
.A1(n_2772),
.A2(n_2778),
.A3(n_2779),
.B(n_2794),
.Y(n_2797)
);

INVxp67_ASAP7_75t_SL g2798 ( 
.A(n_2784),
.Y(n_2798)
);

AOI22xp5_ASAP7_75t_L g2799 ( 
.A1(n_2795),
.A2(n_1894),
.B1(n_1965),
.B2(n_1924),
.Y(n_2799)
);

AOI221xp5_ASAP7_75t_L g2800 ( 
.A1(n_2787),
.A2(n_1920),
.B1(n_1926),
.B2(n_75),
.C(n_76),
.Y(n_2800)
);

OAI322xp33_ASAP7_75t_SL g2801 ( 
.A1(n_2777),
.A2(n_73),
.A3(n_74),
.B1(n_75),
.B2(n_77),
.C1(n_80),
.C2(n_81),
.Y(n_2801)
);

AOI22xp5_ASAP7_75t_L g2802 ( 
.A1(n_2780),
.A2(n_1920),
.B1(n_1926),
.B2(n_1980),
.Y(n_2802)
);

A2O1A1Ixp33_ASAP7_75t_L g2803 ( 
.A1(n_2776),
.A2(n_83),
.B(n_74),
.C(n_82),
.Y(n_2803)
);

O2A1O1Ixp33_ASAP7_75t_L g2804 ( 
.A1(n_2775),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_2804)
);

NOR2xp33_ASAP7_75t_L g2805 ( 
.A(n_2771),
.B(n_85),
.Y(n_2805)
);

OR3x1_ASAP7_75t_L g2806 ( 
.A(n_2788),
.B(n_85),
.C(n_87),
.Y(n_2806)
);

NOR2xp33_ASAP7_75t_L g2807 ( 
.A(n_2773),
.B(n_88),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2792),
.Y(n_2808)
);

AOI22xp5_ASAP7_75t_L g2809 ( 
.A1(n_2775),
.A2(n_1980),
.B1(n_2008),
.B2(n_1996),
.Y(n_2809)
);

NAND4xp25_ASAP7_75t_L g2810 ( 
.A(n_2790),
.B(n_91),
.C(n_88),
.D(n_90),
.Y(n_2810)
);

OAI221xp5_ASAP7_75t_L g2811 ( 
.A1(n_2774),
.A2(n_1980),
.B1(n_94),
.B2(n_97),
.C(n_98),
.Y(n_2811)
);

AOI222xp33_ASAP7_75t_L g2812 ( 
.A1(n_2781),
.A2(n_91),
.B1(n_94),
.B2(n_98),
.C1(n_99),
.C2(n_100),
.Y(n_2812)
);

INVxp67_ASAP7_75t_L g2813 ( 
.A(n_2783),
.Y(n_2813)
);

AOI21xp5_ASAP7_75t_L g2814 ( 
.A1(n_2793),
.A2(n_100),
.B(n_101),
.Y(n_2814)
);

OAI22xp5_ASAP7_75t_L g2815 ( 
.A1(n_2798),
.A2(n_2785),
.B1(n_2786),
.B2(n_2789),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2806),
.Y(n_2816)
);

NAND3xp33_ASAP7_75t_L g2817 ( 
.A(n_2797),
.B(n_2782),
.C(n_102),
.Y(n_2817)
);

NOR2x1_ASAP7_75t_L g2818 ( 
.A(n_2808),
.B(n_104),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2796),
.Y(n_2819)
);

INVxp67_ASAP7_75t_L g2820 ( 
.A(n_2805),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2807),
.Y(n_2821)
);

XOR2xp5_ASAP7_75t_L g2822 ( 
.A(n_2810),
.B(n_105),
.Y(n_2822)
);

HB1xp67_ASAP7_75t_L g2823 ( 
.A(n_2813),
.Y(n_2823)
);

AOI221xp5_ASAP7_75t_L g2824 ( 
.A1(n_2804),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.C(n_108),
.Y(n_2824)
);

AOI211xp5_ASAP7_75t_L g2825 ( 
.A1(n_2803),
.A2(n_2800),
.B(n_2814),
.C(n_2811),
.Y(n_2825)
);

A2O1A1Ixp33_ASAP7_75t_L g2826 ( 
.A1(n_2799),
.A2(n_109),
.B(n_106),
.C(n_107),
.Y(n_2826)
);

O2A1O1Ixp33_ASAP7_75t_L g2827 ( 
.A1(n_2812),
.A2(n_112),
.B(n_110),
.C(n_111),
.Y(n_2827)
);

OAI22xp5_ASAP7_75t_L g2828 ( 
.A1(n_2819),
.A2(n_2809),
.B1(n_2802),
.B2(n_2801),
.Y(n_2828)
);

NAND4xp75_ASAP7_75t_L g2829 ( 
.A(n_2818),
.B(n_114),
.C(n_110),
.D(n_112),
.Y(n_2829)
);

AND3x2_ASAP7_75t_L g2830 ( 
.A(n_2823),
.B(n_115),
.C(n_116),
.Y(n_2830)
);

AOI221xp5_ASAP7_75t_L g2831 ( 
.A1(n_2816),
.A2(n_2815),
.B1(n_2825),
.B2(n_2827),
.C(n_2820),
.Y(n_2831)
);

AO22x2_ASAP7_75t_L g2832 ( 
.A1(n_2822),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_2832)
);

OAI21xp5_ASAP7_75t_SL g2833 ( 
.A1(n_2817),
.A2(n_120),
.B(n_123),
.Y(n_2833)
);

OAI221xp5_ASAP7_75t_L g2834 ( 
.A1(n_2824),
.A2(n_120),
.B1(n_123),
.B2(n_126),
.C(n_127),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2821),
.Y(n_2835)
);

BUFx6f_ASAP7_75t_L g2836 ( 
.A(n_2826),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2818),
.Y(n_2837)
);

A2O1A1Ixp33_ASAP7_75t_L g2838 ( 
.A1(n_2816),
.A2(n_126),
.B(n_128),
.C(n_129),
.Y(n_2838)
);

INVx8_ASAP7_75t_L g2839 ( 
.A(n_2823),
.Y(n_2839)
);

OAI22xp5_ASAP7_75t_L g2840 ( 
.A1(n_2819),
.A2(n_1980),
.B1(n_1996),
.B2(n_1240),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2839),
.Y(n_2841)
);

NOR2xp33_ASAP7_75t_L g2842 ( 
.A(n_2837),
.B(n_130),
.Y(n_2842)
);

OR2x2_ASAP7_75t_L g2843 ( 
.A(n_2838),
.B(n_130),
.Y(n_2843)
);

NAND2x1_ASAP7_75t_L g2844 ( 
.A(n_2835),
.B(n_131),
.Y(n_2844)
);

AND2x4_ASAP7_75t_L g2845 ( 
.A(n_2830),
.B(n_134),
.Y(n_2845)
);

NOR2x1_ASAP7_75t_L g2846 ( 
.A(n_2829),
.B(n_135),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_2832),
.B(n_135),
.Y(n_2847)
);

O2A1O1Ixp33_ASAP7_75t_L g2848 ( 
.A1(n_2833),
.A2(n_136),
.B(n_137),
.C(n_140),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2836),
.Y(n_2849)
);

OAI22xp33_ASAP7_75t_SL g2850 ( 
.A1(n_2828),
.A2(n_2834),
.B1(n_2831),
.B2(n_2840),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2839),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2839),
.Y(n_2852)
);

INVxp67_ASAP7_75t_L g2853 ( 
.A(n_2829),
.Y(n_2853)
);

NOR2x1_ASAP7_75t_L g2854 ( 
.A(n_2838),
.B(n_136),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2839),
.Y(n_2855)
);

INVxp33_ASAP7_75t_SL g2856 ( 
.A(n_2831),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2839),
.Y(n_2857)
);

INVx3_ASAP7_75t_L g2858 ( 
.A(n_2844),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2845),
.Y(n_2859)
);

NOR2x1_ASAP7_75t_L g2860 ( 
.A(n_2841),
.B(n_137),
.Y(n_2860)
);

NOR2xp33_ASAP7_75t_L g2861 ( 
.A(n_2845),
.B(n_140),
.Y(n_2861)
);

AOI22xp33_ASAP7_75t_SL g2862 ( 
.A1(n_2856),
.A2(n_1144),
.B1(n_1165),
.B2(n_1251),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2847),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2846),
.Y(n_2864)
);

NOR2x1_ASAP7_75t_L g2865 ( 
.A(n_2851),
.B(n_141),
.Y(n_2865)
);

INVxp67_ASAP7_75t_SL g2866 ( 
.A(n_2842),
.Y(n_2866)
);

AND2x2_ASAP7_75t_L g2867 ( 
.A(n_2852),
.B(n_141),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2855),
.Y(n_2868)
);

NOR3xp33_ASAP7_75t_L g2869 ( 
.A(n_2857),
.B(n_2850),
.C(n_2849),
.Y(n_2869)
);

NAND4xp75_ASAP7_75t_L g2870 ( 
.A(n_2854),
.B(n_142),
.C(n_144),
.D(n_145),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2843),
.Y(n_2871)
);

NAND4xp75_ASAP7_75t_L g2872 ( 
.A(n_2853),
.B(n_144),
.C(n_146),
.D(n_147),
.Y(n_2872)
);

INVx1_ASAP7_75t_SL g2873 ( 
.A(n_2867),
.Y(n_2873)
);

AOI22xp5_ASAP7_75t_L g2874 ( 
.A1(n_2863),
.A2(n_2858),
.B1(n_2866),
.B2(n_2861),
.Y(n_2874)
);

OAI211xp5_ASAP7_75t_SL g2875 ( 
.A1(n_2869),
.A2(n_2848),
.B(n_148),
.C(n_149),
.Y(n_2875)
);

AOI211xp5_ASAP7_75t_L g2876 ( 
.A1(n_2868),
.A2(n_2864),
.B(n_2859),
.C(n_2858),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2860),
.B(n_147),
.Y(n_2877)
);

AOI21xp5_ASAP7_75t_L g2878 ( 
.A1(n_2865),
.A2(n_149),
.B(n_150),
.Y(n_2878)
);

OAI211xp5_ASAP7_75t_SL g2879 ( 
.A1(n_2871),
.A2(n_151),
.B(n_152),
.C(n_153),
.Y(n_2879)
);

OAI221xp5_ASAP7_75t_SL g2880 ( 
.A1(n_2862),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.C(n_157),
.Y(n_2880)
);

AOI221xp5_ASAP7_75t_L g2881 ( 
.A1(n_2870),
.A2(n_155),
.B1(n_156),
.B2(n_158),
.C(n_159),
.Y(n_2881)
);

AO22x2_ASAP7_75t_L g2882 ( 
.A1(n_2872),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_2882)
);

AOI322xp5_ASAP7_75t_L g2883 ( 
.A1(n_2863),
.A2(n_164),
.A3(n_165),
.B1(n_166),
.B2(n_167),
.C1(n_168),
.C2(n_169),
.Y(n_2883)
);

BUFx2_ASAP7_75t_L g2884 ( 
.A(n_2860),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2884),
.B(n_166),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2882),
.Y(n_2886)
);

NOR2xp33_ASAP7_75t_L g2887 ( 
.A(n_2873),
.B(n_167),
.Y(n_2887)
);

NOR2xp67_ASAP7_75t_L g2888 ( 
.A(n_2878),
.B(n_169),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2876),
.B(n_170),
.Y(n_2889)
);

INVx4_ASAP7_75t_L g2890 ( 
.A(n_2882),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2877),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2874),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2879),
.Y(n_2893)
);

NAND4xp75_ASAP7_75t_L g2894 ( 
.A(n_2881),
.B(n_170),
.C(n_171),
.D(n_173),
.Y(n_2894)
);

XNOR2xp5_ASAP7_75t_L g2895 ( 
.A(n_2875),
.B(n_171),
.Y(n_2895)
);

NAND3x1_ASAP7_75t_L g2896 ( 
.A(n_2885),
.B(n_2880),
.C(n_2883),
.Y(n_2896)
);

NOR2x1_ASAP7_75t_L g2897 ( 
.A(n_2890),
.B(n_173),
.Y(n_2897)
);

INVx2_ASAP7_75t_SL g2898 ( 
.A(n_2892),
.Y(n_2898)
);

XNOR2x1_ASAP7_75t_L g2899 ( 
.A(n_2895),
.B(n_175),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2886),
.Y(n_2900)
);

NOR2x1_ASAP7_75t_L g2901 ( 
.A(n_2889),
.B(n_176),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2891),
.Y(n_2902)
);

OAI21xp5_ASAP7_75t_L g2903 ( 
.A1(n_2888),
.A2(n_1144),
.B(n_1165),
.Y(n_2903)
);

AO22x2_ASAP7_75t_L g2904 ( 
.A1(n_2894),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_SL g2905 ( 
.A(n_2893),
.B(n_177),
.Y(n_2905)
);

AND2x4_ASAP7_75t_L g2906 ( 
.A(n_2887),
.B(n_179),
.Y(n_2906)
);

XNOR2xp5_ASAP7_75t_L g2907 ( 
.A(n_2895),
.B(n_180),
.Y(n_2907)
);

XNOR2xp5_ASAP7_75t_L g2908 ( 
.A(n_2895),
.B(n_181),
.Y(n_2908)
);

OR2x2_ASAP7_75t_L g2909 ( 
.A(n_2898),
.B(n_182),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2897),
.B(n_182),
.Y(n_2910)
);

BUFx2_ASAP7_75t_L g2911 ( 
.A(n_2901),
.Y(n_2911)
);

OAI21x1_ASAP7_75t_L g2912 ( 
.A1(n_2896),
.A2(n_183),
.B(n_185),
.Y(n_2912)
);

INVxp67_ASAP7_75t_SL g2913 ( 
.A(n_2902),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2904),
.Y(n_2914)
);

AOI21x1_ASAP7_75t_L g2915 ( 
.A1(n_2900),
.A2(n_185),
.B(n_187),
.Y(n_2915)
);

INVx3_ASAP7_75t_L g2916 ( 
.A(n_2906),
.Y(n_2916)
);

INVx2_ASAP7_75t_SL g2917 ( 
.A(n_2899),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2911),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2915),
.Y(n_2919)
);

AOI22xp5_ASAP7_75t_L g2920 ( 
.A1(n_2913),
.A2(n_2908),
.B1(n_2907),
.B2(n_2905),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2910),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2916),
.Y(n_2922)
);

INVx2_ASAP7_75t_SL g2923 ( 
.A(n_2909),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2912),
.Y(n_2924)
);

OAI221xp5_ASAP7_75t_L g2925 ( 
.A1(n_2917),
.A2(n_2903),
.B1(n_188),
.B2(n_189),
.C(n_190),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2914),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2911),
.Y(n_2927)
);

AOI22xp5_ASAP7_75t_L g2928 ( 
.A1(n_2913),
.A2(n_1144),
.B1(n_1165),
.B2(n_1251),
.Y(n_2928)
);

NAND2x1p5_ASAP7_75t_L g2929 ( 
.A(n_2912),
.B(n_831),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2911),
.Y(n_2930)
);

XNOR2xp5_ASAP7_75t_L g2931 ( 
.A(n_2917),
.B(n_187),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2911),
.Y(n_2932)
);

AOI22x1_ASAP7_75t_L g2933 ( 
.A1(n_2913),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2911),
.Y(n_2934)
);

OA22x2_ASAP7_75t_L g2935 ( 
.A1(n_2913),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_2935)
);

NAND3xp33_ASAP7_75t_L g2936 ( 
.A(n_2911),
.B(n_831),
.C(n_817),
.Y(n_2936)
);

XOR2xp5_ASAP7_75t_L g2937 ( 
.A(n_2917),
.B(n_193),
.Y(n_2937)
);

AO22x2_ASAP7_75t_L g2938 ( 
.A1(n_2919),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2918),
.Y(n_2939)
);

AO22x2_ASAP7_75t_L g2940 ( 
.A1(n_2924),
.A2(n_2932),
.B1(n_2930),
.B2(n_2927),
.Y(n_2940)
);

OAI22xp5_ASAP7_75t_L g2941 ( 
.A1(n_2934),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_2941)
);

AOI22x1_ASAP7_75t_L g2942 ( 
.A1(n_2926),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2929),
.Y(n_2943)
);

NOR2x1_ASAP7_75t_L g2944 ( 
.A(n_2922),
.B(n_204),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2923),
.B(n_204),
.Y(n_2945)
);

AO22x2_ASAP7_75t_L g2946 ( 
.A1(n_2937),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_2946)
);

OAI21xp5_ASAP7_75t_L g2947 ( 
.A1(n_2920),
.A2(n_1165),
.B(n_1144),
.Y(n_2947)
);

NAND4xp75_ASAP7_75t_L g2948 ( 
.A(n_2921),
.B(n_208),
.C(n_209),
.D(n_210),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2931),
.B(n_210),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2935),
.Y(n_2950)
);

OAI22x1_ASAP7_75t_L g2951 ( 
.A1(n_2933),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_2951)
);

AOI21x1_ASAP7_75t_L g2952 ( 
.A1(n_2936),
.A2(n_214),
.B(n_216),
.Y(n_2952)
);

OAI22x1_ASAP7_75t_L g2953 ( 
.A1(n_2925),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_2953)
);

OAI22xp5_ASAP7_75t_L g2954 ( 
.A1(n_2928),
.A2(n_219),
.B1(n_1154),
.B2(n_1264),
.Y(n_2954)
);

CKINVDCx20_ASAP7_75t_R g2955 ( 
.A(n_2920),
.Y(n_2955)
);

HB1xp67_ASAP7_75t_L g2956 ( 
.A(n_2918),
.Y(n_2956)
);

OAI22xp5_ASAP7_75t_L g2957 ( 
.A1(n_2918),
.A2(n_1195),
.B1(n_1264),
.B2(n_1257),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2918),
.Y(n_2958)
);

INVx2_ASAP7_75t_L g2959 ( 
.A(n_2929),
.Y(n_2959)
);

CKINVDCx20_ASAP7_75t_R g2960 ( 
.A(n_2920),
.Y(n_2960)
);

AOI22xp33_ASAP7_75t_L g2961 ( 
.A1(n_2956),
.A2(n_813),
.B1(n_817),
.B2(n_1165),
.Y(n_2961)
);

OAI21xp5_ASAP7_75t_L g2962 ( 
.A1(n_2939),
.A2(n_1264),
.B(n_1257),
.Y(n_2962)
);

AOI221xp5_ASAP7_75t_L g2963 ( 
.A1(n_2940),
.A2(n_813),
.B1(n_817),
.B2(n_1240),
.C(n_1257),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2940),
.Y(n_2964)
);

AOI21xp5_ASAP7_75t_L g2965 ( 
.A1(n_2958),
.A2(n_2949),
.B(n_2943),
.Y(n_2965)
);

OAI21xp5_ASAP7_75t_L g2966 ( 
.A1(n_2955),
.A2(n_1250),
.B(n_1240),
.Y(n_2966)
);

OAI21x1_ASAP7_75t_L g2967 ( 
.A1(n_2944),
.A2(n_1979),
.B(n_1941),
.Y(n_2967)
);

OAI21x1_ASAP7_75t_L g2968 ( 
.A1(n_2950),
.A2(n_1979),
.B(n_1941),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2946),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2960),
.B(n_221),
.Y(n_2970)
);

NOR2xp33_ASAP7_75t_R g2971 ( 
.A(n_2945),
.B(n_223),
.Y(n_2971)
);

NOR2xp33_ASAP7_75t_L g2972 ( 
.A(n_2959),
.B(n_224),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2938),
.Y(n_2973)
);

AOI22xp5_ASAP7_75t_L g2974 ( 
.A1(n_2948),
.A2(n_1250),
.B1(n_1251),
.B2(n_1185),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2938),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2951),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2942),
.Y(n_2977)
);

OAI22xp5_ASAP7_75t_SL g2978 ( 
.A1(n_2953),
.A2(n_226),
.B1(n_230),
.B2(n_236),
.Y(n_2978)
);

OAI21x1_ASAP7_75t_SL g2979 ( 
.A1(n_2952),
.A2(n_1250),
.B(n_240),
.Y(n_2979)
);

OAI22x1_ASAP7_75t_L g2980 ( 
.A1(n_2941),
.A2(n_238),
.B1(n_241),
.B2(n_243),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2964),
.B(n_2954),
.Y(n_2981)
);

AOI21xp33_ASAP7_75t_L g2982 ( 
.A1(n_2973),
.A2(n_2957),
.B(n_2947),
.Y(n_2982)
);

AOI221xp5_ASAP7_75t_L g2983 ( 
.A1(n_2969),
.A2(n_817),
.B1(n_813),
.B2(n_819),
.C(n_836),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2975),
.B(n_246),
.Y(n_2984)
);

AOI21xp5_ASAP7_75t_L g2985 ( 
.A1(n_2965),
.A2(n_817),
.B(n_813),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2976),
.B(n_247),
.Y(n_2986)
);

OAI21xp5_ASAP7_75t_L g2987 ( 
.A1(n_2977),
.A2(n_836),
.B(n_823),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2979),
.Y(n_2988)
);

AOI31xp33_ASAP7_75t_L g2989 ( 
.A1(n_2970),
.A2(n_249),
.A3(n_258),
.B(n_261),
.Y(n_2989)
);

AO221x2_ASAP7_75t_L g2990 ( 
.A1(n_2978),
.A2(n_262),
.B1(n_265),
.B2(n_267),
.C(n_268),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2971),
.Y(n_2991)
);

AOI22xp5_ASAP7_75t_L g2992 ( 
.A1(n_2988),
.A2(n_2966),
.B1(n_2972),
.B2(n_2980),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2991),
.Y(n_2993)
);

OR2x2_ASAP7_75t_L g2994 ( 
.A(n_2981),
.B(n_2962),
.Y(n_2994)
);

OAI22x1_ASAP7_75t_L g2995 ( 
.A1(n_2984),
.A2(n_2974),
.B1(n_2963),
.B2(n_2961),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2986),
.Y(n_2996)
);

AOI22xp5_ASAP7_75t_L g2997 ( 
.A1(n_2990),
.A2(n_2967),
.B1(n_2968),
.B2(n_813),
.Y(n_2997)
);

OAI22xp5_ASAP7_75t_SL g2998 ( 
.A1(n_2987),
.A2(n_270),
.B1(n_271),
.B2(n_274),
.Y(n_2998)
);

OAI22xp5_ASAP7_75t_SL g2999 ( 
.A1(n_2982),
.A2(n_279),
.B1(n_280),
.B2(n_282),
.Y(n_2999)
);

AOI22xp33_ASAP7_75t_L g3000 ( 
.A1(n_2996),
.A2(n_2985),
.B1(n_2983),
.B2(n_2989),
.Y(n_3000)
);

AOI22xp5_ASAP7_75t_L g3001 ( 
.A1(n_2993),
.A2(n_1251),
.B1(n_1129),
.B2(n_1111),
.Y(n_3001)
);

AOI22xp33_ASAP7_75t_SL g3002 ( 
.A1(n_2994),
.A2(n_836),
.B1(n_823),
.B2(n_819),
.Y(n_3002)
);

AOI22xp5_ASAP7_75t_SL g3003 ( 
.A1(n_2995),
.A2(n_283),
.B1(n_285),
.B2(n_286),
.Y(n_3003)
);

AOI22xp5_ASAP7_75t_L g3004 ( 
.A1(n_2992),
.A2(n_2998),
.B1(n_2997),
.B2(n_2999),
.Y(n_3004)
);

AOI22xp5_ASAP7_75t_L g3005 ( 
.A1(n_2993),
.A2(n_1129),
.B1(n_1111),
.B2(n_836),
.Y(n_3005)
);

AOI22xp33_ASAP7_75t_SL g3006 ( 
.A1(n_2993),
.A2(n_836),
.B1(n_823),
.B2(n_819),
.Y(n_3006)
);

INVx4_ASAP7_75t_L g3007 ( 
.A(n_3004),
.Y(n_3007)
);

HAxp5_ASAP7_75t_L g3008 ( 
.A(n_3000),
.B(n_3006),
.CON(n_3008),
.SN(n_3008)
);

AOI221xp5_ASAP7_75t_L g3009 ( 
.A1(n_3007),
.A2(n_3002),
.B1(n_3005),
.B2(n_3003),
.C(n_3001),
.Y(n_3009)
);

AOI211xp5_ASAP7_75t_L g3010 ( 
.A1(n_3009),
.A2(n_3008),
.B(n_289),
.C(n_290),
.Y(n_3010)
);


endmodule