module fake_netlist_5_1638_n_2427 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_46, n_233, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_239, n_175, n_169, n_59, n_26, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2427);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_239;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2427;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_544;
wire n_1007;
wire n_2369;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2249;
wire n_2180;
wire n_344;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_475;
wire n_1070;
wire n_777;
wire n_422;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1561;
wire n_1267;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1587;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_283;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_407;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_561;
wire n_1319;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_604;
wire n_433;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_2359;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_2346;
wire n_662;
wire n_459;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2399;
wire n_473;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2418;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_2400;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1205;
wire n_1044;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_2266;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_2333;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_378;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_302;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_321;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_2269;
wire n_2309;
wire n_2415;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_323;
wire n_2287;
wire n_356;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1928;
wire n_1848;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_2282;
wire n_510;
wire n_2371;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_2068;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_2363;
wire n_916;
wire n_1081;
wire n_493;
wire n_2332;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_377;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_994;
wire n_386;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_328;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_2278;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_2414;
wire n_246;
wire n_1583;
wire n_2426;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_2273;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;
wire n_2268;

INVx1_ASAP7_75t_L g242 ( 
.A(n_167),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_114),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_46),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_162),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_32),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_121),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_72),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_129),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_141),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_170),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_40),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_8),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_214),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_43),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_192),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_51),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_40),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_110),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_238),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_173),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_160),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_176),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_199),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_210),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_37),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_109),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_201),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_156),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_89),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_64),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_12),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_219),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_64),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_180),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_140),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_28),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_23),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_15),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_187),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_206),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_32),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_9),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_106),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_13),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_97),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_22),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_110),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_15),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_36),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_107),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_108),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_92),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_14),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_175),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_137),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_208),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_158),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_190),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_34),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_16),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_57),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_89),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_193),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_23),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_43),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_150),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_41),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_38),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_54),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_86),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_132),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_13),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_234),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_183),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_107),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_131),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_226),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_79),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_144),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_111),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_19),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_62),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_11),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_17),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_36),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_101),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_149),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_188),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_31),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_2),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_28),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_179),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_233),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_204),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_211),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_92),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_2),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_97),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_55),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_71),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_26),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_227),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_58),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_147),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_181),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_215),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_236),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_171),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_65),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_19),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_139),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_37),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_21),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_60),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_99),
.Y(n_358)
);

BUFx10_ASAP7_75t_L g359 ( 
.A(n_151),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_128),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_59),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_189),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_133),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_237),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_63),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_26),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_69),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_80),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_148),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_230),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_159),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_116),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_146),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_202),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_228),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_4),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_207),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_22),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_41),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_163),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_225),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_10),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_21),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_168),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_136),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_82),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_8),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_126),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_205),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_224),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_38),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_184),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_124),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_9),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_195),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_33),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_155),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_66),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_4),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_29),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_145),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_241),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_80),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_138),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_77),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_45),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_24),
.Y(n_407)
);

BUFx10_ASAP7_75t_L g408 ( 
.A(n_53),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_105),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_68),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_20),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_0),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_50),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_142),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_42),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_70),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_82),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_99),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_161),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_78),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_5),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_70),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_48),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_212),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_174),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_177),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_50),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_90),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_118),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_98),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_74),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_196),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_108),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_56),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_83),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_0),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_29),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_55),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_39),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_83),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_75),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_44),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_185),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_116),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_112),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_231),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_209),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_198),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_10),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_86),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_203),
.Y(n_451)
);

BUFx5_ASAP7_75t_L g452 ( 
.A(n_79),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_48),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_61),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_69),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_25),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_200),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_31),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_104),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_54),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_33),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_106),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_61),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_66),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_77),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_221),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_117),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_57),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_59),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_56),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_112),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_67),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_71),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_328),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_452),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_245),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_452),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_264),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_328),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_336),
.Y(n_480)
);

INVxp33_ASAP7_75t_L g481 ( 
.A(n_312),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_287),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_247),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_452),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_251),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_242),
.B(n_1),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_252),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_255),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_261),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_452),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_393),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_452),
.B(n_1),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_452),
.Y(n_493)
);

INVxp33_ASAP7_75t_L g494 ( 
.A(n_287),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_328),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_452),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_387),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_452),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_242),
.B(n_3),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_301),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_452),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_301),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g503 ( 
.A(n_383),
.B(n_3),
.Y(n_503)
);

CKINVDCx14_ASAP7_75t_R g504 ( 
.A(n_288),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_288),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_262),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_246),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_383),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_387),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_248),
.B(n_5),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_263),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_265),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_246),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_347),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_257),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_347),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_246),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_389),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_266),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_274),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_389),
.Y(n_521)
);

INVxp33_ASAP7_75t_SL g522 ( 
.A(n_243),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_387),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_321),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_447),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_276),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_368),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_368),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_257),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_453),
.B(n_321),
.Y(n_530)
);

INVxp33_ASAP7_75t_L g531 ( 
.A(n_279),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_277),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_282),
.Y(n_533)
);

CKINVDCx16_ASAP7_75t_R g534 ( 
.A(n_447),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_246),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_453),
.B(n_6),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_246),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_246),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_297),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_281),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_453),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_458),
.B(n_6),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_300),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_248),
.B(n_7),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_458),
.B(n_7),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_408),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_306),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_316),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_317),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_281),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_319),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_279),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_320),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_250),
.B(n_11),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_428),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_281),
.B(n_12),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_322),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_330),
.Y(n_558)
);

INVxp67_ASAP7_75t_SL g559 ( 
.A(n_428),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_254),
.B(n_14),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_284),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_331),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_281),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_281),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_281),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_335),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_348),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_284),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_250),
.B(n_16),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_291),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_350),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_351),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_360),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_291),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_364),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_244),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_269),
.B(n_17),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_369),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_370),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_291),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_291),
.Y(n_581)
);

INVxp33_ASAP7_75t_SL g582 ( 
.A(n_249),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_371),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_373),
.Y(n_584)
);

INVxp67_ASAP7_75t_SL g585 ( 
.A(n_285),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_291),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_291),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_375),
.Y(n_588)
);

INVxp67_ASAP7_75t_SL g589 ( 
.A(n_285),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_341),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_377),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_341),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_269),
.B(n_18),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g594 ( 
.A(n_296),
.Y(n_594)
);

INVxp67_ASAP7_75t_SL g595 ( 
.A(n_296),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_257),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_341),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_341),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_341),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_304),
.Y(n_600)
);

INVxp67_ASAP7_75t_SL g601 ( 
.A(n_304),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_305),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_341),
.Y(n_603)
);

INVxp67_ASAP7_75t_SL g604 ( 
.A(n_305),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_522),
.B(n_298),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_475),
.A2(n_278),
.B(n_270),
.Y(n_606)
);

OAI21x1_ASAP7_75t_L g607 ( 
.A1(n_475),
.A2(n_278),
.B(n_270),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_507),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_527),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_507),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_476),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_513),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_513),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_483),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_485),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_582),
.B(n_298),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_477),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_R g618 ( 
.A(n_549),
.B(n_380),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_487),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_488),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_477),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_489),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_517),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_500),
.B(n_259),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_506),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_511),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_478),
.B(n_353),
.Y(n_627)
);

CKINVDCx16_ASAP7_75t_R g628 ( 
.A(n_528),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_512),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_519),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_517),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_560),
.B(n_264),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_535),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_576),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_504),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_535),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_482),
.A2(n_290),
.B1(n_293),
.B2(n_275),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_478),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_537),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_520),
.Y(n_640)
);

OA21x2_ASAP7_75t_L g641 ( 
.A1(n_492),
.A2(n_299),
.B(n_283),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_534),
.B(n_546),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_526),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_537),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_532),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_R g646 ( 
.A(n_553),
.B(n_381),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_533),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_560),
.B(n_264),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_538),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_484),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_480),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_478),
.B(n_353),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_474),
.B(n_353),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_482),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_508),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_474),
.B(n_353),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_539),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_479),
.B(n_353),
.Y(n_658)
);

AND3x1_ASAP7_75t_L g659 ( 
.A(n_486),
.B(n_310),
.C(n_308),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_538),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_R g661 ( 
.A(n_562),
.B(n_566),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_540),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_479),
.B(n_353),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_540),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_495),
.B(n_372),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_543),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_550),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_547),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_550),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_505),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_563),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_484),
.Y(n_672)
);

NOR2xp67_ASAP7_75t_L g673 ( 
.A(n_490),
.B(n_283),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_534),
.B(n_359),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_563),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_559),
.B(n_372),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_495),
.B(n_349),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_505),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_564),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_564),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_548),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_565),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_565),
.Y(n_683)
);

OA21x2_ASAP7_75t_L g684 ( 
.A1(n_492),
.A2(n_309),
.B(n_299),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_570),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_490),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_551),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_570),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_493),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_574),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_491),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_530),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_557),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_574),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_567),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_558),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_580),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_573),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_580),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_575),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_578),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_579),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_581),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_621),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_654),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_R g706 ( 
.A(n_695),
.B(n_583),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_692),
.B(n_591),
.Y(n_707)
);

AO22x2_ASAP7_75t_L g708 ( 
.A1(n_674),
.A2(n_559),
.B1(n_441),
.B2(n_416),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_605),
.B(n_571),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_617),
.Y(n_710)
);

BUFx8_ASAP7_75t_SL g711 ( 
.A(n_651),
.Y(n_711)
);

NOR2x1p5_ASAP7_75t_L g712 ( 
.A(n_611),
.B(n_542),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_605),
.B(n_546),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_638),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_692),
.B(n_497),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_639),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_692),
.B(n_581),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_661),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_621),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_616),
.B(n_572),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_639),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_639),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_680),
.Y(n_723)
);

AND2x6_ASAP7_75t_L g724 ( 
.A(n_632),
.B(n_388),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_680),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_617),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_617),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_616),
.B(n_528),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_680),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_634),
.B(n_584),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_621),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_638),
.B(n_677),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_621),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_649),
.Y(n_734)
);

OR2x2_ASAP7_75t_L g735 ( 
.A(n_654),
.B(n_494),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_635),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_638),
.B(n_349),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_634),
.A2(n_588),
.B1(n_502),
.B2(n_516),
.Y(n_738)
);

OAI21xp33_ASAP7_75t_L g739 ( 
.A1(n_676),
.A2(n_531),
.B(n_510),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_677),
.Y(n_740)
);

AO22x2_ASAP7_75t_L g741 ( 
.A1(n_659),
.A2(n_441),
.B1(n_416),
.B2(n_542),
.Y(n_741)
);

AND3x4_ASAP7_75t_L g742 ( 
.A(n_628),
.B(n_503),
.C(n_260),
.Y(n_742)
);

AND2x4_ASAP7_75t_SL g743 ( 
.A(n_691),
.B(n_514),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_670),
.B(n_481),
.Y(n_744)
);

INVxp67_ASAP7_75t_SL g745 ( 
.A(n_653),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_635),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_689),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_676),
.B(n_497),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_617),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_628),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_677),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_677),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_649),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_648),
.B(n_349),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_689),
.Y(n_755)
);

INVx5_ASAP7_75t_L g756 ( 
.A(n_617),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_689),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_614),
.B(n_518),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_649),
.Y(n_759)
);

NAND2x1p5_ASAP7_75t_L g760 ( 
.A(n_641),
.B(n_374),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_648),
.B(n_586),
.Y(n_761)
);

OAI21xp33_ASAP7_75t_L g762 ( 
.A1(n_655),
.A2(n_544),
.B(n_499),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_632),
.B(n_509),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_641),
.A2(n_569),
.B1(n_577),
.B2(n_554),
.Y(n_764)
);

AO21x2_ASAP7_75t_L g765 ( 
.A1(n_606),
.A2(n_556),
.B(n_314),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_689),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_641),
.A2(n_593),
.B1(n_536),
.B2(n_556),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_648),
.B(n_374),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_615),
.B(n_521),
.Y(n_769)
);

NAND3xp33_ASAP7_75t_L g770 ( 
.A(n_659),
.B(n_555),
.C(n_508),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_627),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_632),
.B(n_509),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_627),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_652),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_652),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_609),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_608),
.Y(n_777)
);

INVx4_ASAP7_75t_SL g778 ( 
.A(n_617),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_619),
.B(n_525),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_617),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_620),
.B(n_545),
.Y(n_781)
);

BUFx8_ASAP7_75t_SL g782 ( 
.A(n_622),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_625),
.B(n_545),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_662),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_670),
.B(n_555),
.Y(n_785)
);

AO22x2_ASAP7_75t_L g786 ( 
.A1(n_655),
.A2(n_310),
.B1(n_329),
.B2(n_308),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_608),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_626),
.A2(n_503),
.B1(n_589),
.B2(n_585),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_650),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_610),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_610),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_612),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_612),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_629),
.B(n_585),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_648),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_630),
.B(n_589),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_640),
.B(n_359),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_662),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_662),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_613),
.Y(n_800)
);

INVx4_ASAP7_75t_L g801 ( 
.A(n_650),
.Y(n_801)
);

NOR2x1p5_ASAP7_75t_L g802 ( 
.A(n_643),
.B(n_594),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_613),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_L g804 ( 
.A(n_650),
.B(n_388),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_623),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_650),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_623),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_631),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_631),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_633),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_633),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_636),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_636),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_664),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_653),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_609),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_644),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_656),
.B(n_586),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_R g819 ( 
.A(n_645),
.B(n_647),
.Y(n_819)
);

AND2x6_ASAP7_75t_L g820 ( 
.A(n_650),
.B(n_388),
.Y(n_820)
);

BUFx10_ASAP7_75t_L g821 ( 
.A(n_657),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_664),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_650),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_644),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_656),
.B(n_587),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_664),
.Y(n_826)
);

INVx4_ASAP7_75t_L g827 ( 
.A(n_650),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_660),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_660),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_669),
.Y(n_830)
);

BUFx8_ASAP7_75t_SL g831 ( 
.A(n_666),
.Y(n_831)
);

OR2x6_ASAP7_75t_L g832 ( 
.A(n_642),
.B(n_536),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_658),
.B(n_587),
.Y(n_833)
);

BUFx10_ASAP7_75t_L g834 ( 
.A(n_668),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_667),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_681),
.B(n_359),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_658),
.B(n_590),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_667),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_687),
.B(n_359),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_669),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_663),
.B(n_523),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_693),
.B(n_594),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_696),
.B(n_698),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_663),
.B(n_523),
.Y(n_844)
);

INVxp33_ASAP7_75t_L g845 ( 
.A(n_678),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_669),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_665),
.B(n_541),
.Y(n_847)
);

NOR3xp33_ASAP7_75t_L g848 ( 
.A(n_678),
.B(n_530),
.C(n_595),
.Y(n_848)
);

INVx5_ASAP7_75t_L g849 ( 
.A(n_672),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_675),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_671),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_672),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_665),
.B(n_590),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_624),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_675),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_700),
.B(n_595),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_606),
.B(n_374),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_701),
.A2(n_604),
.B1(n_601),
.B2(n_385),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_SL g859 ( 
.A(n_702),
.B(n_363),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_671),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_679),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_637),
.B(n_524),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_679),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_672),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_618),
.B(n_363),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_672),
.B(n_592),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_675),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_705),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_745),
.B(n_672),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_790),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_815),
.B(n_672),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_815),
.B(n_672),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_751),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_751),
.B(n_426),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_819),
.Y(n_875)
);

OR2x6_ASAP7_75t_L g876 ( 
.A(n_705),
.B(n_600),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_795),
.A2(n_684),
.B1(n_641),
.B2(n_390),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_SL g878 ( 
.A(n_718),
.B(n_358),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_795),
.Y(n_879)
);

OR2x6_ASAP7_75t_L g880 ( 
.A(n_816),
.B(n_600),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_SL g881 ( 
.A(n_718),
.B(n_782),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_715),
.B(n_637),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_740),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_790),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_740),
.B(n_752),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_752),
.A2(n_314),
.B1(n_337),
.B2(n_309),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_714),
.B(n_426),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_781),
.B(n_646),
.Y(n_888)
);

NAND2xp33_ASAP7_75t_L g889 ( 
.A(n_764),
.B(n_257),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_841),
.B(n_686),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_707),
.B(n_601),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_794),
.B(n_604),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_832),
.A2(n_684),
.B1(n_641),
.B2(n_392),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_761),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_723),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_SL g896 ( 
.A1(n_859),
.A2(n_720),
.B1(n_709),
.B2(n_708),
.Y(n_896)
);

INVx5_ASAP7_75t_L g897 ( 
.A(n_820),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_754),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_841),
.B(n_686),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_725),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_796),
.B(n_684),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_844),
.B(n_686),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_715),
.B(n_524),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_R g904 ( 
.A(n_750),
.B(n_624),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_754),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_791),
.Y(n_906)
);

NAND2x1_ASAP7_75t_L g907 ( 
.A(n_704),
.B(n_684),
.Y(n_907)
);

NOR2x2_ASAP7_75t_L g908 ( 
.A(n_832),
.B(n_394),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_732),
.A2(n_673),
.B(n_684),
.Y(n_909)
);

NAND2x1_ASAP7_75t_L g910 ( 
.A(n_704),
.B(n_682),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_842),
.B(n_253),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_739),
.A2(n_541),
.B(n_561),
.C(n_552),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_783),
.B(n_686),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_763),
.B(n_552),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_844),
.B(n_847),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_832),
.A2(n_397),
.B1(n_401),
.B2(n_384),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_SL g917 ( 
.A1(n_854),
.A2(n_750),
.B1(n_410),
.B2(n_439),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_847),
.B(n_686),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_762),
.A2(n_607),
.B(n_606),
.C(n_673),
.Y(n_919)
);

BUFx6f_ASAP7_75t_SL g920 ( 
.A(n_821),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_767),
.A2(n_771),
.B1(n_774),
.B2(n_773),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_748),
.B(n_686),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_832),
.A2(n_404),
.B1(n_414),
.B2(n_402),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_748),
.B(n_686),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_775),
.A2(n_607),
.B1(n_338),
.B2(n_345),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_856),
.B(n_256),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_763),
.B(n_682),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_772),
.B(n_388),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_729),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_SL g930 ( 
.A1(n_738),
.A2(n_462),
.B1(n_471),
.B2(n_396),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_772),
.B(n_717),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_714),
.B(n_683),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_848),
.A2(n_568),
.B(n_602),
.C(n_561),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_760),
.A2(n_607),
.B(n_496),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_791),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_735),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_735),
.B(n_568),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_818),
.B(n_683),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_754),
.B(n_426),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_768),
.Y(n_940)
);

NOR2x1p5_ASAP7_75t_L g941 ( 
.A(n_862),
.B(n_254),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_809),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_857),
.A2(n_338),
.B1(n_345),
.B2(n_337),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_809),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_816),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_810),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_742),
.A2(n_425),
.B1(n_429),
.B2(n_424),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_825),
.B(n_690),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_833),
.B(n_690),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_837),
.B(n_694),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_853),
.B(n_694),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_810),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_777),
.B(n_697),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_811),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_787),
.B(n_697),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_768),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_744),
.B(n_602),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_742),
.A2(n_443),
.B1(n_448),
.B2(n_432),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_845),
.B(n_408),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_811),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_728),
.A2(n_362),
.B1(n_395),
.B2(n_354),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_812),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_857),
.A2(n_708),
.B1(n_768),
.B2(n_724),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_760),
.A2(n_362),
.B1(n_395),
.B2(n_354),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_792),
.B(n_699),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_812),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_813),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_813),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_817),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_746),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_845),
.B(n_408),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_858),
.B(n_258),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_817),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_793),
.B(n_699),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_713),
.B(n_267),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_788),
.B(n_268),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_800),
.B(n_703),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_737),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_760),
.B(n_388),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_862),
.B(n_271),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_857),
.B(n_388),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_863),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_803),
.B(n_703),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_863),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_805),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_719),
.B(n_257),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_SL g987 ( 
.A(n_782),
.B(n_472),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_807),
.B(n_419),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_712),
.A2(n_446),
.B1(n_451),
.B2(n_419),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_808),
.B(n_824),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_802),
.A2(n_737),
.B1(n_708),
.B2(n_797),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_719),
.B(n_257),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_828),
.B(n_446),
.Y(n_993)
);

OR2x6_ASAP7_75t_L g994 ( 
.A(n_746),
.B(n_254),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_829),
.B(n_451),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_831),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_737),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_835),
.B(n_457),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_838),
.B(n_457),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_747),
.B(n_257),
.Y(n_1000)
);

AOI22x1_ASAP7_75t_L g1001 ( 
.A1(n_708),
.A2(n_466),
.B1(n_496),
.B2(n_493),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_724),
.A2(n_466),
.B1(n_372),
.B2(n_498),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_770),
.B(n_272),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_710),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_851),
.B(n_688),
.Y(n_1005)
);

BUFx12f_ASAP7_75t_L g1006 ( 
.A(n_821),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_747),
.B(n_257),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_724),
.A2(n_372),
.B1(n_501),
.B2(n_498),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_755),
.B(n_257),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_860),
.B(n_688),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_861),
.B(n_688),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_716),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_755),
.B(n_260),
.Y(n_1013)
);

INVxp67_ASAP7_75t_SL g1014 ( 
.A(n_710),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_744),
.B(n_408),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_731),
.B(n_501),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_865),
.B(n_273),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_733),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_757),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_766),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_776),
.B(n_280),
.Y(n_1021)
);

O2A1O1Ixp5_ASAP7_75t_L g1022 ( 
.A1(n_823),
.A2(n_852),
.B(n_827),
.C(n_801),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_710),
.B(n_515),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_823),
.B(n_685),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_823),
.B(n_685),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_852),
.B(n_685),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_710),
.B(n_515),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_836),
.B(n_292),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_839),
.A2(n_363),
.B1(n_599),
.B2(n_598),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_852),
.B(n_592),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_716),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_724),
.A2(n_765),
.B1(n_741),
.B2(n_786),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_785),
.A2(n_352),
.B(n_418),
.C(n_470),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_710),
.B(n_515),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_724),
.B(n_597),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_724),
.B(n_597),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_726),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_785),
.B(n_294),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_726),
.B(n_727),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_726),
.B(n_598),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_726),
.B(n_599),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_831),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_730),
.B(n_295),
.Y(n_1043)
);

INVxp67_ASAP7_75t_SL g1044 ( 
.A(n_873),
.Y(n_1044)
);

OR2x4_ASAP7_75t_L g1045 ( 
.A(n_972),
.B(n_329),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_870),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_892),
.B(n_741),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_996),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_905),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_914),
.B(n_741),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_870),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_905),
.Y(n_1052)
);

INVxp67_ASAP7_75t_SL g1053 ( 
.A(n_873),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_1001),
.A2(n_889),
.B1(n_896),
.B2(n_901),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_884),
.Y(n_1055)
);

INVxp33_ASAP7_75t_SL g1056 ( 
.A(n_881),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_905),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_884),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_945),
.Y(n_1059)
);

AND2x6_ASAP7_75t_SL g1060 ( 
.A(n_1043),
.B(n_333),
.Y(n_1060)
);

INVx3_ASAP7_75t_SL g1061 ( 
.A(n_1042),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_906),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_906),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_892),
.B(n_741),
.Y(n_1064)
);

AND2x4_ASAP7_75t_SL g1065 ( 
.A(n_970),
.B(n_821),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_928),
.A2(n_804),
.B(n_866),
.C(n_722),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_935),
.Y(n_1067)
);

NAND3xp33_ASAP7_75t_L g1068 ( 
.A(n_911),
.B(n_769),
.C(n_758),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_891),
.B(n_834),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_935),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_876),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_891),
.B(n_765),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_944),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_903),
.B(n_786),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_R g1075 ( 
.A(n_875),
.B(n_834),
.Y(n_1075)
);

AND2x6_ASAP7_75t_SL g1076 ( 
.A(n_1043),
.B(n_333),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_905),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_944),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_1006),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_946),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_946),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_876),
.Y(n_1082)
);

OR2x2_ASAP7_75t_SL g1083 ( 
.A(n_957),
.B(n_340),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_915),
.A2(n_827),
.B(n_801),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_931),
.B(n_765),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_937),
.Y(n_1086)
);

INVx5_ASAP7_75t_L g1087 ( 
.A(n_940),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_954),
.Y(n_1088)
);

CKINVDCx11_ASAP7_75t_R g1089 ( 
.A(n_1006),
.Y(n_1089)
);

NOR2xp67_ASAP7_75t_L g1090 ( 
.A(n_868),
.B(n_843),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_894),
.B(n_726),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_940),
.B(n_991),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_954),
.Y(n_1093)
);

NAND2xp33_ASAP7_75t_SL g1094 ( 
.A(n_888),
.B(n_706),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_978),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_940),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_940),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_960),
.Y(n_1098)
);

CKINVDCx16_ASAP7_75t_R g1099 ( 
.A(n_904),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_876),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_882),
.B(n_786),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_997),
.Y(n_1102)
);

INVx5_ASAP7_75t_L g1103 ( 
.A(n_1004),
.Y(n_1103)
);

INVx4_ASAP7_75t_L g1104 ( 
.A(n_1004),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_911),
.B(n_727),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_960),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_962),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_936),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_901),
.B(n_786),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_926),
.A2(n_779),
.B1(n_736),
.B2(n_834),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_962),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_926),
.B(n_727),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_969),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_927),
.B(n_727),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_921),
.B(n_727),
.Y(n_1115)
);

INVxp33_ASAP7_75t_L g1116 ( 
.A(n_904),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_898),
.B(n_743),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_942),
.B(n_749),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_1004),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_898),
.B(n_743),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_956),
.A2(n_827),
.B1(n_801),
.B2(n_780),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_880),
.Y(n_1122)
);

NOR3xp33_ASAP7_75t_SL g1123 ( 
.A(n_917),
.B(n_303),
.C(n_302),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_880),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_952),
.B(n_749),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_880),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_874),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_966),
.B(n_749),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_967),
.B(n_749),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_968),
.B(n_749),
.Y(n_1130)
);

INVx5_ASAP7_75t_L g1131 ( 
.A(n_1004),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_969),
.Y(n_1132)
);

NOR3xp33_ASAP7_75t_SL g1133 ( 
.A(n_930),
.B(n_311),
.C(n_307),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_R g1134 ( 
.A(n_878),
.B(n_711),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_982),
.B(n_780),
.Y(n_1135)
);

AND2x2_ASAP7_75t_SL g1136 ( 
.A(n_1032),
.B(n_372),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_956),
.B(n_778),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_972),
.A2(n_721),
.B1(n_734),
.B2(n_722),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_984),
.B(n_780),
.Y(n_1139)
);

CKINVDCx16_ASAP7_75t_R g1140 ( 
.A(n_920),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_973),
.Y(n_1141)
);

CKINVDCx8_ASAP7_75t_R g1142 ( 
.A(n_994),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1037),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_922),
.B(n_780),
.Y(n_1144)
);

NAND2x1p5_ASAP7_75t_L g1145 ( 
.A(n_897),
.B(n_780),
.Y(n_1145)
);

NOR3xp33_ASAP7_75t_SL g1146 ( 
.A(n_1033),
.B(n_980),
.C(n_976),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_924),
.B(n_789),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_973),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_907),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1012),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1012),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1037),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1031),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_879),
.A2(n_806),
.B1(n_864),
.B2(n_789),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_890),
.B(n_789),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1031),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_1037),
.Y(n_1157)
);

AOI21xp33_ASAP7_75t_L g1158 ( 
.A1(n_976),
.A2(n_315),
.B(n_313),
.Y(n_1158)
);

NOR3xp33_ASAP7_75t_SL g1159 ( 
.A(n_1033),
.B(n_323),
.C(n_318),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_SL g1160 ( 
.A1(n_980),
.A2(n_325),
.B1(n_326),
.B2(n_324),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1037),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1018),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_874),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_994),
.Y(n_1164)
);

INVxp67_ASAP7_75t_SL g1165 ( 
.A(n_885),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1019),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_899),
.B(n_789),
.Y(n_1167)
);

NOR3xp33_ASAP7_75t_SL g1168 ( 
.A(n_1003),
.B(n_332),
.C(n_327),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_941),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_994),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_963),
.A2(n_893),
.B1(n_883),
.B2(n_877),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1020),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_902),
.B(n_789),
.Y(n_1173)
);

NOR3xp33_ASAP7_75t_SL g1174 ( 
.A(n_1003),
.B(n_339),
.C(n_334),
.Y(n_1174)
);

INVx4_ASAP7_75t_L g1175 ( 
.A(n_897),
.Y(n_1175)
);

NOR3xp33_ASAP7_75t_L g1176 ( 
.A(n_888),
.B(n_344),
.C(n_343),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_918),
.B(n_806),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1013),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_939),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_928),
.A2(n_804),
.B(n_855),
.C(n_850),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_897),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_897),
.Y(n_1182)
);

INVxp33_ASAP7_75t_SL g1183 ( 
.A(n_987),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_985),
.B(n_806),
.Y(n_1184)
);

INVx4_ASAP7_75t_L g1185 ( 
.A(n_939),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1005),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_910),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_975),
.A2(n_806),
.B1(n_864),
.B2(n_820),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_990),
.B(n_806),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1013),
.Y(n_1190)
);

BUFx12f_ASAP7_75t_L g1191 ( 
.A(n_1015),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1013),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_895),
.Y(n_1193)
);

NOR3xp33_ASAP7_75t_SL g1194 ( 
.A(n_1038),
.B(n_356),
.C(n_355),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_939),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1017),
.B(n_864),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_900),
.Y(n_1197)
);

OR2x6_ASAP7_75t_L g1198 ( 
.A(n_874),
.B(n_372),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1010),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_975),
.A2(n_864),
.B1(n_820),
.B2(n_855),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1017),
.B(n_864),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1038),
.B(n_721),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_920),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_943),
.A2(n_867),
.B1(n_850),
.B2(n_759),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_R g1205 ( 
.A(n_1028),
.B(n_1021),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_887),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_929),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1028),
.A2(n_867),
.B(n_734),
.C(n_846),
.Y(n_1208)
);

CKINVDCx8_ASAP7_75t_R g1209 ( 
.A(n_887),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_887),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_871),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_872),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_947),
.B(n_778),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1011),
.Y(n_1214)
);

NOR3xp33_ASAP7_75t_SL g1215 ( 
.A(n_1021),
.B(n_361),
.C(n_357),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_913),
.B(n_869),
.Y(n_1216)
);

NAND3xp33_ASAP7_75t_L g1217 ( 
.A(n_961),
.B(n_366),
.C(n_365),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_959),
.B(n_753),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1016),
.Y(n_1219)
);

NAND2x1p5_ASAP7_75t_L g1220 ( 
.A(n_981),
.B(n_756),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1016),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1024),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1025),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1026),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_964),
.A2(n_784),
.B1(n_846),
.B2(n_840),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1014),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1040),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_908),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1041),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1030),
.Y(n_1230)
);

NAND3xp33_ASAP7_75t_SL g1231 ( 
.A(n_958),
.B(n_379),
.C(n_376),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_913),
.B(n_753),
.Y(n_1232)
);

INVxp67_ASAP7_75t_SL g1233 ( 
.A(n_1039),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_979),
.A2(n_820),
.B1(n_840),
.B2(n_830),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_953),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_971),
.B(n_759),
.Y(n_1236)
);

NOR3xp33_ASAP7_75t_SL g1237 ( 
.A(n_933),
.B(n_399),
.C(n_382),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_938),
.B(n_784),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1108),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1171),
.A2(n_1072),
.A3(n_919),
.B(n_1085),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1143),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1208),
.A2(n_909),
.A3(n_886),
.B(n_988),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1071),
.Y(n_1243)
);

CKINVDCx16_ASAP7_75t_R g1244 ( 
.A(n_1075),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1054),
.A2(n_979),
.B(n_934),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1115),
.A2(n_981),
.B(n_925),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1235),
.B(n_948),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1235),
.B(n_949),
.Y(n_1248)
);

NAND3xp33_ASAP7_75t_SL g1249 ( 
.A(n_1205),
.B(n_1029),
.C(n_923),
.Y(n_1249)
);

OA21x2_ASAP7_75t_L g1250 ( 
.A1(n_1216),
.A2(n_1022),
.B(n_992),
.Y(n_1250)
);

INVx4_ASAP7_75t_L g1251 ( 
.A(n_1077),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1149),
.A2(n_1039),
.B(n_992),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1175),
.A2(n_951),
.B(n_950),
.Y(n_1253)
);

NAND2x1_ASAP7_75t_L g1254 ( 
.A(n_1175),
.B(n_798),
.Y(n_1254)
);

INVxp67_ASAP7_75t_SL g1255 ( 
.A(n_1049),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1048),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1046),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1136),
.A2(n_916),
.B1(n_932),
.B2(n_1008),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1218),
.B(n_1236),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1218),
.B(n_912),
.Y(n_1260)
);

AOI21xp33_ASAP7_75t_L g1261 ( 
.A1(n_1068),
.A2(n_989),
.B(n_965),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_SL g1262 ( 
.A(n_1048),
.B(n_711),
.Y(n_1262)
);

OA22x2_ASAP7_75t_L g1263 ( 
.A1(n_1110),
.A2(n_442),
.B1(n_342),
.B2(n_346),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1086),
.B(n_993),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1236),
.B(n_955),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1047),
.A2(n_995),
.A3(n_998),
.B(n_999),
.Y(n_1266)
);

NAND2x1p5_ASAP7_75t_L g1267 ( 
.A(n_1077),
.B(n_1023),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1134),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1070),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1149),
.A2(n_1000),
.B(n_986),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1202),
.B(n_974),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1175),
.A2(n_1027),
.B(n_1023),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1082),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1100),
.Y(n_1274)
);

NAND2x1p5_ASAP7_75t_L g1275 ( 
.A(n_1077),
.B(n_1027),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1136),
.A2(n_977),
.B(n_983),
.C(n_1000),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1061),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1182),
.A2(n_1131),
.B(n_1103),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1070),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1077),
.B(n_986),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1209),
.A2(n_1002),
.B1(n_1035),
.B2(n_1036),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1182),
.A2(n_1034),
.B(n_849),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1182),
.A2(n_1034),
.B(n_849),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1127),
.B(n_1007),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_1077),
.Y(n_1285)
);

OR2x6_ASAP7_75t_L g1286 ( 
.A(n_1185),
.B(n_1009),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1164),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1209),
.A2(n_1009),
.B1(n_1007),
.B2(n_798),
.Y(n_1288)
);

AOI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1196),
.A2(n_814),
.B(n_799),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1144),
.A2(n_1147),
.B(n_1155),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1101),
.B(n_1074),
.Y(n_1291)
);

AO21x2_ASAP7_75t_L g1292 ( 
.A1(n_1092),
.A2(n_814),
.B(n_799),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1143),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1064),
.A2(n_830),
.A3(n_826),
.B(n_822),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1103),
.A2(n_849),
.B(n_756),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1164),
.Y(n_1296)
);

OA21x2_ASAP7_75t_L g1297 ( 
.A1(n_1167),
.A2(n_826),
.B(n_822),
.Y(n_1297)
);

BUFx4_ASAP7_75t_SL g1298 ( 
.A(n_1079),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1149),
.A2(n_596),
.B(n_529),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1103),
.A2(n_849),
.B(n_756),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1211),
.A2(n_596),
.B(n_529),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1211),
.A2(n_596),
.B(n_529),
.Y(n_1302)
);

AO22x1_ASAP7_75t_L g1303 ( 
.A1(n_1183),
.A2(n_473),
.B1(n_417),
.B2(n_415),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1202),
.B(n_778),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1143),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1103),
.A2(n_849),
.B(n_756),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1186),
.B(n_778),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1046),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1211),
.A2(n_1212),
.B(n_1232),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1101),
.B(n_260),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1212),
.A2(n_603),
.B(n_342),
.Y(n_1311)
);

O2A1O1Ixp5_ASAP7_75t_L g1312 ( 
.A1(n_1201),
.A2(n_413),
.B(n_367),
.C(n_470),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_SL g1313 ( 
.A(n_1079),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1212),
.A2(n_603),
.B(n_346),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1051),
.Y(n_1315)
);

AO31x2_ASAP7_75t_L g1316 ( 
.A1(n_1105),
.A2(n_418),
.A3(n_464),
.B(n_461),
.Y(n_1316)
);

AO21x2_ASAP7_75t_L g1317 ( 
.A1(n_1112),
.A2(n_352),
.B(n_340),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1173),
.A2(n_386),
.B(n_367),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1103),
.A2(n_756),
.B(n_820),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1177),
.A2(n_1114),
.B(n_1066),
.Y(n_1320)
);

INVx4_ASAP7_75t_L g1321 ( 
.A(n_1087),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1127),
.B(n_119),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1131),
.A2(n_820),
.B(n_398),
.Y(n_1323)
);

NAND3xp33_ASAP7_75t_SL g1324 ( 
.A(n_1176),
.B(n_405),
.C(n_403),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1094),
.A2(n_363),
.B1(n_468),
.B2(n_467),
.Y(n_1325)
);

OA21x2_ASAP7_75t_L g1326 ( 
.A1(n_1051),
.A2(n_398),
.B(n_386),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1165),
.A2(n_434),
.B1(n_465),
.B2(n_411),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1186),
.B(n_406),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1084),
.A2(n_400),
.B(n_464),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1180),
.A2(n_400),
.B(n_461),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1078),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1227),
.A2(n_409),
.B(n_460),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1199),
.B(n_407),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1219),
.A2(n_1221),
.B(n_1214),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1227),
.A2(n_1229),
.B(n_1081),
.Y(n_1335)
);

NOR2xp67_ASAP7_75t_L g1336 ( 
.A(n_1191),
.B(n_120),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1219),
.A2(n_413),
.B(n_420),
.Y(n_1337)
);

NAND2x1_ASAP7_75t_L g1338 ( 
.A(n_1104),
.B(n_409),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1227),
.A2(n_420),
.B(n_460),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1229),
.A2(n_1081),
.B(n_1078),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1146),
.A2(n_469),
.B(n_289),
.C(n_378),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1221),
.A2(n_440),
.B(n_437),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1131),
.A2(n_437),
.B(n_456),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1098),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1229),
.A2(n_440),
.B(n_456),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1049),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1143),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1199),
.A2(n_442),
.B(n_463),
.Y(n_1348)
);

O2A1O1Ixp33_ASAP7_75t_SL g1349 ( 
.A1(n_1213),
.A2(n_18),
.B(n_20),
.C(n_24),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1050),
.B(n_412),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1214),
.B(n_421),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1069),
.B(n_422),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1131),
.A2(n_469),
.B(n_445),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1098),
.A2(n_122),
.B(n_235),
.Y(n_1354)
);

OA22x2_ASAP7_75t_L g1355 ( 
.A1(n_1122),
.A2(n_459),
.B1(n_455),
.B2(n_454),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1107),
.A2(n_1148),
.B(n_1125),
.Y(n_1356)
);

AO21x2_ASAP7_75t_L g1357 ( 
.A1(n_1200),
.A2(n_186),
.B(n_125),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1107),
.A2(n_191),
.B(n_127),
.Y(n_1358)
);

AOI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1055),
.A2(n_1062),
.B(n_1058),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1148),
.A2(n_194),
.B(n_130),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1118),
.A2(n_197),
.B(n_134),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1055),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1091),
.A2(n_433),
.B(n_450),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1074),
.B(n_423),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1128),
.A2(n_1130),
.B(n_1129),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1135),
.A2(n_213),
.B(n_135),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_1087),
.B(n_427),
.Y(n_1367)
);

AND2x6_ASAP7_75t_L g1368 ( 
.A(n_1181),
.B(n_286),
.Y(n_1368)
);

A2O1A1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1050),
.A2(n_469),
.B(n_289),
.C(n_445),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1206),
.B(n_430),
.Y(n_1370)
);

NOR2xp67_ASAP7_75t_L g1371 ( 
.A(n_1191),
.B(n_123),
.Y(n_1371)
);

AO31x2_ASAP7_75t_L g1372 ( 
.A1(n_1058),
.A2(n_25),
.A3(n_27),
.B(n_30),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1062),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1193),
.B(n_431),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1131),
.A2(n_286),
.B(n_445),
.Y(n_1375)
);

OA22x2_ASAP7_75t_L g1376 ( 
.A1(n_1160),
.A2(n_449),
.B1(n_444),
.B2(n_438),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1193),
.B(n_435),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1139),
.A2(n_182),
.B(n_152),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1063),
.A2(n_216),
.B(n_153),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1087),
.B(n_436),
.Y(n_1380)
);

NAND2x1p5_ASAP7_75t_L g1381 ( 
.A(n_1087),
.B(n_391),
.Y(n_1381)
);

OA22x2_ASAP7_75t_L g1382 ( 
.A1(n_1124),
.A2(n_27),
.B1(n_30),
.B2(n_34),
.Y(n_1382)
);

AND2x2_ASAP7_75t_SL g1383 ( 
.A(n_1109),
.B(n_143),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1169),
.B(n_286),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1109),
.A2(n_391),
.B(n_378),
.C(n_289),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1197),
.B(n_1207),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1197),
.B(n_378),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1143),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1138),
.A2(n_391),
.B(n_232),
.Y(n_1389)
);

NAND2xp33_ASAP7_75t_L g1390 ( 
.A(n_1049),
.B(n_229),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1087),
.A2(n_223),
.B(n_222),
.Y(n_1391)
);

AOI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1063),
.A2(n_220),
.B(n_218),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1234),
.A2(n_217),
.B(n_178),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1067),
.A2(n_172),
.B(n_169),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1067),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1158),
.B(n_35),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1126),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1207),
.B(n_35),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1238),
.A2(n_166),
.B(n_165),
.Y(n_1399)
);

AO31x2_ASAP7_75t_L g1400 ( 
.A1(n_1073),
.A2(n_39),
.A3(n_42),
.B(n_44),
.Y(n_1400)
);

AO31x2_ASAP7_75t_L g1401 ( 
.A1(n_1073),
.A2(n_45),
.A3(n_46),
.B(n_47),
.Y(n_1401)
);

NOR2xp67_ASAP7_75t_SL g1402 ( 
.A(n_1142),
.B(n_47),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1099),
.B(n_49),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1210),
.A2(n_164),
.B1(n_157),
.B2(n_154),
.Y(n_1404)
);

INVxp67_ASAP7_75t_SL g1405 ( 
.A(n_1049),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1166),
.B(n_49),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1080),
.A2(n_51),
.B(n_52),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1166),
.B(n_52),
.Y(n_1408)
);

AO31x2_ASAP7_75t_L g1409 ( 
.A1(n_1341),
.A2(n_1106),
.A3(n_1113),
.B(n_1080),
.Y(n_1409)
);

BUFx12f_ASAP7_75t_L g1410 ( 
.A(n_1277),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1395),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1340),
.A2(n_1106),
.B(n_1088),
.Y(n_1412)
);

AO31x2_ASAP7_75t_L g1413 ( 
.A1(n_1341),
.A2(n_1088),
.A3(n_1113),
.B(n_1132),
.Y(n_1413)
);

AO31x2_ASAP7_75t_L g1414 ( 
.A1(n_1276),
.A2(n_1132),
.A3(n_1111),
.B(n_1093),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1396),
.B(n_1194),
.C(n_1215),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1251),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1359),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1269),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1348),
.A2(n_1231),
.B(n_1133),
.C(n_1174),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1247),
.B(n_1195),
.Y(n_1420)
);

AOI221xp5_ASAP7_75t_L g1421 ( 
.A1(n_1303),
.A2(n_1094),
.B1(n_1123),
.B2(n_1183),
.C(n_1228),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1248),
.B(n_1116),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1322),
.B(n_1195),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1271),
.B(n_1179),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1322),
.B(n_1210),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1340),
.A2(n_1093),
.B(n_1111),
.Y(n_1426)
);

AOI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1289),
.A2(n_1189),
.B(n_1141),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1259),
.A2(n_1226),
.B1(n_1163),
.B2(n_1044),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1335),
.A2(n_1141),
.B(n_1184),
.Y(n_1429)
);

INVx2_ASAP7_75t_SL g1430 ( 
.A(n_1239),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1291),
.B(n_1364),
.Y(n_1431)
);

AO21x2_ASAP7_75t_L g1432 ( 
.A1(n_1389),
.A2(n_1154),
.B(n_1188),
.Y(n_1432)
);

OAI211xp5_ASAP7_75t_SL g1433 ( 
.A1(n_1325),
.A2(n_1168),
.B(n_1237),
.C(n_1159),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1276),
.A2(n_1233),
.B(n_1162),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1335),
.A2(n_1222),
.B(n_1223),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1386),
.Y(n_1436)
);

NAND2x1p5_ASAP7_75t_L g1437 ( 
.A(n_1251),
.B(n_1049),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1239),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_L g1439 ( 
.A(n_1352),
.B(n_1261),
.C(n_1402),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1269),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1356),
.A2(n_1222),
.B(n_1223),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_1244),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1257),
.Y(n_1443)
);

NOR4xp25_ASAP7_75t_L g1444 ( 
.A(n_1249),
.B(n_1217),
.C(n_1060),
.D(n_1076),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1356),
.A2(n_1224),
.B(n_1225),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1287),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1308),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1265),
.B(n_1291),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1258),
.A2(n_1162),
.B(n_1230),
.Y(n_1449)
);

OAI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1352),
.A2(n_1228),
.B1(n_1090),
.B2(n_1328),
.C(n_1333),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1296),
.Y(n_1451)
);

O2A1O1Ixp33_ASAP7_75t_L g1452 ( 
.A1(n_1369),
.A2(n_1170),
.B(n_1056),
.C(n_1172),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1301),
.A2(n_1224),
.B(n_1150),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1315),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1362),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1279),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1301),
.A2(n_1302),
.B(n_1309),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1245),
.A2(n_1226),
.B1(n_1163),
.B2(n_1053),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1383),
.B(n_1178),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1383),
.B(n_1178),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1302),
.A2(n_1309),
.B(n_1299),
.Y(n_1461)
);

BUFx8_ASAP7_75t_L g1462 ( 
.A(n_1313),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1256),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1273),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1331),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1256),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1322),
.B(n_1284),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1331),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1344),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1344),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1393),
.A2(n_1172),
.B(n_1190),
.C(n_1192),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1260),
.B(n_1083),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_1277),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1264),
.B(n_1117),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1310),
.B(n_1117),
.Y(n_1475)
);

OR2x6_ASAP7_75t_L g1476 ( 
.A(n_1334),
.B(n_1286),
.Y(n_1476)
);

NAND2x1p5_ASAP7_75t_L g1477 ( 
.A(n_1251),
.B(n_1052),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1373),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1241),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1284),
.B(n_1117),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1246),
.A2(n_1226),
.B1(n_1190),
.B2(n_1185),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1284),
.B(n_1120),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1299),
.A2(n_1151),
.B(n_1150),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1292),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1253),
.A2(n_1230),
.B(n_1192),
.Y(n_1485)
);

OAI221xp5_ASAP7_75t_L g1486 ( 
.A1(n_1351),
.A2(n_1142),
.B1(n_1059),
.B2(n_1045),
.C(n_1203),
.Y(n_1486)
);

BUFx2_ASAP7_75t_R g1487 ( 
.A(n_1268),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1274),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1298),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1292),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1387),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1311),
.A2(n_1151),
.B(n_1220),
.Y(n_1492)
);

AO21x2_ASAP7_75t_L g1493 ( 
.A1(n_1320),
.A2(n_1121),
.B(n_1156),
.Y(n_1493)
);

NOR2xp67_ASAP7_75t_L g1494 ( 
.A(n_1268),
.B(n_1059),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1241),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1281),
.A2(n_1204),
.B(n_1190),
.Y(n_1496)
);

OAI211xp5_ASAP7_75t_SL g1497 ( 
.A1(n_1403),
.A2(n_1089),
.B(n_1045),
.C(n_1083),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1266),
.B(n_1120),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1311),
.A2(n_1220),
.B(n_1152),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1310),
.B(n_1198),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1243),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1326),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1397),
.B(n_1056),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1314),
.A2(n_1220),
.B(n_1152),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1255),
.A2(n_1405),
.B1(n_1185),
.B2(n_1045),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1314),
.A2(n_1161),
.B(n_1157),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1326),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1350),
.B(n_1198),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1326),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1374),
.B(n_1120),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1294),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1294),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1290),
.A2(n_1181),
.B(n_1145),
.Y(n_1513)
);

AO31x2_ASAP7_75t_L g1514 ( 
.A1(n_1385),
.A2(n_1156),
.A3(n_1153),
.B(n_1119),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1241),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1294),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1285),
.B(n_1095),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1286),
.A2(n_1052),
.B1(n_1057),
.B2(n_1097),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1398),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1294),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1406),
.Y(n_1521)
);

NAND2x1p5_ASAP7_75t_L g1522 ( 
.A(n_1285),
.B(n_1052),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1408),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1329),
.A2(n_1365),
.B(n_1330),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1337),
.B(n_1198),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1332),
.Y(n_1526)
);

OAI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1262),
.A2(n_1140),
.B1(n_1203),
.B2(n_1095),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_SL g1528 ( 
.A1(n_1392),
.A2(n_1119),
.B(n_1104),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1241),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1377),
.B(n_1102),
.Y(n_1530)
);

INVx2_ASAP7_75t_SL g1531 ( 
.A(n_1293),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1329),
.A2(n_1365),
.B(n_1330),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1285),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1332),
.Y(n_1534)
);

AND2x6_ASAP7_75t_L g1535 ( 
.A(n_1293),
.B(n_1052),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1339),
.Y(n_1536)
);

O2A1O1Ixp33_ASAP7_75t_SL g1537 ( 
.A1(n_1385),
.A2(n_1369),
.B(n_1367),
.C(n_1380),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1293),
.Y(n_1538)
);

AO21x2_ASAP7_75t_L g1539 ( 
.A1(n_1318),
.A2(n_1153),
.B(n_1137),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1370),
.B(n_1102),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1324),
.A2(n_1198),
.B1(n_1096),
.B2(n_1052),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1339),
.A2(n_1161),
.B(n_1157),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1321),
.B(n_1096),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1321),
.A2(n_1181),
.B(n_1145),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1338),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1345),
.A2(n_1161),
.B(n_1157),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1321),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1263),
.Y(n_1548)
);

OAI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1312),
.A2(n_1096),
.B(n_1137),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_SL g1550 ( 
.A1(n_1399),
.A2(n_1119),
.B(n_1104),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1345),
.A2(n_1152),
.B(n_1145),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1297),
.Y(n_1552)
);

NAND2xp33_ASAP7_75t_L g1553 ( 
.A(n_1293),
.B(n_1057),
.Y(n_1553)
);

O2A1O1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1342),
.A2(n_1061),
.B(n_1137),
.C(n_1065),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1266),
.B(n_1240),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1266),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1266),
.Y(n_1557)
);

OAI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1304),
.A2(n_1187),
.B(n_1097),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1327),
.B(n_1065),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1305),
.Y(n_1560)
);

AOI222xp33_ASAP7_75t_L g1561 ( 
.A1(n_1384),
.A2(n_1089),
.B1(n_1097),
.B2(n_1057),
.C1(n_1187),
.C2(n_63),
.Y(n_1561)
);

INVx3_ASAP7_75t_L g1562 ( 
.A(n_1305),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1305),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1297),
.Y(n_1564)
);

AO31x2_ASAP7_75t_L g1565 ( 
.A1(n_1288),
.A2(n_1187),
.A3(n_1097),
.B(n_1057),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_SL g1566 ( 
.A1(n_1391),
.A2(n_1097),
.B(n_1057),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1305),
.Y(n_1567)
);

NOR3xp33_ASAP7_75t_SL g1568 ( 
.A(n_1363),
.B(n_53),
.C(n_58),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1252),
.A2(n_1187),
.B(n_1181),
.Y(n_1569)
);

AOI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1390),
.A2(n_1181),
.B(n_1187),
.Y(n_1570)
);

OAI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1270),
.A2(n_117),
.B(n_62),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1263),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1252),
.A2(n_60),
.B(n_65),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1354),
.A2(n_67),
.B(n_68),
.Y(n_1574)
);

OAI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1270),
.A2(n_115),
.B(n_73),
.Y(n_1575)
);

OR2x6_ASAP7_75t_L g1576 ( 
.A(n_1286),
.B(n_72),
.Y(n_1576)
);

A2O1A1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1390),
.A2(n_73),
.B(n_74),
.C(n_75),
.Y(n_1577)
);

O2A1O1Ixp33_ASAP7_75t_SL g1578 ( 
.A1(n_1367),
.A2(n_76),
.B(n_78),
.C(n_81),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1313),
.Y(n_1579)
);

AO21x2_ASAP7_75t_L g1580 ( 
.A1(n_1318),
.A2(n_76),
.B(n_81),
.Y(n_1580)
);

A2O1A1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1380),
.A2(n_84),
.B(n_85),
.C(n_87),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1382),
.B(n_84),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1280),
.A2(n_1272),
.B(n_1278),
.Y(n_1583)
);

OAI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1354),
.A2(n_1360),
.B(n_1358),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1297),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1347),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1286),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1250),
.Y(n_1588)
);

A2O1A1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1343),
.A2(n_88),
.B(n_90),
.C(n_91),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1346),
.B(n_91),
.Y(n_1590)
);

OAI21x1_ASAP7_75t_L g1591 ( 
.A1(n_1358),
.A2(n_93),
.B(n_94),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1376),
.B(n_93),
.Y(n_1592)
);

OAI21x1_ASAP7_75t_L g1593 ( 
.A1(n_1360),
.A2(n_94),
.B(n_95),
.Y(n_1593)
);

BUFx8_ASAP7_75t_SL g1594 ( 
.A(n_1489),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1443),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1570),
.A2(n_1280),
.B(n_1250),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_L g1597 ( 
.A(n_1479),
.Y(n_1597)
);

AND2x6_ASAP7_75t_L g1598 ( 
.A(n_1459),
.B(n_1460),
.Y(n_1598)
);

A2O1A1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1439),
.A2(n_1407),
.B(n_1371),
.C(n_1336),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1422),
.B(n_1376),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1447),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_1479),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1561),
.A2(n_1382),
.B1(n_1355),
.B2(n_1404),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1409),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1409),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1448),
.B(n_1240),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_SL g1607 ( 
.A(n_1487),
.B(n_1313),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1582),
.B(n_1355),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1517),
.Y(n_1609)
);

OAI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1576),
.A2(n_1472),
.B1(n_1431),
.B2(n_1450),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1409),
.Y(n_1611)
);

OR2x6_ASAP7_75t_L g1612 ( 
.A(n_1576),
.B(n_1379),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1521),
.B(n_1240),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1444),
.A2(n_1349),
.B1(n_1353),
.B2(n_1375),
.C(n_1317),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1454),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1464),
.Y(n_1616)
);

AOI221xp5_ASAP7_75t_L g1617 ( 
.A1(n_1592),
.A2(n_1349),
.B1(n_1317),
.B2(n_1357),
.C(n_1307),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1472),
.A2(n_1381),
.B1(n_1346),
.B2(n_1275),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1582),
.A2(n_1357),
.B1(n_1407),
.B2(n_1368),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1423),
.B(n_1425),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1455),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1478),
.Y(n_1622)
);

NAND3xp33_ASAP7_75t_L g1623 ( 
.A(n_1568),
.B(n_1323),
.C(n_1250),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1431),
.B(n_1381),
.Y(n_1624)
);

A2O1A1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1571),
.A2(n_1379),
.B(n_1394),
.C(n_1366),
.Y(n_1625)
);

AOI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1419),
.A2(n_1283),
.B1(n_1282),
.B2(n_1347),
.C(n_1388),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1478),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1411),
.Y(n_1628)
);

INVx4_ASAP7_75t_L g1629 ( 
.A(n_1489),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1523),
.B(n_1240),
.Y(n_1630)
);

A2O1A1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1575),
.A2(n_1394),
.B(n_1378),
.C(n_1361),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1587),
.A2(n_1368),
.B1(n_1378),
.B2(n_1366),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1420),
.B(n_1316),
.Y(n_1633)
);

NAND2xp33_ASAP7_75t_R g1634 ( 
.A(n_1459),
.B(n_1361),
.Y(n_1634)
);

OR2x6_ASAP7_75t_L g1635 ( 
.A(n_1576),
.B(n_1347),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1411),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1418),
.Y(n_1637)
);

OAI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1449),
.A2(n_1368),
.B(n_1267),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1474),
.B(n_1316),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1475),
.B(n_1275),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_SL g1641 ( 
.A1(n_1576),
.A2(n_1368),
.B1(n_1400),
.B2(n_1372),
.Y(n_1641)
);

OA21x2_ASAP7_75t_L g1642 ( 
.A1(n_1524),
.A2(n_1319),
.B(n_1316),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1503),
.A2(n_1267),
.B1(n_1388),
.B2(n_1347),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1468),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1423),
.A2(n_1388),
.B1(n_1254),
.B2(n_1295),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1468),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_1410),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1423),
.A2(n_1388),
.B1(n_1300),
.B2(n_1306),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_SL g1649 ( 
.A(n_1410),
.B(n_1368),
.Y(n_1649)
);

OR2x6_ASAP7_75t_L g1650 ( 
.A(n_1554),
.B(n_1401),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1467),
.B(n_1480),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1424),
.B(n_1316),
.Y(n_1652)
);

BUFx12f_ASAP7_75t_L g1653 ( 
.A(n_1462),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1446),
.B(n_1401),
.Y(n_1654)
);

CKINVDCx16_ASAP7_75t_R g1655 ( 
.A(n_1442),
.Y(n_1655)
);

INVx3_ASAP7_75t_L g1656 ( 
.A(n_1517),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1479),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1433),
.A2(n_1401),
.B1(n_1400),
.B2(n_1372),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1471),
.A2(n_1242),
.B(n_1400),
.Y(n_1659)
);

AOI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1485),
.A2(n_1242),
.B(n_1400),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1425),
.B(n_1242),
.Y(n_1661)
);

BUFx4f_ASAP7_75t_SL g1662 ( 
.A(n_1462),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1440),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1446),
.Y(n_1664)
);

OR2x6_ASAP7_75t_L g1665 ( 
.A(n_1476),
.B(n_1467),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1425),
.B(n_1242),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1519),
.B(n_1401),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1460),
.B(n_1372),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1553),
.A2(n_1372),
.B(n_96),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1553),
.A2(n_95),
.B(n_96),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1469),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1469),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1548),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1479),
.Y(n_1674)
);

NAND2x1p5_ASAP7_75t_L g1675 ( 
.A(n_1416),
.B(n_100),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1470),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_SL g1677 ( 
.A1(n_1590),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1572),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1436),
.B(n_109),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1470),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1510),
.B(n_111),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1456),
.Y(n_1682)
);

OAI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1584),
.A2(n_115),
.B(n_113),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1480),
.B(n_113),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1409),
.Y(n_1685)
);

NAND2xp33_ASAP7_75t_R g1686 ( 
.A(n_1525),
.B(n_114),
.Y(n_1686)
);

INVx5_ASAP7_75t_L g1687 ( 
.A(n_1535),
.Y(n_1687)
);

AOI21x1_ASAP7_75t_L g1688 ( 
.A1(n_1427),
.A2(n_1583),
.B(n_1526),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1451),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1480),
.B(n_1482),
.Y(n_1690)
);

O2A1O1Ixp33_ASAP7_75t_SL g1691 ( 
.A1(n_1577),
.A2(n_1581),
.B(n_1589),
.C(n_1452),
.Y(n_1691)
);

INVx3_ASAP7_75t_L g1692 ( 
.A(n_1517),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1543),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1530),
.B(n_1451),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1421),
.A2(n_1540),
.B1(n_1415),
.B2(n_1497),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1491),
.B(n_1482),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_1442),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1456),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1482),
.B(n_1579),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1501),
.Y(n_1700)
);

AO31x2_ASAP7_75t_L g1701 ( 
.A1(n_1511),
.A2(n_1516),
.A3(n_1520),
.B(n_1512),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1465),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1488),
.B(n_1501),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_R g1704 ( 
.A(n_1463),
.B(n_1466),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1476),
.A2(n_1559),
.B1(n_1486),
.B2(n_1541),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1409),
.Y(n_1706)
);

NAND2x1p5_ASAP7_75t_L g1707 ( 
.A(n_1416),
.B(n_1533),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_SL g1708 ( 
.A1(n_1590),
.A2(n_1432),
.B1(n_1496),
.B2(n_1462),
.Y(n_1708)
);

CKINVDCx14_ASAP7_75t_R g1709 ( 
.A(n_1463),
.Y(n_1709)
);

A2O1A1Ixp33_ASAP7_75t_SL g1710 ( 
.A1(n_1434),
.A2(n_1558),
.B(n_1549),
.C(n_1556),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1438),
.B(n_1430),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1465),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1508),
.B(n_1500),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1430),
.B(n_1466),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1498),
.B(n_1473),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1494),
.B(n_1473),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1417),
.Y(n_1717)
);

INVx4_ASAP7_75t_L g1718 ( 
.A(n_1535),
.Y(n_1718)
);

CKINVDCx6p67_ASAP7_75t_R g1719 ( 
.A(n_1515),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1412),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1508),
.A2(n_1432),
.B1(n_1590),
.B2(n_1476),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1498),
.B(n_1500),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1413),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_SL g1724 ( 
.A1(n_1432),
.A2(n_1580),
.B1(n_1505),
.B2(n_1573),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1527),
.B(n_1537),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1426),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1580),
.A2(n_1493),
.B1(n_1556),
.B2(n_1557),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1529),
.B(n_1560),
.Y(n_1728)
);

AO21x2_ASAP7_75t_L g1729 ( 
.A1(n_1584),
.A2(n_1524),
.B(n_1532),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1518),
.A2(n_1428),
.B1(n_1458),
.B2(n_1481),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1560),
.B(n_1567),
.Y(n_1731)
);

NAND3xp33_ASAP7_75t_SL g1732 ( 
.A(n_1545),
.B(n_1513),
.C(n_1522),
.Y(n_1732)
);

INVx2_ASAP7_75t_SL g1733 ( 
.A(n_1586),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1580),
.A2(n_1493),
.B1(n_1557),
.B2(n_1555),
.Y(n_1734)
);

NAND2xp33_ASAP7_75t_R g1735 ( 
.A(n_1416),
.B(n_1533),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1437),
.A2(n_1477),
.B1(n_1522),
.B2(n_1567),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_1543),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_SL g1738 ( 
.A(n_1543),
.B(n_1529),
.Y(n_1738)
);

OAI21xp33_ASAP7_75t_L g1739 ( 
.A1(n_1573),
.A2(n_1512),
.B(n_1516),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1426),
.Y(n_1740)
);

NAND2xp33_ASAP7_75t_R g1741 ( 
.A(n_1533),
.B(n_1547),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1413),
.B(n_1414),
.Y(n_1742)
);

CKINVDCx16_ASAP7_75t_R g1743 ( 
.A(n_1586),
.Y(n_1743)
);

OAI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1507),
.A2(n_1509),
.B1(n_1502),
.B2(n_1520),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1437),
.A2(n_1477),
.B1(n_1522),
.B2(n_1547),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1437),
.A2(n_1477),
.B1(n_1547),
.B2(n_1562),
.Y(n_1746)
);

OAI21x1_ASAP7_75t_L g1747 ( 
.A1(n_1457),
.A2(n_1461),
.B(n_1441),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1435),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1562),
.B(n_1563),
.Y(n_1749)
);

OAI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1507),
.A2(n_1509),
.B1(n_1502),
.B2(n_1534),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1563),
.B(n_1531),
.Y(n_1751)
);

AOI221xp5_ASAP7_75t_SL g1752 ( 
.A1(n_1526),
.A2(n_1534),
.B1(n_1536),
.B2(n_1544),
.C(n_1495),
.Y(n_1752)
);

A2O1A1Ixp33_ASAP7_75t_L g1753 ( 
.A1(n_1574),
.A2(n_1593),
.B(n_1591),
.C(n_1445),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1435),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1413),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1479),
.Y(n_1756)
);

NAND3xp33_ASAP7_75t_L g1757 ( 
.A(n_1578),
.B(n_1536),
.C(n_1490),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1495),
.Y(n_1758)
);

CKINVDCx6p67_ASAP7_75t_R g1759 ( 
.A(n_1495),
.Y(n_1759)
);

INVx4_ASAP7_75t_L g1760 ( 
.A(n_1535),
.Y(n_1760)
);

BUFx12f_ASAP7_75t_L g1761 ( 
.A(n_1495),
.Y(n_1761)
);

OAI21xp5_ASAP7_75t_SL g1762 ( 
.A1(n_1531),
.A2(n_1538),
.B(n_1427),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1413),
.B(n_1414),
.Y(n_1763)
);

AO21x2_ASAP7_75t_L g1764 ( 
.A1(n_1532),
.A2(n_1550),
.B(n_1528),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1495),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1538),
.B(n_1514),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1514),
.B(n_1413),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1484),
.A2(n_1490),
.B1(n_1588),
.B2(n_1585),
.Y(n_1768)
);

INVxp33_ASAP7_75t_L g1769 ( 
.A(n_1542),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1535),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1514),
.Y(n_1771)
);

INVx4_ASAP7_75t_L g1772 ( 
.A(n_1535),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1414),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1493),
.A2(n_1550),
.B1(n_1574),
.B2(n_1591),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1514),
.B(n_1414),
.Y(n_1775)
);

A2O1A1Ixp33_ASAP7_75t_L g1776 ( 
.A1(n_1593),
.A2(n_1445),
.B(n_1441),
.C(n_1429),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1535),
.A2(n_1539),
.B1(n_1484),
.B2(n_1551),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1414),
.Y(n_1778)
);

BUFx12f_ASAP7_75t_L g1779 ( 
.A(n_1566),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1483),
.Y(n_1780)
);

O2A1O1Ixp33_ASAP7_75t_L g1781 ( 
.A1(n_1566),
.A2(n_1528),
.B(n_1539),
.C(n_1564),
.Y(n_1781)
);

OAI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1588),
.A2(n_1585),
.B1(n_1564),
.B2(n_1552),
.Y(n_1782)
);

INVx3_ASAP7_75t_L g1783 ( 
.A(n_1514),
.Y(n_1783)
);

NOR2x1_ASAP7_75t_SL g1784 ( 
.A(n_1539),
.B(n_1552),
.Y(n_1784)
);

INVx2_ASAP7_75t_SL g1785 ( 
.A(n_1565),
.Y(n_1785)
);

BUFx2_ASAP7_75t_L g1786 ( 
.A(n_1565),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1429),
.A2(n_1483),
.B1(n_1453),
.B2(n_1492),
.Y(n_1787)
);

AOI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1453),
.A2(n_1492),
.B1(n_1546),
.B2(n_1542),
.Y(n_1788)
);

OAI211xp5_ASAP7_75t_L g1789 ( 
.A1(n_1546),
.A2(n_1506),
.B(n_1504),
.C(n_1499),
.Y(n_1789)
);

OAI21xp33_ASAP7_75t_L g1790 ( 
.A1(n_1603),
.A2(n_1506),
.B(n_1504),
.Y(n_1790)
);

OAI211xp5_ASAP7_75t_SL g1791 ( 
.A1(n_1695),
.A2(n_1565),
.B(n_1499),
.C(n_1569),
.Y(n_1791)
);

OAI221xp5_ASAP7_75t_L g1792 ( 
.A1(n_1603),
.A2(n_1565),
.B1(n_1569),
.B2(n_1551),
.C(n_1457),
.Y(n_1792)
);

AOI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1691),
.A2(n_1461),
.B1(n_1565),
.B2(n_1610),
.C(n_1673),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1673),
.A2(n_1678),
.B1(n_1681),
.B2(n_1677),
.Y(n_1794)
);

INVx3_ASAP7_75t_L g1795 ( 
.A(n_1761),
.Y(n_1795)
);

OAI211xp5_ASAP7_75t_L g1796 ( 
.A1(n_1678),
.A2(n_1677),
.B(n_1670),
.C(n_1681),
.Y(n_1796)
);

OAI22xp33_ASAP7_75t_SL g1797 ( 
.A1(n_1725),
.A2(n_1705),
.B1(n_1675),
.B2(n_1650),
.Y(n_1797)
);

NOR3xp33_ASAP7_75t_L g1798 ( 
.A(n_1610),
.B(n_1600),
.C(n_1691),
.Y(n_1798)
);

AOI21xp33_ASAP7_75t_L g1799 ( 
.A1(n_1624),
.A2(n_1640),
.B(n_1652),
.Y(n_1799)
);

BUFx2_ASAP7_75t_L g1800 ( 
.A(n_1700),
.Y(n_1800)
);

OAI33xp33_ASAP7_75t_L g1801 ( 
.A1(n_1679),
.A2(n_1654),
.A3(n_1667),
.B1(n_1616),
.B2(n_1668),
.B3(n_1621),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1694),
.B(n_1696),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1635),
.A2(n_1708),
.B1(n_1709),
.B2(n_1714),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1622),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1708),
.A2(n_1694),
.B1(n_1639),
.B2(n_1684),
.Y(n_1805)
);

OAI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1635),
.A2(n_1709),
.B1(n_1715),
.B2(n_1664),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1731),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1701),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1616),
.B(n_1689),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1624),
.A2(n_1662),
.B1(n_1699),
.B2(n_1653),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1703),
.B(n_1651),
.Y(n_1811)
);

OAI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1686),
.A2(n_1635),
.B1(n_1735),
.B2(n_1741),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1722),
.B(n_1728),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1662),
.A2(n_1699),
.B1(n_1669),
.B2(n_1614),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1633),
.B(n_1613),
.Y(n_1815)
);

BUFx2_ASAP7_75t_L g1816 ( 
.A(n_1704),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1630),
.B(n_1606),
.Y(n_1817)
);

OR2x6_ASAP7_75t_L g1818 ( 
.A(n_1665),
.B(n_1779),
.Y(n_1818)
);

OAI221xp5_ASAP7_75t_L g1819 ( 
.A1(n_1686),
.A2(n_1599),
.B1(n_1617),
.B2(n_1632),
.C(n_1675),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1627),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1730),
.A2(n_1658),
.B1(n_1641),
.B2(n_1650),
.Y(n_1821)
);

AOI221xp5_ASAP7_75t_L g1822 ( 
.A1(n_1658),
.A2(n_1660),
.B1(n_1659),
.B2(n_1641),
.C(n_1668),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1717),
.Y(n_1823)
);

OAI221xp5_ASAP7_75t_L g1824 ( 
.A1(n_1599),
.A2(n_1632),
.B1(n_1638),
.B2(n_1619),
.C(n_1649),
.Y(n_1824)
);

OAI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1735),
.A2(n_1741),
.B1(n_1607),
.B2(n_1738),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1620),
.B(n_1711),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1620),
.B(n_1609),
.Y(n_1827)
);

AOI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1623),
.A2(n_1619),
.B1(n_1710),
.B2(n_1721),
.C(n_1734),
.Y(n_1828)
);

INVxp67_ASAP7_75t_L g1829 ( 
.A(n_1595),
.Y(n_1829)
);

OAI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1640),
.A2(n_1724),
.B1(n_1625),
.B2(n_1631),
.C(n_1626),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1721),
.A2(n_1716),
.B1(n_1743),
.B2(n_1770),
.Y(n_1831)
);

INVxp67_ASAP7_75t_SL g1832 ( 
.A(n_1750),
.Y(n_1832)
);

OAI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1716),
.A2(n_1697),
.B1(n_1650),
.B2(n_1643),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1601),
.A2(n_1615),
.B1(n_1661),
.B2(n_1666),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1661),
.A2(n_1666),
.B1(n_1690),
.B2(n_1665),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1690),
.A2(n_1665),
.B1(n_1598),
.B2(n_1612),
.Y(n_1836)
);

OA21x2_ASAP7_75t_L g1837 ( 
.A1(n_1776),
.A2(n_1752),
.B(n_1625),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1598),
.A2(n_1612),
.B1(n_1629),
.B2(n_1628),
.Y(n_1838)
);

OAI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1687),
.A2(n_1656),
.B1(n_1692),
.B2(n_1719),
.Y(n_1839)
);

AOI222xp33_ASAP7_75t_L g1840 ( 
.A1(n_1598),
.A2(n_1618),
.B1(n_1710),
.B2(n_1647),
.C1(n_1629),
.C2(n_1636),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1732),
.A2(n_1693),
.B1(n_1737),
.B2(n_1634),
.Y(n_1841)
);

OA21x2_ASAP7_75t_L g1842 ( 
.A1(n_1776),
.A2(n_1753),
.B(n_1631),
.Y(n_1842)
);

AOI221xp5_ASAP7_75t_L g1843 ( 
.A1(n_1734),
.A2(n_1724),
.B1(n_1774),
.B2(n_1727),
.C(n_1773),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1693),
.B(n_1737),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1612),
.A2(n_1671),
.B1(n_1646),
.B2(n_1672),
.Y(n_1845)
);

INVx5_ASAP7_75t_SL g1846 ( 
.A(n_1759),
.Y(n_1846)
);

OAI221xp5_ASAP7_75t_SL g1847 ( 
.A1(n_1774),
.A2(n_1753),
.B1(n_1727),
.B2(n_1762),
.C(n_1596),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_SL g1848 ( 
.A(n_1594),
.B(n_1756),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1644),
.B(n_1676),
.Y(n_1849)
);

OAI222xp33_ASAP7_75t_L g1850 ( 
.A1(n_1718),
.A2(n_1772),
.B1(n_1760),
.B2(n_1680),
.C1(n_1786),
.C2(n_1749),
.Y(n_1850)
);

OAI211xp5_ASAP7_75t_L g1851 ( 
.A1(n_1683),
.A2(n_1739),
.B(n_1757),
.C(n_1763),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1637),
.B(n_1663),
.Y(n_1852)
);

NOR2x1_ASAP7_75t_L g1853 ( 
.A(n_1751),
.B(n_1765),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1687),
.A2(n_1772),
.B1(n_1760),
.B2(n_1718),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1687),
.A2(n_1733),
.B1(n_1707),
.B2(n_1736),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_SL g1856 ( 
.A1(n_1745),
.A2(n_1775),
.B(n_1777),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_SL g1857 ( 
.A1(n_1648),
.A2(n_1645),
.B1(n_1746),
.B2(n_1767),
.Y(n_1857)
);

AOI222xp33_ASAP7_75t_L g1858 ( 
.A1(n_1682),
.A2(n_1712),
.B1(n_1702),
.B2(n_1698),
.C1(n_1778),
.C2(n_1742),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1634),
.A2(n_1766),
.B1(n_1764),
.B2(n_1707),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1701),
.B(n_1723),
.Y(n_1860)
);

AO21x2_ASAP7_75t_L g1861 ( 
.A1(n_1688),
.A2(n_1789),
.B(n_1750),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1597),
.B(n_1758),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_SL g1863 ( 
.A1(n_1785),
.A2(n_1771),
.B1(n_1723),
.B2(n_1685),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1597),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_SL g1865 ( 
.A1(n_1771),
.A2(n_1706),
.B1(n_1604),
.B2(n_1605),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1701),
.B(n_1611),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_SL g1867 ( 
.A1(n_1604),
.A2(n_1706),
.B1(n_1605),
.B2(n_1611),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1602),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_R g1869 ( 
.A(n_1602),
.B(n_1758),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1602),
.B(n_1657),
.Y(n_1870)
);

OAI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1755),
.A2(n_1685),
.B1(n_1602),
.B2(n_1657),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1768),
.Y(n_1872)
);

O2A1O1Ixp33_ASAP7_75t_L g1873 ( 
.A1(n_1781),
.A2(n_1783),
.B(n_1740),
.C(n_1720),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1657),
.B(n_1674),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1594),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1764),
.A2(n_1657),
.B1(n_1674),
.B2(n_1783),
.Y(n_1876)
);

AOI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1744),
.A2(n_1784),
.B(n_1787),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1782),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1787),
.A2(n_1674),
.B1(n_1788),
.B2(n_1769),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1726),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1780),
.A2(n_1748),
.B1(n_1754),
.B2(n_1744),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1642),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1642),
.A2(n_1769),
.B1(n_1729),
.B2(n_1788),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1747),
.B(n_1729),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1642),
.A2(n_1561),
.B1(n_896),
.B2(n_1205),
.Y(n_1885)
);

AOI221xp5_ASAP7_75t_L g1886 ( 
.A1(n_1691),
.A2(n_1158),
.B1(n_1444),
.B2(n_762),
.C(n_720),
.Y(n_1886)
);

AOI21xp33_ASAP7_75t_L g1887 ( 
.A1(n_1610),
.A2(n_1439),
.B(n_1419),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1713),
.B(n_1608),
.Y(n_1888)
);

INVx4_ASAP7_75t_L g1889 ( 
.A(n_1761),
.Y(n_1889)
);

OAI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1686),
.A2(n_1576),
.B1(n_1382),
.B2(n_1439),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1700),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1603),
.A2(n_1561),
.B1(n_896),
.B2(n_1205),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1603),
.A2(n_896),
.B1(n_1695),
.B2(n_720),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1713),
.B(n_1608),
.Y(n_1894)
);

AOI221xp5_ASAP7_75t_L g1895 ( 
.A1(n_1691),
.A2(n_1158),
.B1(n_1444),
.B2(n_762),
.C(n_720),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1610),
.B(n_1439),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_L g1897 ( 
.A1(n_1603),
.A2(n_1561),
.B1(n_896),
.B2(n_1205),
.Y(n_1897)
);

OAI221xp5_ASAP7_75t_L g1898 ( 
.A1(n_1695),
.A2(n_720),
.B1(n_709),
.B2(n_1444),
.C(n_896),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1603),
.A2(n_1561),
.B1(n_896),
.B2(n_1205),
.Y(n_1899)
);

AOI222xp33_ASAP7_75t_L g1900 ( 
.A1(n_1603),
.A2(n_930),
.B1(n_980),
.B2(n_674),
.C1(n_1160),
.C2(n_917),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1603),
.A2(n_1561),
.B1(n_896),
.B2(n_1205),
.Y(n_1901)
);

OAI211xp5_ASAP7_75t_SL g1902 ( 
.A1(n_1695),
.A2(n_1450),
.B(n_762),
.C(n_896),
.Y(n_1902)
);

INVx4_ASAP7_75t_SL g1903 ( 
.A(n_1635),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1722),
.B(n_1715),
.Y(n_1904)
);

OAI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1603),
.A2(n_896),
.B1(n_1695),
.B2(n_720),
.Y(n_1905)
);

INVx4_ASAP7_75t_L g1906 ( 
.A(n_1761),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1722),
.B(n_1715),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1722),
.B(n_1715),
.Y(n_1908)
);

OR2x6_ASAP7_75t_L g1909 ( 
.A(n_1635),
.B(n_1665),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1603),
.A2(n_1561),
.B1(n_896),
.B2(n_1205),
.Y(n_1910)
);

OAI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1603),
.A2(n_896),
.B1(n_1695),
.B2(n_720),
.Y(n_1911)
);

BUFx6f_ASAP7_75t_SL g1912 ( 
.A(n_1629),
.Y(n_1912)
);

NAND3xp33_ASAP7_75t_SL g1913 ( 
.A(n_1695),
.B(n_1205),
.C(n_720),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1622),
.Y(n_1914)
);

O2A1O1Ixp33_ASAP7_75t_L g1915 ( 
.A1(n_1691),
.A2(n_709),
.B(n_720),
.C(n_1450),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1695),
.A2(n_709),
.B1(n_720),
.B2(n_1439),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1681),
.B(n_1694),
.Y(n_1917)
);

BUFx6f_ASAP7_75t_L g1918 ( 
.A(n_1597),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1722),
.B(n_1715),
.Y(n_1919)
);

AOI22xp33_ASAP7_75t_L g1920 ( 
.A1(n_1603),
.A2(n_1561),
.B1(n_896),
.B2(n_1205),
.Y(n_1920)
);

OAI221xp5_ASAP7_75t_L g1921 ( 
.A1(n_1695),
.A2(n_720),
.B1(n_709),
.B2(n_1444),
.C(n_896),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1620),
.B(n_1609),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_SL g1923 ( 
.A(n_1594),
.B(n_1487),
.Y(n_1923)
);

AO31x2_ASAP7_75t_L g1924 ( 
.A1(n_1776),
.A2(n_1753),
.A3(n_1631),
.B(n_1625),
.Y(n_1924)
);

AOI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1596),
.A2(n_1389),
.B(n_1245),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1603),
.A2(n_1561),
.B1(n_896),
.B2(n_1205),
.Y(n_1926)
);

NAND3xp33_ASAP7_75t_L g1927 ( 
.A(n_1686),
.B(n_720),
.C(n_709),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1681),
.B(n_1694),
.Y(n_1928)
);

OAI221xp5_ASAP7_75t_L g1929 ( 
.A1(n_1695),
.A2(n_720),
.B1(n_709),
.B2(n_1444),
.C(n_896),
.Y(n_1929)
);

OAI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1686),
.A2(n_1576),
.B1(n_1382),
.B2(n_1439),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1622),
.Y(n_1931)
);

INVx3_ASAP7_75t_L g1932 ( 
.A(n_1761),
.Y(n_1932)
);

CKINVDCx16_ASAP7_75t_R g1933 ( 
.A(n_1655),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1603),
.A2(n_1561),
.B1(n_896),
.B2(n_1205),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1610),
.B(n_1439),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1681),
.B(n_1694),
.Y(n_1936)
);

AOI211xp5_ASAP7_75t_L g1937 ( 
.A1(n_1610),
.A2(n_709),
.B(n_720),
.C(n_1444),
.Y(n_1937)
);

OAI221xp5_ASAP7_75t_L g1938 ( 
.A1(n_1695),
.A2(n_720),
.B1(n_709),
.B2(n_1444),
.C(n_896),
.Y(n_1938)
);

AOI221xp5_ASAP7_75t_L g1939 ( 
.A1(n_1691),
.A2(n_1158),
.B1(n_1444),
.B2(n_762),
.C(n_720),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1603),
.A2(n_896),
.B1(n_1695),
.B2(n_720),
.Y(n_1940)
);

AOI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1603),
.A2(n_1561),
.B1(n_896),
.B2(n_1205),
.Y(n_1941)
);

OAI211xp5_ASAP7_75t_SL g1942 ( 
.A1(n_1695),
.A2(n_1450),
.B(n_762),
.C(n_896),
.Y(n_1942)
);

INVx3_ASAP7_75t_L g1943 ( 
.A(n_1761),
.Y(n_1943)
);

AO21x2_ASAP7_75t_L g1944 ( 
.A1(n_1631),
.A2(n_1625),
.B(n_1753),
.Y(n_1944)
);

OA21x2_ASAP7_75t_L g1945 ( 
.A1(n_1776),
.A2(n_1659),
.B(n_1660),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1731),
.Y(n_1946)
);

AOI222xp33_ASAP7_75t_L g1947 ( 
.A1(n_1603),
.A2(n_930),
.B1(n_980),
.B2(n_674),
.C1(n_1160),
.C2(n_917),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1603),
.A2(n_1561),
.B1(n_896),
.B2(n_1205),
.Y(n_1948)
);

OAI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1603),
.A2(n_896),
.B1(n_1695),
.B2(n_720),
.Y(n_1949)
);

OAI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1686),
.A2(n_1576),
.B1(n_1382),
.B2(n_1439),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1817),
.B(n_1815),
.Y(n_1951)
);

OAI211xp5_ASAP7_75t_L g1952 ( 
.A1(n_1900),
.A2(n_1947),
.B(n_1927),
.C(n_1916),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1860),
.B(n_1866),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1945),
.B(n_1944),
.Y(n_1954)
);

BUFx2_ASAP7_75t_L g1955 ( 
.A(n_1884),
.Y(n_1955)
);

INVxp67_ASAP7_75t_L g1956 ( 
.A(n_1853),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1882),
.Y(n_1957)
);

INVx1_ASAP7_75t_SL g1958 ( 
.A(n_1800),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1904),
.B(n_1907),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1888),
.B(n_1894),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1884),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1823),
.Y(n_1962)
);

INVx3_ASAP7_75t_L g1963 ( 
.A(n_1842),
.Y(n_1963)
);

BUFx2_ASAP7_75t_L g1964 ( 
.A(n_1876),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1813),
.B(n_1822),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1808),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1799),
.B(n_1821),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1808),
.Y(n_1968)
);

INVx3_ASAP7_75t_L g1969 ( 
.A(n_1842),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1804),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1820),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1914),
.Y(n_1972)
);

BUFx6f_ASAP7_75t_L g1973 ( 
.A(n_1918),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1821),
.B(n_1931),
.Y(n_1974)
);

AOI21xp5_ASAP7_75t_L g1975 ( 
.A1(n_1925),
.A2(n_1945),
.B(n_1944),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1908),
.B(n_1919),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1856),
.B(n_1880),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1880),
.B(n_1859),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1924),
.B(n_1945),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1872),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1878),
.B(n_1802),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1832),
.B(n_1858),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1849),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1842),
.B(n_1924),
.Y(n_1984)
);

OR2x2_ASAP7_75t_L g1985 ( 
.A(n_1924),
.B(n_1872),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1873),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1829),
.Y(n_1987)
);

BUFx3_ASAP7_75t_L g1988 ( 
.A(n_1818),
.Y(n_1988)
);

AND2x4_ASAP7_75t_L g1989 ( 
.A(n_1909),
.B(n_1903),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1924),
.B(n_1837),
.Y(n_1990)
);

HB1xp67_ASAP7_75t_L g1991 ( 
.A(n_1861),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1832),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1843),
.B(n_1834),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1837),
.B(n_1883),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1837),
.B(n_1883),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1861),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1867),
.B(n_1881),
.Y(n_1997)
);

OA21x2_ASAP7_75t_L g1998 ( 
.A1(n_1877),
.A2(n_1790),
.B(n_1828),
.Y(n_1998)
);

HB1xp67_ASAP7_75t_L g1999 ( 
.A(n_1879),
.Y(n_1999)
);

OR2x2_ASAP7_75t_L g2000 ( 
.A(n_1807),
.B(n_1946),
.Y(n_2000)
);

INVxp67_ASAP7_75t_L g2001 ( 
.A(n_1801),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1917),
.B(n_1928),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1852),
.Y(n_2003)
);

OR2x6_ASAP7_75t_L g2004 ( 
.A(n_1818),
.B(n_1854),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1881),
.B(n_1865),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1792),
.Y(n_2006)
);

AOI22xp33_ASAP7_75t_SL g2007 ( 
.A1(n_1893),
.A2(n_1911),
.B1(n_1905),
.B2(n_1940),
.Y(n_2007)
);

INVxp67_ASAP7_75t_SL g2008 ( 
.A(n_1841),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1847),
.B(n_1845),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1834),
.B(n_1805),
.Y(n_2010)
);

INVx2_ASAP7_75t_SL g2011 ( 
.A(n_1818),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1805),
.B(n_1845),
.Y(n_2012)
);

AOI22xp33_ASAP7_75t_L g2013 ( 
.A1(n_1949),
.A2(n_1913),
.B1(n_1929),
.B2(n_1921),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1836),
.B(n_1857),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1936),
.B(n_1935),
.Y(n_2015)
);

BUFx2_ASAP7_75t_L g2016 ( 
.A(n_1869),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1836),
.B(n_1835),
.Y(n_2017)
);

AND2x4_ASAP7_75t_L g2018 ( 
.A(n_1903),
.B(n_1838),
.Y(n_2018)
);

INVx2_ASAP7_75t_SL g2019 ( 
.A(n_1869),
.Y(n_2019)
);

INVx1_ASAP7_75t_SL g2020 ( 
.A(n_1891),
.Y(n_2020)
);

AOI221xp5_ASAP7_75t_L g2021 ( 
.A1(n_1898),
.A2(n_1938),
.B1(n_1794),
.B2(n_1915),
.C(n_1948),
.Y(n_2021)
);

INVxp67_ASAP7_75t_L g2022 ( 
.A(n_1935),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1835),
.B(n_1863),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1903),
.B(n_1838),
.Y(n_2024)
);

NOR2x1_ASAP7_75t_SL g2025 ( 
.A(n_1851),
.B(n_1896),
.Y(n_2025)
);

BUFx3_ASAP7_75t_L g2026 ( 
.A(n_1816),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1798),
.B(n_1896),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1830),
.Y(n_2028)
);

INVx2_ASAP7_75t_R g2029 ( 
.A(n_1791),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1892),
.A2(n_1899),
.B1(n_1920),
.B2(n_1948),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1871),
.Y(n_2031)
);

HB1xp67_ASAP7_75t_L g2032 ( 
.A(n_1855),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1871),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1798),
.B(n_1812),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1812),
.B(n_1887),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1937),
.B(n_1793),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1862),
.B(n_1870),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1824),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1811),
.B(n_1826),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_1833),
.B(n_1809),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1819),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_1850),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1803),
.B(n_1840),
.Y(n_2043)
);

OR2x2_ASAP7_75t_L g2044 ( 
.A(n_1959),
.B(n_1933),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1962),
.Y(n_2045)
);

NOR2x1_ASAP7_75t_L g2046 ( 
.A(n_2026),
.B(n_1986),
.Y(n_2046)
);

OA21x2_ASAP7_75t_L g2047 ( 
.A1(n_1975),
.A2(n_1814),
.B(n_1885),
.Y(n_2047)
);

INVx2_ASAP7_75t_SL g2048 ( 
.A(n_2037),
.Y(n_2048)
);

AOI221xp5_ASAP7_75t_L g2049 ( 
.A1(n_1952),
.A2(n_1886),
.B1(n_1895),
.B2(n_1939),
.C(n_1902),
.Y(n_2049)
);

HB1xp67_ASAP7_75t_L g2050 ( 
.A(n_1966),
.Y(n_2050)
);

AOI221xp5_ASAP7_75t_L g2051 ( 
.A1(n_1952),
.A2(n_1942),
.B1(n_1950),
.B2(n_1930),
.C(n_1890),
.Y(n_2051)
);

AOI33xp33_ASAP7_75t_L g2052 ( 
.A1(n_2007),
.A2(n_1910),
.A3(n_1941),
.B1(n_1934),
.B2(n_1926),
.B3(n_1920),
.Y(n_2052)
);

AOI22xp33_ASAP7_75t_L g2053 ( 
.A1(n_2007),
.A2(n_1910),
.B1(n_1941),
.B2(n_1934),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1962),
.Y(n_2054)
);

AND4x1_ASAP7_75t_L g2055 ( 
.A(n_2021),
.B(n_1923),
.C(n_1848),
.D(n_1901),
.Y(n_2055)
);

NOR3xp33_ASAP7_75t_L g2056 ( 
.A(n_2021),
.B(n_1796),
.C(n_1890),
.Y(n_2056)
);

INVx4_ASAP7_75t_L g2057 ( 
.A(n_1973),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_1966),
.Y(n_2058)
);

BUFx3_ASAP7_75t_L g2059 ( 
.A(n_2026),
.Y(n_2059)
);

OAI33xp33_ASAP7_75t_L g2060 ( 
.A1(n_2022),
.A2(n_1930),
.A3(n_1950),
.B1(n_1806),
.B2(n_1797),
.B3(n_1825),
.Y(n_2060)
);

AOI221xp5_ASAP7_75t_SL g2061 ( 
.A1(n_2022),
.A2(n_1926),
.B1(n_1892),
.B2(n_1897),
.C(n_1899),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1970),
.Y(n_2062)
);

INVx3_ASAP7_75t_L g2063 ( 
.A(n_2026),
.Y(n_2063)
);

OR2x2_ASAP7_75t_L g2064 ( 
.A(n_1959),
.B(n_1976),
.Y(n_2064)
);

OAI221xp5_ASAP7_75t_L g2065 ( 
.A1(n_2013),
.A2(n_1897),
.B1(n_1901),
.B2(n_1794),
.C(n_1810),
.Y(n_2065)
);

INVxp67_ASAP7_75t_L g2066 ( 
.A(n_1978),
.Y(n_2066)
);

OAI211xp5_ASAP7_75t_L g2067 ( 
.A1(n_2036),
.A2(n_1885),
.B(n_1814),
.C(n_1810),
.Y(n_2067)
);

INVx4_ASAP7_75t_L g2068 ( 
.A(n_1973),
.Y(n_2068)
);

AOI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_2030),
.A2(n_1831),
.B1(n_1825),
.B2(n_1912),
.Y(n_2069)
);

OAI221xp5_ASAP7_75t_L g2070 ( 
.A1(n_2036),
.A2(n_1906),
.B1(n_1889),
.B2(n_1839),
.C(n_1943),
.Y(n_2070)
);

INVxp67_ASAP7_75t_SL g2071 ( 
.A(n_1980),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1972),
.Y(n_2072)
);

OAI221xp5_ASAP7_75t_L g2073 ( 
.A1(n_2027),
.A2(n_1906),
.B1(n_1889),
.B2(n_1943),
.C(n_1795),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1951),
.B(n_2037),
.Y(n_2074)
);

AOI21xp5_ASAP7_75t_L g2075 ( 
.A1(n_2027),
.A2(n_1827),
.B(n_1922),
.Y(n_2075)
);

AOI22xp33_ASAP7_75t_L g2076 ( 
.A1(n_2041),
.A2(n_1912),
.B1(n_1922),
.B2(n_1844),
.Y(n_2076)
);

OAI211xp5_ASAP7_75t_SL g2077 ( 
.A1(n_2015),
.A2(n_1795),
.B(n_1932),
.C(n_1864),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_SL g2078 ( 
.A(n_1958),
.B(n_1875),
.Y(n_2078)
);

AOI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_2041),
.A2(n_1932),
.B1(n_1864),
.B2(n_1868),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_L g2080 ( 
.A(n_2015),
.B(n_1874),
.Y(n_2080)
);

AOI221xp5_ASAP7_75t_L g2081 ( 
.A1(n_2038),
.A2(n_1846),
.B1(n_1874),
.B2(n_1918),
.C(n_2028),
.Y(n_2081)
);

AOI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_2028),
.A2(n_1846),
.B1(n_2038),
.B2(n_2014),
.Y(n_2082)
);

OAI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_2028),
.A2(n_2009),
.B1(n_2034),
.B2(n_2043),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1951),
.B(n_2039),
.Y(n_2084)
);

AOI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_2014),
.A2(n_2043),
.B1(n_2008),
.B2(n_1967),
.Y(n_2085)
);

NAND2x1p5_ASAP7_75t_L g2086 ( 
.A(n_1989),
.B(n_2016),
.Y(n_2086)
);

NAND3xp33_ASAP7_75t_SL g2087 ( 
.A(n_2043),
.B(n_2035),
.C(n_2009),
.Y(n_2087)
);

OAI22xp5_ASAP7_75t_L g2088 ( 
.A1(n_2034),
.A2(n_1982),
.B1(n_2040),
.B2(n_2035),
.Y(n_2088)
);

INVxp67_ASAP7_75t_SL g2089 ( 
.A(n_1980),
.Y(n_2089)
);

OR2x6_ASAP7_75t_L g2090 ( 
.A(n_2004),
.B(n_1989),
.Y(n_2090)
);

INVx5_ASAP7_75t_SL g2091 ( 
.A(n_2004),
.Y(n_2091)
);

AOI211x1_ASAP7_75t_L g2092 ( 
.A1(n_2002),
.A2(n_1981),
.B(n_1982),
.C(n_1987),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_1957),
.Y(n_2093)
);

NAND4xp25_ASAP7_75t_L g2094 ( 
.A(n_2002),
.B(n_2001),
.C(n_1981),
.D(n_1967),
.Y(n_2094)
);

AOI221xp5_ASAP7_75t_L g2095 ( 
.A1(n_2001),
.A2(n_2008),
.B1(n_1993),
.B2(n_2012),
.C(n_1999),
.Y(n_2095)
);

AOI322xp5_ASAP7_75t_L g2096 ( 
.A1(n_1993),
.A2(n_2012),
.A3(n_2010),
.B1(n_1965),
.B2(n_1997),
.C1(n_2005),
.C2(n_1999),
.Y(n_2096)
);

NAND3xp33_ASAP7_75t_L g2097 ( 
.A(n_1998),
.B(n_1975),
.C(n_1986),
.Y(n_2097)
);

AOI221xp5_ASAP7_75t_L g2098 ( 
.A1(n_2006),
.A2(n_2010),
.B1(n_1997),
.B2(n_2005),
.C(n_1987),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_1953),
.B(n_1978),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2003),
.B(n_2000),
.Y(n_2100)
);

HB1xp67_ASAP7_75t_L g2101 ( 
.A(n_1957),
.Y(n_2101)
);

NOR2xp33_ASAP7_75t_R g2102 ( 
.A(n_2019),
.B(n_2016),
.Y(n_2102)
);

AOI22xp33_ASAP7_75t_SL g2103 ( 
.A1(n_2025),
.A2(n_1998),
.B1(n_2005),
.B2(n_1997),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2003),
.B(n_2000),
.Y(n_2104)
);

OAI22xp5_ASAP7_75t_L g2105 ( 
.A1(n_2040),
.A2(n_2020),
.B1(n_1998),
.B2(n_2032),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1971),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1971),
.Y(n_2107)
);

AOI221xp5_ASAP7_75t_L g2108 ( 
.A1(n_2006),
.A2(n_1965),
.B1(n_1974),
.B2(n_2042),
.C(n_2032),
.Y(n_2108)
);

AOI22xp33_ASAP7_75t_L g2109 ( 
.A1(n_2006),
.A2(n_1998),
.B1(n_2029),
.B2(n_1974),
.Y(n_2109)
);

AOI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_1998),
.A2(n_2029),
.B1(n_2023),
.B2(n_2042),
.Y(n_2110)
);

AND2x4_ASAP7_75t_SL g2111 ( 
.A(n_1989),
.B(n_1960),
.Y(n_2111)
);

OAI31xp33_ASAP7_75t_L g2112 ( 
.A1(n_1988),
.A2(n_2023),
.A3(n_2017),
.B(n_2025),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2093),
.Y(n_2113)
);

OR2x2_ASAP7_75t_L g2114 ( 
.A(n_2066),
.B(n_1979),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2106),
.B(n_1954),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_2066),
.B(n_1979),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2099),
.B(n_1983),
.Y(n_2117)
);

AND2x4_ASAP7_75t_SL g2118 ( 
.A(n_2090),
.B(n_2018),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_2101),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2071),
.B(n_1983),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2101),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2107),
.Y(n_2122)
);

AND2x4_ASAP7_75t_L g2123 ( 
.A(n_2090),
.B(n_1961),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2071),
.B(n_1992),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2074),
.B(n_1984),
.Y(n_2125)
);

NAND2x1p5_ASAP7_75t_L g2126 ( 
.A(n_2047),
.B(n_1963),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2045),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2054),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2090),
.B(n_1984),
.Y(n_2129)
);

AND2x4_ASAP7_75t_L g2130 ( 
.A(n_2057),
.B(n_1961),
.Y(n_2130)
);

INVx1_ASAP7_75t_SL g2131 ( 
.A(n_2046),
.Y(n_2131)
);

OR2x2_ASAP7_75t_L g2132 ( 
.A(n_2097),
.B(n_1985),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_SL g2133 ( 
.A(n_2103),
.B(n_2112),
.Y(n_2133)
);

HB1xp67_ASAP7_75t_L g2134 ( 
.A(n_2050),
.Y(n_2134)
);

INVx3_ASAP7_75t_L g2135 ( 
.A(n_2057),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2089),
.B(n_1992),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2062),
.Y(n_2137)
);

AND2x4_ASAP7_75t_L g2138 ( 
.A(n_2068),
.B(n_1961),
.Y(n_2138)
);

BUFx2_ASAP7_75t_L g2139 ( 
.A(n_2102),
.Y(n_2139)
);

AND2x4_ASAP7_75t_SL g2140 ( 
.A(n_2068),
.B(n_2018),
.Y(n_2140)
);

OR2x2_ASAP7_75t_L g2141 ( 
.A(n_2050),
.B(n_2058),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2091),
.B(n_1969),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2072),
.Y(n_2143)
);

INVxp33_ASAP7_75t_L g2144 ( 
.A(n_2102),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2109),
.B(n_1990),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2089),
.B(n_2105),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2109),
.B(n_1990),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2092),
.B(n_1953),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2048),
.B(n_1994),
.Y(n_2149)
);

OR2x2_ASAP7_75t_L g2150 ( 
.A(n_2058),
.B(n_1985),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2110),
.B(n_1995),
.Y(n_2151)
);

OR2x2_ASAP7_75t_L g2152 ( 
.A(n_2064),
.B(n_1991),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2110),
.B(n_1995),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2100),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2084),
.B(n_1996),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2047),
.B(n_1996),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_2104),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2047),
.B(n_1991),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2088),
.B(n_1964),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2086),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2103),
.B(n_1957),
.Y(n_2161)
);

BUFx2_ASAP7_75t_L g2162 ( 
.A(n_2139),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2161),
.B(n_2029),
.Y(n_2163)
);

NOR2x1p5_ASAP7_75t_L g2164 ( 
.A(n_2159),
.B(n_2087),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2161),
.B(n_1964),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_2119),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2127),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2119),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2161),
.B(n_2086),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2161),
.B(n_1955),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_2119),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2127),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2127),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2127),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2159),
.B(n_2080),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2143),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2143),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2154),
.B(n_2080),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_2129),
.B(n_1955),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2129),
.B(n_2063),
.Y(n_2180)
);

AOI32xp33_ASAP7_75t_L g2181 ( 
.A1(n_2151),
.A2(n_2056),
.A3(n_2049),
.B1(n_2095),
.B2(n_2051),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2119),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2143),
.Y(n_2183)
);

BUFx2_ASAP7_75t_L g2184 ( 
.A(n_2139),
.Y(n_2184)
);

AND2x2_ASAP7_75t_SL g2185 ( 
.A(n_2132),
.B(n_2056),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2143),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2129),
.B(n_2063),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2115),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2154),
.B(n_2108),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2115),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2154),
.B(n_2094),
.Y(n_2191)
);

OR2x2_ASAP7_75t_L g2192 ( 
.A(n_2114),
.B(n_1968),
.Y(n_2192)
);

OR2x2_ASAP7_75t_L g2193 ( 
.A(n_2114),
.B(n_1968),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2122),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2115),
.Y(n_2195)
);

AND2x2_ASAP7_75t_SL g2196 ( 
.A(n_2132),
.B(n_2055),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2122),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2154),
.B(n_2098),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2129),
.B(n_2111),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2115),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2157),
.B(n_2085),
.Y(n_2201)
);

OAI33xp33_ASAP7_75t_L g2202 ( 
.A1(n_2133),
.A2(n_2083),
.A3(n_2044),
.B1(n_1956),
.B2(n_2031),
.B3(n_2033),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2156),
.Y(n_2203)
);

NOR2xp33_ASAP7_75t_L g2204 ( 
.A(n_2148),
.B(n_2070),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_2149),
.B(n_2059),
.Y(n_2205)
);

INVx1_ASAP7_75t_SL g2206 ( 
.A(n_2131),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2122),
.Y(n_2207)
);

AND2x4_ASAP7_75t_L g2208 ( 
.A(n_2123),
.B(n_1989),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2113),
.Y(n_2209)
);

OR2x2_ASAP7_75t_L g2210 ( 
.A(n_2114),
.B(n_1977),
.Y(n_2210)
);

OR2x2_ASAP7_75t_L g2211 ( 
.A(n_2114),
.B(n_1977),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2128),
.Y(n_2212)
);

INVxp67_ASAP7_75t_L g2213 ( 
.A(n_2185),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2188),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2199),
.B(n_2139),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2199),
.B(n_2169),
.Y(n_2216)
);

OR2x2_ASAP7_75t_L g2217 ( 
.A(n_2201),
.B(n_2191),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2185),
.B(n_2148),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2185),
.B(n_2204),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2185),
.B(n_2146),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2204),
.B(n_2146),
.Y(n_2221)
);

NAND3xp33_ASAP7_75t_L g2222 ( 
.A(n_2181),
.B(n_2133),
.C(n_2096),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2212),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2212),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2175),
.B(n_2157),
.Y(n_2225)
);

NOR2x1_ASAP7_75t_L g2226 ( 
.A(n_2164),
.B(n_2206),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_SL g2227 ( 
.A(n_2196),
.B(n_2131),
.Y(n_2227)
);

OR2x2_ASAP7_75t_L g2228 ( 
.A(n_2201),
.B(n_2191),
.Y(n_2228)
);

AND2x4_ASAP7_75t_L g2229 ( 
.A(n_2162),
.B(n_2118),
.Y(n_2229)
);

OR2x2_ASAP7_75t_L g2230 ( 
.A(n_2178),
.B(n_2117),
.Y(n_2230)
);

OR2x2_ASAP7_75t_L g2231 ( 
.A(n_2178),
.B(n_2117),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2175),
.B(n_2157),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2194),
.Y(n_2233)
);

NOR2xp33_ASAP7_75t_L g2234 ( 
.A(n_2202),
.B(n_2078),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2194),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2199),
.B(n_2125),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2194),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2164),
.B(n_2157),
.Y(n_2238)
);

OR2x2_ASAP7_75t_L g2239 ( 
.A(n_2189),
.B(n_2151),
.Y(n_2239)
);

INVx2_ASAP7_75t_SL g2240 ( 
.A(n_2162),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2207),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2207),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2188),
.Y(n_2243)
);

NOR2xp67_ASAP7_75t_L g2244 ( 
.A(n_2169),
.B(n_2160),
.Y(n_2244)
);

NAND4xp25_ASAP7_75t_SL g2245 ( 
.A(n_2181),
.B(n_2053),
.C(n_2052),
.D(n_2061),
.Y(n_2245)
);

NOR3xp33_ASAP7_75t_SL g2246 ( 
.A(n_2202),
.B(n_2073),
.C(n_2060),
.Y(n_2246)
);

OR2x2_ASAP7_75t_L g2247 ( 
.A(n_2189),
.B(n_2151),
.Y(n_2247)
);

OR2x2_ASAP7_75t_L g2248 ( 
.A(n_2198),
.B(n_2151),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_2169),
.B(n_2160),
.Y(n_2249)
);

OAI33xp33_ASAP7_75t_L g2250 ( 
.A1(n_2198),
.A2(n_2132),
.A3(n_2124),
.B1(n_2136),
.B2(n_2141),
.B3(n_2116),
.Y(n_2250)
);

INVx2_ASAP7_75t_SL g2251 ( 
.A(n_2162),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2207),
.Y(n_2252)
);

BUFx2_ASAP7_75t_L g2253 ( 
.A(n_2184),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2197),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2197),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2209),
.Y(n_2256)
);

AOI32xp33_ASAP7_75t_L g2257 ( 
.A1(n_2163),
.A2(n_2153),
.A3(n_2145),
.B1(n_2147),
.B2(n_2144),
.Y(n_2257)
);

NAND2x1p5_ASAP7_75t_L g2258 ( 
.A(n_2196),
.B(n_2135),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2209),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2209),
.Y(n_2260)
);

AOI22xp33_ASAP7_75t_L g2261 ( 
.A1(n_2196),
.A2(n_2053),
.B1(n_2065),
.B2(n_2069),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2196),
.B(n_2155),
.Y(n_2262)
);

NAND2xp33_ASAP7_75t_R g2263 ( 
.A(n_2184),
.B(n_2153),
.Y(n_2263)
);

AND2x4_ASAP7_75t_L g2264 ( 
.A(n_2240),
.B(n_2184),
.Y(n_2264)
);

HB1xp67_ASAP7_75t_L g2265 ( 
.A(n_2240),
.Y(n_2265)
);

OR2x2_ASAP7_75t_L g2266 ( 
.A(n_2230),
.B(n_2210),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2253),
.Y(n_2267)
);

XNOR2xp5_ASAP7_75t_L g2268 ( 
.A(n_2222),
.B(n_2082),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2233),
.Y(n_2269)
);

HB1xp67_ASAP7_75t_L g2270 ( 
.A(n_2251),
.Y(n_2270)
);

O2A1O1Ixp33_ASAP7_75t_L g2271 ( 
.A1(n_2227),
.A2(n_2206),
.B(n_2163),
.C(n_2132),
.Y(n_2271)
);

AOI32xp33_ASAP7_75t_L g2272 ( 
.A1(n_2226),
.A2(n_2234),
.A3(n_2219),
.B1(n_2227),
.B2(n_2221),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2235),
.Y(n_2273)
);

OAI322xp33_ASAP7_75t_L g2274 ( 
.A1(n_2213),
.A2(n_2211),
.A3(n_2210),
.B1(n_2163),
.B2(n_2116),
.C1(n_2165),
.C2(n_2150),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2234),
.B(n_2165),
.Y(n_2275)
);

OAI22xp5_ASAP7_75t_L g2276 ( 
.A1(n_2261),
.A2(n_2144),
.B1(n_2069),
.B2(n_2165),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2237),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2241),
.Y(n_2278)
);

NOR2xp33_ASAP7_75t_L g2279 ( 
.A(n_2245),
.B(n_2208),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2242),
.Y(n_2280)
);

NAND2x1_ASAP7_75t_SL g2281 ( 
.A(n_2229),
.B(n_2170),
.Y(n_2281)
);

AOI22xp33_ASAP7_75t_L g2282 ( 
.A1(n_2261),
.A2(n_2153),
.B1(n_2145),
.B2(n_2147),
.Y(n_2282)
);

OAI221xp5_ASAP7_75t_L g2283 ( 
.A1(n_2213),
.A2(n_2067),
.B1(n_2210),
.B2(n_2211),
.C(n_2153),
.Y(n_2283)
);

AOI221xp5_ASAP7_75t_L g2284 ( 
.A1(n_2250),
.A2(n_2145),
.B1(n_2147),
.B2(n_2158),
.C(n_2203),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2258),
.B(n_2208),
.Y(n_2285)
);

AOI21xp5_ASAP7_75t_L g2286 ( 
.A1(n_2220),
.A2(n_2075),
.B(n_2145),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2252),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2223),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2224),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2251),
.Y(n_2290)
);

INVx1_ASAP7_75t_SL g2291 ( 
.A(n_2215),
.Y(n_2291)
);

NOR2xp33_ASAP7_75t_L g2292 ( 
.A(n_2218),
.B(n_2208),
.Y(n_2292)
);

OAI21xp33_ASAP7_75t_L g2293 ( 
.A1(n_2246),
.A2(n_2147),
.B(n_2211),
.Y(n_2293)
);

AOI21xp33_ASAP7_75t_L g2294 ( 
.A1(n_2263),
.A2(n_2158),
.B(n_2011),
.Y(n_2294)
);

OAI221xp5_ASAP7_75t_L g2295 ( 
.A1(n_2257),
.A2(n_2076),
.B1(n_2160),
.B2(n_2081),
.C(n_2116),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2246),
.B(n_2170),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2217),
.B(n_2170),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2258),
.B(n_2216),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2254),
.Y(n_2299)
);

OAI32xp33_ASAP7_75t_L g2300 ( 
.A1(n_2263),
.A2(n_2158),
.A3(n_2203),
.B1(n_2126),
.B2(n_2116),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2228),
.B(n_2125),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2238),
.B(n_2125),
.Y(n_2302)
);

INVxp67_ASAP7_75t_L g2303 ( 
.A(n_2248),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2229),
.B(n_2208),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2298),
.B(n_2229),
.Y(n_2305)
);

AOI22xp5_ASAP7_75t_L g2306 ( 
.A1(n_2293),
.A2(n_2250),
.B1(n_2262),
.B2(n_2239),
.Y(n_2306)
);

NAND3xp33_ASAP7_75t_SL g2307 ( 
.A(n_2272),
.B(n_2247),
.C(n_2231),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2269),
.Y(n_2308)
);

AOI22xp5_ASAP7_75t_L g2309 ( 
.A1(n_2296),
.A2(n_2244),
.B1(n_2225),
.B2(n_2232),
.Y(n_2309)
);

O2A1O1Ixp33_ASAP7_75t_SL g2310 ( 
.A1(n_2268),
.A2(n_2134),
.B(n_2077),
.C(n_2019),
.Y(n_2310)
);

OAI32xp33_ASAP7_75t_L g2311 ( 
.A1(n_2275),
.A2(n_2203),
.A3(n_2249),
.B1(n_2158),
.B2(n_2126),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2273),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2277),
.Y(n_2313)
);

OR2x2_ASAP7_75t_L g2314 ( 
.A(n_2297),
.B(n_2236),
.Y(n_2314)
);

OR2x2_ASAP7_75t_L g2315 ( 
.A(n_2291),
.B(n_2249),
.Y(n_2315)
);

XNOR2xp5_ASAP7_75t_L g2316 ( 
.A(n_2268),
.B(n_2076),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2278),
.Y(n_2317)
);

NAND2xp33_ASAP7_75t_SL g2318 ( 
.A(n_2281),
.B(n_2160),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2280),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2287),
.Y(n_2320)
);

O2A1O1Ixp5_ASAP7_75t_SL g2321 ( 
.A1(n_2267),
.A2(n_2260),
.B(n_2259),
.C(n_2256),
.Y(n_2321)
);

AOI32xp33_ASAP7_75t_L g2322 ( 
.A1(n_2279),
.A2(n_2187),
.A3(n_2180),
.B1(n_2205),
.B2(n_2179),
.Y(n_2322)
);

OR2x2_ASAP7_75t_L g2323 ( 
.A(n_2303),
.B(n_2255),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_L g2324 ( 
.A(n_2279),
.B(n_2208),
.Y(n_2324)
);

INVx1_ASAP7_75t_SL g2325 ( 
.A(n_2264),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2288),
.Y(n_2326)
);

OAI22xp33_ASAP7_75t_SL g2327 ( 
.A1(n_2283),
.A2(n_2203),
.B1(n_2214),
.B2(n_2243),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2289),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2282),
.B(n_2214),
.Y(n_2329)
);

XNOR2x2_ASAP7_75t_L g2330 ( 
.A(n_2276),
.B(n_2141),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2282),
.B(n_2243),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2299),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2265),
.Y(n_2333)
);

AOI322xp5_ASAP7_75t_L g2334 ( 
.A1(n_2284),
.A2(n_2179),
.A3(n_2195),
.B1(n_2190),
.B2(n_2188),
.C1(n_2200),
.C2(n_2156),
.Y(n_2334)
);

AOI32xp33_ASAP7_75t_L g2335 ( 
.A1(n_2298),
.A2(n_2180),
.A3(n_2187),
.B1(n_2205),
.B2(n_2179),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2325),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2305),
.B(n_2304),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2325),
.Y(n_2338)
);

AOI221xp5_ASAP7_75t_L g2339 ( 
.A1(n_2307),
.A2(n_2271),
.B1(n_2300),
.B2(n_2274),
.C(n_2294),
.Y(n_2339)
);

OAI21xp33_ASAP7_75t_L g2340 ( 
.A1(n_2306),
.A2(n_2281),
.B(n_2292),
.Y(n_2340)
);

INVxp67_ASAP7_75t_L g2341 ( 
.A(n_2333),
.Y(n_2341)
);

OAI21xp5_ASAP7_75t_L g2342 ( 
.A1(n_2321),
.A2(n_2286),
.B(n_2270),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2308),
.Y(n_2343)
);

AOI22xp5_ASAP7_75t_L g2344 ( 
.A1(n_2324),
.A2(n_2292),
.B1(n_2285),
.B2(n_2304),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_2316),
.B(n_2264),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2326),
.B(n_2290),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2328),
.B(n_2290),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2312),
.Y(n_2348)
);

XOR2x2_ASAP7_75t_L g2349 ( 
.A(n_2330),
.B(n_2295),
.Y(n_2349)
);

NOR3x1_ASAP7_75t_L g2350 ( 
.A(n_2329),
.B(n_2301),
.C(n_2302),
.Y(n_2350)
);

AOI21xp33_ASAP7_75t_L g2351 ( 
.A1(n_2327),
.A2(n_2331),
.B(n_2329),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2313),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2317),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2319),
.Y(n_2354)
);

NAND2xp33_ASAP7_75t_SL g2355 ( 
.A(n_2331),
.B(n_2264),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2320),
.Y(n_2356)
);

NAND2xp33_ASAP7_75t_SL g2357 ( 
.A(n_2323),
.B(n_2285),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2332),
.Y(n_2358)
);

OR3x1_ASAP7_75t_L g2359 ( 
.A(n_2311),
.B(n_2177),
.C(n_2176),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2322),
.B(n_2266),
.Y(n_2360)
);

NOR2xp33_ASAP7_75t_L g2361 ( 
.A(n_2345),
.B(n_2314),
.Y(n_2361)
);

O2A1O1Ixp33_ASAP7_75t_SL g2362 ( 
.A1(n_2342),
.A2(n_2334),
.B(n_2315),
.C(n_2309),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_2337),
.B(n_2266),
.Y(n_2363)
);

NOR2x1_ASAP7_75t_L g2364 ( 
.A(n_2345),
.B(n_2318),
.Y(n_2364)
);

NAND3xp33_ASAP7_75t_L g2365 ( 
.A(n_2355),
.B(n_2335),
.C(n_2310),
.Y(n_2365)
);

NOR2xp33_ASAP7_75t_L g2366 ( 
.A(n_2341),
.B(n_2208),
.Y(n_2366)
);

INVx1_ASAP7_75t_SL g2367 ( 
.A(n_2357),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2336),
.B(n_2180),
.Y(n_2368)
);

NOR3xp33_ASAP7_75t_L g2369 ( 
.A(n_2351),
.B(n_2011),
.C(n_2135),
.Y(n_2369)
);

AOI22xp5_ASAP7_75t_L g2370 ( 
.A1(n_2349),
.A2(n_2140),
.B1(n_2118),
.B2(n_2011),
.Y(n_2370)
);

AOI22xp5_ASAP7_75t_L g2371 ( 
.A1(n_2340),
.A2(n_2140),
.B1(n_2118),
.B2(n_2187),
.Y(n_2371)
);

NOR2xp67_ASAP7_75t_SL g2372 ( 
.A(n_2338),
.B(n_1988),
.Y(n_2372)
);

OAI21xp5_ASAP7_75t_L g2373 ( 
.A1(n_2339),
.A2(n_1956),
.B(n_2135),
.Y(n_2373)
);

NOR3x1_ASAP7_75t_L g2374 ( 
.A(n_2346),
.B(n_2347),
.C(n_2360),
.Y(n_2374)
);

NOR3xp33_ASAP7_75t_L g2375 ( 
.A(n_2355),
.B(n_2156),
.C(n_2135),
.Y(n_2375)
);

AOI221x1_ASAP7_75t_L g2376 ( 
.A1(n_2369),
.A2(n_2357),
.B1(n_2358),
.B2(n_2353),
.C(n_2356),
.Y(n_2376)
);

NAND4xp25_ASAP7_75t_L g2377 ( 
.A(n_2361),
.B(n_2350),
.C(n_2341),
.D(n_2344),
.Y(n_2377)
);

AOI221xp5_ASAP7_75t_L g2378 ( 
.A1(n_2362),
.A2(n_2354),
.B1(n_2352),
.B2(n_2348),
.C(n_2343),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2367),
.B(n_2359),
.Y(n_2379)
);

NAND3xp33_ASAP7_75t_L g2380 ( 
.A(n_2364),
.B(n_2365),
.C(n_2375),
.Y(n_2380)
);

AOI221x1_ASAP7_75t_L g2381 ( 
.A1(n_2375),
.A2(n_2166),
.B1(n_2168),
.B2(n_2171),
.C(n_2182),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2363),
.B(n_2366),
.Y(n_2382)
);

OAI221xp5_ASAP7_75t_L g2383 ( 
.A1(n_2371),
.A2(n_1988),
.B1(n_2135),
.B2(n_2079),
.C(n_2188),
.Y(n_2383)
);

AOI322xp5_ASAP7_75t_L g2384 ( 
.A1(n_2370),
.A2(n_2156),
.A3(n_2195),
.B1(n_2190),
.B2(n_2200),
.C1(n_2134),
.C2(n_2205),
.Y(n_2384)
);

OAI21xp33_ASAP7_75t_L g2385 ( 
.A1(n_2368),
.A2(n_2140),
.B(n_2118),
.Y(n_2385)
);

AOI221xp5_ASAP7_75t_L g2386 ( 
.A1(n_2373),
.A2(n_2171),
.B1(n_2166),
.B2(n_2168),
.C(n_2182),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_L g2387 ( 
.A(n_2372),
.B(n_2192),
.Y(n_2387)
);

NOR3xp33_ASAP7_75t_SL g2388 ( 
.A(n_2377),
.B(n_2374),
.C(n_2120),
.Y(n_2388)
);

AOI222xp33_ASAP7_75t_L g2389 ( 
.A1(n_2380),
.A2(n_2124),
.B1(n_2136),
.B2(n_2171),
.C1(n_2166),
.C2(n_2168),
.Y(n_2389)
);

AOI21xp33_ASAP7_75t_SL g2390 ( 
.A1(n_2379),
.A2(n_2182),
.B(n_2168),
.Y(n_2390)
);

AOI22xp33_ASAP7_75t_L g2391 ( 
.A1(n_2378),
.A2(n_2004),
.B1(n_2024),
.B2(n_2018),
.Y(n_2391)
);

OAI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_2376),
.A2(n_2166),
.B(n_2171),
.Y(n_2392)
);

NAND2xp33_ASAP7_75t_SL g2393 ( 
.A(n_2382),
.B(n_2135),
.Y(n_2393)
);

OAI31xp33_ASAP7_75t_L g2394 ( 
.A1(n_2383),
.A2(n_2140),
.A3(n_2126),
.B(n_2182),
.Y(n_2394)
);

OAI211xp5_ASAP7_75t_SL g2395 ( 
.A1(n_2388),
.A2(n_2384),
.B(n_2385),
.C(n_2387),
.Y(n_2395)
);

INVx3_ASAP7_75t_L g2396 ( 
.A(n_2393),
.Y(n_2396)
);

AOI22xp5_ASAP7_75t_L g2397 ( 
.A1(n_2391),
.A2(n_2386),
.B1(n_2130),
.B2(n_2138),
.Y(n_2397)
);

NOR2xp67_ASAP7_75t_L g2398 ( 
.A(n_2390),
.B(n_2381),
.Y(n_2398)
);

NOR3xp33_ASAP7_75t_L g2399 ( 
.A(n_2392),
.B(n_2120),
.C(n_2142),
.Y(n_2399)
);

INVxp67_ASAP7_75t_SL g2400 ( 
.A(n_2389),
.Y(n_2400)
);

OR2x2_ASAP7_75t_L g2401 ( 
.A(n_2394),
.B(n_2190),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2388),
.B(n_2190),
.Y(n_2402)
);

AOI22xp5_ASAP7_75t_L g2403 ( 
.A1(n_2395),
.A2(n_2130),
.B1(n_2138),
.B2(n_2200),
.Y(n_2403)
);

AOI22xp5_ASAP7_75t_L g2404 ( 
.A1(n_2400),
.A2(n_2130),
.B1(n_2138),
.B2(n_2200),
.Y(n_2404)
);

NAND3xp33_ASAP7_75t_SL g2405 ( 
.A(n_2399),
.B(n_2079),
.C(n_2141),
.Y(n_2405)
);

OAI322xp33_ASAP7_75t_L g2406 ( 
.A1(n_2402),
.A2(n_2192),
.A3(n_2193),
.B1(n_2141),
.B2(n_2195),
.C1(n_2177),
.C2(n_2176),
.Y(n_2406)
);

NOR3x1_ASAP7_75t_L g2407 ( 
.A(n_2401),
.B(n_2192),
.C(n_2193),
.Y(n_2407)
);

NAND3xp33_ASAP7_75t_SL g2408 ( 
.A(n_2397),
.B(n_2126),
.C(n_2152),
.Y(n_2408)
);

NAND3xp33_ASAP7_75t_L g2409 ( 
.A(n_2396),
.B(n_2176),
.C(n_2174),
.Y(n_2409)
);

INVx3_ASAP7_75t_L g2410 ( 
.A(n_2407),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2403),
.B(n_2398),
.Y(n_2411)
);

HB1xp67_ASAP7_75t_L g2412 ( 
.A(n_2409),
.Y(n_2412)
);

OR3x2_ASAP7_75t_L g2413 ( 
.A(n_2408),
.B(n_2152),
.C(n_2150),
.Y(n_2413)
);

OAI22xp33_ASAP7_75t_L g2414 ( 
.A1(n_2410),
.A2(n_2404),
.B1(n_2405),
.B2(n_2406),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2411),
.Y(n_2415)
);

XOR2xp5_ASAP7_75t_L g2416 ( 
.A(n_2415),
.B(n_2412),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2414),
.B(n_2413),
.Y(n_2417)
);

NOR3xp33_ASAP7_75t_L g2418 ( 
.A(n_2417),
.B(n_2174),
.C(n_2177),
.Y(n_2418)
);

CKINVDCx20_ASAP7_75t_R g2419 ( 
.A(n_2416),
.Y(n_2419)
);

BUFx2_ASAP7_75t_L g2420 ( 
.A(n_2417),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2420),
.B(n_2174),
.Y(n_2421)
);

AOI22xp5_ASAP7_75t_SL g2422 ( 
.A1(n_2419),
.A2(n_2019),
.B1(n_2195),
.B2(n_2183),
.Y(n_2422)
);

OA21x2_ASAP7_75t_L g2423 ( 
.A1(n_2421),
.A2(n_2418),
.B(n_2167),
.Y(n_2423)
);

AOI22xp33_ASAP7_75t_SL g2424 ( 
.A1(n_2422),
.A2(n_2173),
.B1(n_2167),
.B2(n_2186),
.Y(n_2424)
);

AOI22xp5_ASAP7_75t_L g2425 ( 
.A1(n_2424),
.A2(n_2183),
.B1(n_2172),
.B2(n_2173),
.Y(n_2425)
);

AOI221xp5_ASAP7_75t_L g2426 ( 
.A1(n_2425),
.A2(n_2423),
.B1(n_2186),
.B2(n_2172),
.C(n_2121),
.Y(n_2426)
);

AOI211xp5_ASAP7_75t_L g2427 ( 
.A1(n_2426),
.A2(n_2193),
.B(n_2152),
.C(n_2137),
.Y(n_2427)
);


endmodule