module fake_jpeg_23199_n_202 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_0),
.C(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_31),
.Y(n_41)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_19),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_25),
.B1(n_14),
.B2(n_17),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_45),
.B1(n_26),
.B2(n_22),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_14),
.B1(n_17),
.B2(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_24),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_52),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_23),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_54),
.Y(n_70)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_29),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_23),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_69),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_14),
.B1(n_22),
.B2(n_15),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_58),
.A2(n_15),
.B1(n_48),
.B2(n_42),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_43),
.B1(n_41),
.B2(n_26),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_36),
.B1(n_16),
.B2(n_20),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_34),
.B1(n_44),
.B2(n_39),
.Y(n_91)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_67),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_68),
.Y(n_73)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_29),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_36),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_76),
.B(n_57),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_81),
.B1(n_65),
.B2(n_56),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_78),
.B(n_71),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_57),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_53),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_85),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_34),
.B1(n_54),
.B2(n_39),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_91),
.B1(n_44),
.B2(n_66),
.Y(n_101)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_90),
.B1(n_48),
.B2(n_66),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_97),
.B(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_71),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_28),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_83),
.B(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_101),
.A2(n_108),
.B1(n_81),
.B2(n_38),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_105),
.C(n_92),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_109),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_68),
.C(n_65),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_30),
.B1(n_80),
.B2(n_87),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_38),
.B1(n_56),
.B2(n_37),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_88),
.B(n_79),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_110),
.A2(n_111),
.B(n_113),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_79),
.B(n_77),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_118),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_93),
.B(n_105),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_120),
.B1(n_125),
.B2(n_127),
.Y(n_143)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_86),
.B(n_107),
.C(n_99),
.D(n_101),
.Y(n_117)
);

AOI221xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_104),
.B1(n_94),
.B2(n_72),
.C(n_37),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_100),
.A2(n_91),
.B(n_75),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_126),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_107),
.A2(n_67),
.B1(n_52),
.B2(n_51),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_80),
.B1(n_72),
.B2(n_37),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_141),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_137),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_127),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_134),
.Y(n_145)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_28),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_125),
.C(n_126),
.Y(n_144)
);

XNOR2x1_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_28),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_113),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_28),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_114),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_148),
.C(n_30),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_135),
.B(n_117),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_149),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_110),
.B(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_153),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_112),
.C(n_116),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_96),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_129),
.B1(n_137),
.B2(n_142),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_30),
.B1(n_19),
.B2(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_139),
.Y(n_159)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_1),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_143),
.B1(n_140),
.B2(n_139),
.Y(n_157)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_162),
.C(n_163),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_130),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_19),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_159),
.C(n_163),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_145),
.A2(n_13),
.B1(n_12),
.B2(n_3),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_166),
.A2(n_156),
.B1(n_144),
.B2(n_148),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_4),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_164),
.B(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_174),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_147),
.B(n_156),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_177),
.Y(n_180)
);

NOR2xp67_ASAP7_75t_SL g173 ( 
.A(n_168),
.B(n_150),
.Y(n_173)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_178),
.B(n_161),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_2),
.B(n_3),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_176),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_4),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_5),
.C(n_6),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_177),
.B(n_160),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_179),
.B(n_185),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_11),
.B1(n_8),
.B2(n_9),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_169),
.B(n_5),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_184),
.A2(n_169),
.B1(n_178),
.B2(n_8),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_189),
.C(n_191),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_5),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_190),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_181),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_180),
.A2(n_7),
.B(n_9),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_7),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_195),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_10),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_SL g197 ( 
.A(n_193),
.B(n_191),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_11),
.B(n_196),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_192),
.A2(n_10),
.B(n_11),
.Y(n_198)
);

BUFx24_ASAP7_75t_SL g199 ( 
.A(n_198),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_199),
.Y(n_202)
);


endmodule