module fake_jpeg_20811_n_302 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_35),
.Y(n_44)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_7),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_28),
.B(n_18),
.Y(n_51)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_43),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_53),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_24),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_21),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_30),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_68),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_34),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_49),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_28),
.B1(n_25),
.B2(n_18),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_63),
.B1(n_66),
.B2(n_77),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_28),
.B1(n_32),
.B2(n_25),
.Y(n_63)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_28),
.B1(n_25),
.B2(n_17),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_67),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_24),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_71),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_20),
.Y(n_100)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_74),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_18),
.B1(n_20),
.B2(n_19),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_78),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_37),
.B1(n_33),
.B2(n_38),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_81),
.A2(n_76),
.B1(n_92),
.B2(n_55),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_37),
.B(n_33),
.C(n_22),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_98),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_21),
.B1(n_15),
.B2(n_20),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_27),
.B1(n_17),
.B2(n_18),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_102),
.B1(n_78),
.B2(n_61),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_27),
.B1(n_17),
.B2(n_15),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_99),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_64),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_22),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_54),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_100),
.B(n_22),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_58),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_72),
.A2(n_58),
.B1(n_74),
.B2(n_70),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_106),
.Y(n_131)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_27),
.A3(n_30),
.B1(n_21),
.B2(n_23),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_14),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

OR2x4_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_30),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_29),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_110),
.B(n_116),
.Y(n_154)
);

INVx2_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_R g145 ( 
.A(n_113),
.B(n_122),
.Y(n_145)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_56),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_118),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_99),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_107),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_121),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_94),
.Y(n_121)
);

OR2x2_ASAP7_75t_SL g122 ( 
.A(n_82),
.B(n_14),
.Y(n_122)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_85),
.B(n_23),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_129),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_126),
.A2(n_97),
.B(n_89),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_88),
.B1(n_81),
.B2(n_87),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_85),
.B(n_23),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_94),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_81),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_101),
.Y(n_135)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_135),
.Y(n_183)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_138),
.A2(n_114),
.B1(n_96),
.B2(n_124),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_132),
.A2(n_116),
.B1(n_122),
.B2(n_113),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_142),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_84),
.C(n_103),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_150),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_89),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_146),
.B(n_147),
.Y(n_190)
);

XOR2x1_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_13),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_83),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_155),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_127),
.B(n_115),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_112),
.A2(n_123),
.B1(n_128),
.B2(n_113),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_151),
.A2(n_164),
.B1(n_133),
.B2(n_111),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_111),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_158),
.C(n_119),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_127),
.A2(n_92),
.B(n_76),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_157),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_112),
.A2(n_55),
.B1(n_83),
.B2(n_96),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_159),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_165),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_80),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_163),
.B(n_134),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_96),
.B1(n_86),
.B2(n_80),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_65),
.C(n_62),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_175),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_153),
.B(n_130),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_149),
.B(n_121),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_179),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_161),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_186),
.B1(n_159),
.B2(n_144),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_139),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_188),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_138),
.A2(n_124),
.B1(n_26),
.B2(n_14),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_162),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_14),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_189),
.B(n_193),
.Y(n_203)
);

NAND2x1_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_0),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_192),
.Y(n_207)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_148),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_194),
.B(n_195),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_154),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_160),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_198),
.A2(n_206),
.B1(n_219),
.B2(n_191),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_143),
.C(n_146),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_215),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_172),
.A2(n_140),
.B1(n_144),
.B2(n_145),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_205),
.A2(n_173),
.B1(n_193),
.B2(n_190),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_159),
.B1(n_145),
.B2(n_142),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_8),
.Y(n_210)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_26),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_216),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_29),
.C(n_26),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_26),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_218),
.A2(n_207),
.B1(n_167),
.B2(n_215),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_180),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_226),
.B1(n_208),
.B2(n_168),
.Y(n_251)
);

NOR3xp33_ASAP7_75t_SL g221 ( 
.A(n_209),
.B(n_191),
.C(n_185),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_225),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_199),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_237),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_201),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_SL g226 ( 
.A1(n_198),
.A2(n_206),
.B(n_172),
.C(n_205),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_227),
.A2(n_169),
.B1(n_214),
.B2(n_204),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_182),
.Y(n_228)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_169),
.B1(n_179),
.B2(n_171),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_238),
.Y(n_245)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_231),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_197),
.Y(n_231)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_167),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_234),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_184),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_236),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_173),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_192),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_242),
.B1(n_253),
.B2(n_226),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_218),
.C(n_168),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_2),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_237),
.B(n_214),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_222),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_219),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_250),
.Y(n_254)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_253),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_245),
.A2(n_226),
.B(n_208),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_255),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_246),
.A2(n_221),
.B(n_235),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_SL g257 ( 
.A1(n_240),
.A2(n_226),
.A3(n_224),
.B1(n_222),
.B2(n_9),
.C1(n_11),
.C2(n_5),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_259),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_244),
.Y(n_258)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_261),
.A2(n_262),
.B1(n_247),
.B2(n_3),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_243),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_252),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_241),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_265),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_260),
.A2(n_250),
.B1(n_245),
.B2(n_251),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_267),
.A2(n_274),
.B1(n_276),
.B2(n_4),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_249),
.C(n_248),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_262),
.C(n_6),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_270),
.B(n_272),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_254),
.A2(n_266),
.B1(n_255),
.B2(n_258),
.Y(n_274)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_259),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_275),
.C(n_276),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_268),
.B(n_10),
.Y(n_279)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_277),
.B(n_6),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_280),
.B(n_283),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_281),
.B(n_282),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_271),
.B(n_7),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_13),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_285),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_269),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_291),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_287),
.B(n_286),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g296 ( 
.A1(n_293),
.A2(n_294),
.B(n_288),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_292),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_295),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_289),
.C(n_267),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_289),
.B(n_281),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_9),
.Y(n_300)
);

AOI221xp5_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.C(n_4),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_12),
.Y(n_302)
);


endmodule