module real_jpeg_28144_n_18 (n_17, n_8, n_0, n_2, n_341, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_342, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_341;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_342;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_0),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_0),
.A2(n_27),
.B1(n_60),
.B2(n_61),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_0),
.A2(n_27),
.B1(n_54),
.B2(n_56),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_1),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_175),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_1),
.A2(n_60),
.B1(n_61),
.B2(n_175),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_1),
.A2(n_54),
.B1(n_56),
.B2(n_175),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_2),
.B(n_54),
.Y(n_92)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_2),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_3),
.A2(n_37),
.B1(n_60),
.B2(n_61),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_3),
.A2(n_37),
.B1(n_54),
.B2(n_56),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_4),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_4),
.A2(n_60),
.B1(n_61),
.B2(n_101),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_101),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_4),
.A2(n_54),
.B1(n_56),
.B2(n_101),
.Y(n_245)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_6),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_SL g178 ( 
.A1(n_6),
.A2(n_29),
.B(n_33),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_6),
.B(n_31),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_6),
.A2(n_60),
.B(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_6),
.B(n_60),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_6),
.B(n_75),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_6),
.A2(n_91),
.B1(n_95),
.B2(n_257),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_6),
.A2(n_32),
.B(n_273),
.Y(n_272)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_9),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_133),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_9),
.A2(n_54),
.B1(n_56),
.B2(n_133),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_9),
.A2(n_60),
.B1(n_61),
.B2(n_133),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_10),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

OAI32xp33_ASAP7_75t_L g233 ( 
.A1(n_10),
.A2(n_56),
.A3(n_60),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_11),
.A2(n_51),
.B1(n_60),
.B2(n_61),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_51),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_11),
.A2(n_51),
.B1(n_54),
.B2(n_56),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_49),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_12),
.A2(n_49),
.B1(n_60),
.B2(n_61),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_12),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_180)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g163 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_15),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_164),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_15),
.A2(n_60),
.B1(n_61),
.B2(n_164),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_15),
.A2(n_54),
.B1(n_56),
.B2(n_164),
.Y(n_251)
);

INVx11_ASAP7_75t_SL g55 ( 
.A(n_16),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_17),
.A2(n_25),
.B1(n_26),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_17),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_103),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g170 ( 
.A1(n_17),
.A2(n_60),
.B1(n_61),
.B2(n_103),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_17),
.A2(n_54),
.B1(n_56),
.B2(n_103),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_22),
.B(n_43),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_24),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_79)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_29),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_26),
.A2(n_35),
.B(n_173),
.C(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_31),
.B(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_31),
.B1(n_47),
.B2(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_28),
.A2(n_31),
.B1(n_100),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_28),
.A2(n_31),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_28),
.A2(n_31),
.B1(n_132),
.B2(n_204),
.Y(n_218)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_31),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_32),
.A2(n_68),
.B(n_70),
.C(n_73),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_71),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g281 ( 
.A1(n_32),
.A2(n_61),
.A3(n_71),
.B1(n_274),
.B2(n_282),
.Y(n_281)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_33),
.B(n_173),
.Y(n_274)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_83),
.B(n_337),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_76),
.C(n_78),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_44),
.A2(n_45),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.C(n_64),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_46),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_48),
.A2(n_80),
.B1(n_82),
.B2(n_102),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_50),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_52),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_52),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_52),
.A2(n_64),
.B1(n_142),
.B2(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_58),
.B(n_63),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_53),
.A2(n_58),
.B1(n_63),
.B2(n_112),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_53),
.A2(n_58),
.B1(n_109),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_53),
.A2(n_58),
.B1(n_128),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_53),
.A2(n_58),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_53),
.A2(n_58),
.B1(n_231),
.B2(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_53),
.B(n_173),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_53),
.A2(n_58),
.B1(n_169),
.B2(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_54),
.B(n_57),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_54),
.B(n_262),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_61),
.B1(n_71),
.B2(n_72),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_60),
.B(n_283),
.Y(n_282)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_64),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_74),
.B2(n_75),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_65),
.A2(n_66),
.B1(n_75),
.B2(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_66),
.A2(n_75),
.B1(n_118),
.B2(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_66),
.A2(n_75),
.B1(n_163),
.B2(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_66),
.A2(n_75),
.B1(n_130),
.B2(n_207),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_73),
.B(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_67),
.A2(n_73),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_67),
.A2(n_73),
.B1(n_162),
.B2(n_165),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_67),
.A2(n_73),
.B1(n_165),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_67),
.A2(n_73),
.B1(n_187),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_71),
.Y(n_283)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_74),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_76),
.A2(n_78),
.B1(n_79),
.B2(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_76),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_82),
.B1(n_99),
.B2(n_102),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_80),
.A2(n_82),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_330),
.B(n_336),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_145),
.A3(n_154),
.B1(n_328),
.B2(n_329),
.C(n_341),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_134),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_86),
.B(n_134),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_115),
.C(n_122),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_87),
.B(n_115),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_104),
.B1(n_105),
.B2(n_114),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_97),
.B2(n_98),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_89),
.A2(n_98),
.B(n_104),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_89),
.A2(n_90),
.B1(n_106),
.B2(n_107),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_93),
.B(n_96),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_93),
.B1(n_96),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_91),
.A2(n_93),
.B1(n_126),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_91),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_91),
.A2(n_95),
.B1(n_251),
.B2(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_91),
.A2(n_93),
.B1(n_245),
.B2(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_92),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_92),
.A2(n_94),
.B1(n_180),
.B2(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_92),
.A2(n_94),
.B1(n_250),
.B2(n_252),
.Y(n_249)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_93),
.Y(n_181)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_SL g246 ( 
.A(n_94),
.Y(n_246)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_110),
.A2(n_113),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_110),
.A2(n_113),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_120),
.B(n_121),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_120),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_119),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_121),
.B(n_135),
.CI(n_144),
.CON(n_134),
.SN(n_134)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_135),
.C(n_144),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_122),
.A2(n_123),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.C(n_131),
.Y(n_123)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_124),
.B(n_129),
.CI(n_131),
.CON(n_311),
.SN(n_311)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_125),
.B(n_127),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_134),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_143),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_137),
.B1(n_149),
.B2(n_152),
.Y(n_148)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_139),
.C(n_142),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_137),
.B(n_152),
.C(n_153),
.Y(n_331)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_146),
.B(n_147),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_153),
.Y(n_147)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_149),
.Y(n_152)
);

AOI321xp33_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_309),
.A3(n_317),
.B1(n_322),
.B2(n_327),
.C(n_342),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_209),
.C(n_221),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_191),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_157),
.B(n_191),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_176),
.C(n_183),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_158),
.B(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_171),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_166),
.B2(n_167),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_167),
.C(n_171),
.Y(n_198)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_170),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_173),
.B(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_174),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_176),
.A2(n_183),
.B1(n_184),
.B2(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_176),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_179),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_182),
.Y(n_197)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.C(n_190),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_185),
.B(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_188),
.B(n_190),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_189),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_199),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_198),
.C(n_199),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_196),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_208),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_205),
.C(n_208),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g323 ( 
.A1(n_210),
.A2(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_211),
.B(n_212),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_220),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_214),
.B(n_215),
.C(n_220),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_216),
.B(n_218),
.C(n_219),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_303),
.B(n_308),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_289),
.B(n_302),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_267),
.B(n_288),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_247),
.B(n_266),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_236),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_226),
.B(n_236),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_232),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_227),
.A2(n_228),
.B1(n_232),
.B2(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_230),
.Y(n_234)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_243),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_241),
.C(n_243),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_242),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_244),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_254),
.B(n_265),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_253),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_259),
.B(n_264),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_256),
.B(n_258),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_268),
.B(n_269),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_280),
.B1(n_286),
.B2(n_287),
.Y(n_269)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_275),
.B1(n_278),
.B2(n_279),
.Y(n_270)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_279),
.C(n_287),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_277),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_280),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_284),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_284),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_290),
.B(n_291),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_298),
.C(n_300),
.Y(n_304)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_300),
.B2(n_301),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_297),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_298),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_314),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_314),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.C(n_313),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_312),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_311),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_318),
.A2(n_323),
.B(n_326),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_319),
.B(n_320),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);


endmodule