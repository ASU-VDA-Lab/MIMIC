module fake_jpeg_267_n_57 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_57);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_57;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx11_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_21),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_18),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

AO22x2_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_25),
.A2(n_21),
.B1(n_18),
.B2(n_19),
.Y(n_26)
);

A2O1A1O1Ixp25_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_28),
.B(n_30),
.C(n_19),
.D(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_18),
.Y(n_28)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_34),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_22),
.B1(n_20),
.B2(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_40),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_24),
.B1(n_16),
.B2(n_20),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_16),
.B1(n_17),
.B2(n_12),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_19),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_16),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_2),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_44),
.B(n_3),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_39),
.B(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_3),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_41),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_49),
.C(n_5),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_10),
.B(n_6),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_4),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_51),
.C(n_46),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_5),
.B(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

NOR3xp33_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_54),
.C(n_9),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_10),
.B(n_8),
.Y(n_57)
);


endmodule