module real_jpeg_12840_n_27 (n_17, n_123, n_8, n_0, n_21, n_2, n_125, n_10, n_9, n_12, n_124, n_24, n_6, n_121, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_127, n_119, n_5, n_4, n_122, n_1, n_26, n_20, n_19, n_118, n_126, n_16, n_15, n_13, n_120, n_27);

input n_17;
input n_123;
input n_8;
input n_0;
input n_21;
input n_2;
input n_125;
input n_10;
input n_9;
input n_12;
input n_124;
input n_24;
input n_6;
input n_121;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_127;
input n_119;
input n_5;
input n_4;
input n_122;
input n_1;
input n_26;
input n_20;
input n_19;
input n_118;
input n_126;
input n_16;
input n_15;
input n_13;
input n_120;

output n_27;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_116;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_0),
.Y(n_111)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_1),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_2),
.B(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_3),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_4),
.B(n_66),
.C(n_77),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_5),
.B(n_46),
.C(n_94),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_6),
.B(n_54),
.C(n_83),
.Y(n_53)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

MAJx2_ASAP7_75t_L g43 ( 
.A(n_8),
.B(n_44),
.C(n_100),
.Y(n_43)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_9),
.B(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_10),
.B(n_56),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_12),
.Y(n_76)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_12),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_14),
.B(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_14),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_15),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_43),
.C(n_103),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_17),
.Y(n_108)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_18),
.B(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_41),
.C(n_110),
.Y(n_40)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_48),
.C(n_86),
.Y(n_47)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_60),
.C(n_80),
.Y(n_59)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_39),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_33),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_33),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_33),
.B(n_104),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_33),
.B(n_111),
.Y(n_110)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_34),
.B(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_36),
.B(n_81),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_37),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_37),
.B(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_105),
.C(n_106),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_96),
.C(n_97),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_90),
.C(n_91),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_52),
.B(n_53),
.C(n_85),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_58),
.B(n_59),
.C(n_82),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_64),
.B(n_65),
.C(n_79),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_72),
.C(n_73),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_118),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_119),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_120),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_121),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_122),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_123),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_124),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_125),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_126),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_127),
.Y(n_93)
);


endmodule