module fake_jpeg_9660_n_331 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_5),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_26),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_38),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx3_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_18),
.Y(n_46)
);

OR2x2_ASAP7_75t_SL g80 ( 
.A(n_46),
.B(n_20),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_23),
.B1(n_21),
.B2(n_32),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_59),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_32),
.B1(n_21),
.B2(n_23),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_56),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_23),
.B1(n_21),
.B2(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_57),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_63),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_23),
.B1(n_22),
.B2(n_33),
.Y(n_59)
);

CKINVDCx6p67_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_20),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_52),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_26),
.B1(n_33),
.B2(n_25),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_25),
.B1(n_33),
.B2(n_20),
.Y(n_89)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_45),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_31),
.B1(n_26),
.B2(n_25),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_94),
.B1(n_89),
.B2(n_74),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_76),
.Y(n_102)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_43),
.C(n_39),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_90),
.C(n_47),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_43),
.C(n_19),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_81),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_46),
.Y(n_98)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_93),
.Y(n_101)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_96),
.B1(n_73),
.B2(n_88),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_65),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_46),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_92),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_53),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_31),
.B1(n_34),
.B2(n_19),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_28),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_86),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_46),
.Y(n_96)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_107),
.C(n_112),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_79),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_106),
.B1(n_104),
.B2(n_111),
.Y(n_131)
);

AOI32xp33_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_61),
.A3(n_53),
.B1(n_60),
.B2(n_36),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_119),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_60),
.B1(n_53),
.B2(n_47),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_68),
.C(n_58),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_124),
.Y(n_132)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_116),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_70),
.C(n_56),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_80),
.B1(n_73),
.B2(n_85),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_68),
.C(n_39),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_54),
.Y(n_146)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_120),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_82),
.A2(n_60),
.B1(n_68),
.B2(n_67),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_118),
.A2(n_84),
.B1(n_80),
.B2(n_93),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_36),
.A3(n_27),
.B1(n_34),
.B2(n_42),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_121),
.A2(n_123),
.B1(n_83),
.B2(n_81),
.Y(n_134)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_137),
.B1(n_144),
.B2(n_119),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_124),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_128),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_78),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_77),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_138),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_131),
.A2(n_133),
.B1(n_144),
.B2(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_135),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_72),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_140),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_71),
.B(n_77),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_147),
.B(n_30),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_98),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_76),
.B1(n_83),
.B2(n_84),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_99),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_145),
.A2(n_118),
.B1(n_97),
.B2(n_98),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_115),
.C(n_127),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_0),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_148),
.A2(n_117),
.B1(n_105),
.B2(n_103),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_110),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_24),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_67),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_151),
.B(n_110),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_153),
.B(n_159),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_176),
.C(n_180),
.Y(n_188)
);

NAND4xp25_ASAP7_75t_SL g156 ( 
.A(n_135),
.B(n_62),
.C(n_55),
.D(n_17),
.Y(n_156)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_163),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_131),
.B1(n_141),
.B2(n_145),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_162),
.A2(n_175),
.B1(n_34),
.B2(n_27),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_132),
.B(n_104),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_129),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_178),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_172),
.B1(n_173),
.B2(n_149),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_166),
.A2(n_142),
.B(n_147),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_34),
.B1(n_31),
.B2(n_27),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_130),
.B(n_112),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_168),
.B(n_171),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_128),
.A2(n_42),
.B1(n_41),
.B2(n_19),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_177),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_137),
.A2(n_42),
.B1(n_41),
.B2(n_30),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_127),
.B(n_39),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_54),
.C(n_62),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_181),
.B(n_171),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_183),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_149),
.Y(n_184)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

A2O1A1O1Ixp25_ASAP7_75t_L g185 ( 
.A1(n_168),
.A2(n_142),
.B(n_125),
.C(n_147),
.D(n_54),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_201),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g186 ( 
.A1(n_178),
.A2(n_41),
.B(n_148),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_191),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_54),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_180),
.C(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_192),
.B(n_196),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_194),
.A2(n_197),
.B(n_207),
.Y(n_215)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_169),
.Y(n_202)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_165),
.A2(n_143),
.B1(n_24),
.B2(n_30),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_167),
.A2(n_143),
.B1(n_24),
.B2(n_55),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_154),
.A2(n_31),
.B1(n_34),
.B2(n_54),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_29),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_221),
.C(n_227),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_154),
.B1(n_175),
.B2(n_174),
.Y(n_211)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_187),
.A2(n_170),
.B1(n_160),
.B2(n_162),
.Y(n_214)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_157),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_223),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_157),
.Y(n_221)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_199),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_226),
.B(n_228),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_177),
.C(n_45),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_189),
.A2(n_161),
.B(n_179),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_179),
.B1(n_31),
.B2(n_2),
.Y(n_229)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_45),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_232),
.C(n_190),
.Y(n_243)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_45),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_183),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_233),
.A2(n_0),
.B(n_1),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_219),
.B(n_195),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_252),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_199),
.B(n_186),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_240),
.A2(n_251),
.B(n_14),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_226),
.A2(n_195),
.B1(n_205),
.B2(n_194),
.Y(n_241)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_249),
.C(n_250),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_184),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_184),
.C(n_204),
.Y(n_250)
);

XOR2x2_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_182),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_29),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_254),
.C(n_255),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_29),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_213),
.B(n_29),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_220),
.B(n_16),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_256),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_227),
.C(n_210),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_263),
.C(n_267),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_247),
.A2(n_215),
.B(n_212),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_261),
.A2(n_264),
.B(n_234),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_251),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_255),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_232),
.C(n_223),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_212),
.B(n_222),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_222),
.C(n_233),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_268),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_235),
.A2(n_224),
.B1(n_231),
.B2(n_15),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_269),
.B(n_273),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_236),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_270),
.A2(n_248),
.B1(n_241),
.B2(n_252),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_237),
.B(n_244),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_245),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_29),
.C(n_3),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_257),
.C(n_258),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_262),
.A2(n_260),
.B1(n_266),
.B2(n_246),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_275),
.A2(n_283),
.B(n_284),
.Y(n_296)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_274),
.B1(n_270),
.B2(n_258),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_242),
.C(n_243),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_289),
.C(n_29),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_268),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_287),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_286),
.B(n_288),
.Y(n_298)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_267),
.A2(n_242),
.B1(n_253),
.B2(n_254),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_261),
.C(n_263),
.Y(n_289)
);

OAI21x1_ASAP7_75t_SL g291 ( 
.A1(n_279),
.A2(n_271),
.B(n_265),
.Y(n_291)
);

OAI22x1_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_292),
.B1(n_284),
.B2(n_281),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_272),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_12),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_297),
.C(n_300),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_2),
.C(n_3),
.Y(n_297)
);

FAx1_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_3),
.CI(n_4),
.CON(n_299),
.SN(n_299)
);

NAND2x1p5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_301),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_4),
.C(n_5),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_275),
.A2(n_14),
.B(n_13),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_301),
.A2(n_278),
.B(n_299),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_308),
.Y(n_314)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_304),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_276),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_306),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_289),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_311),
.C(n_299),
.Y(n_315)
);

OAI33xp33_ASAP7_75t_L g308 ( 
.A1(n_290),
.A2(n_283),
.A3(n_280),
.B1(n_288),
.B2(n_282),
.B3(n_11),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_302),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_310),
.A2(n_303),
.B1(n_296),
.B2(n_7),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_298),
.A2(n_13),
.B(n_12),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_11),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_319),
.C(n_320),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_318),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_294),
.B(n_295),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_310),
.A2(n_296),
.B(n_6),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_316),
.A2(n_5),
.B(n_7),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_321),
.B(n_323),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_313),
.A2(n_8),
.B(n_9),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_8),
.C(n_9),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_324),
.A2(n_317),
.B1(n_314),
.B2(n_10),
.Y(n_327)
);

AO21x1_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_325),
.B(n_322),
.Y(n_328)
);

NAND3xp33_ASAP7_75t_SL g329 ( 
.A(n_328),
.B(n_326),
.C(n_9),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_8),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_10),
.B(n_317),
.Y(n_331)
);


endmodule