module fake_jpeg_26116_n_83 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_42),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_1),
.B(n_2),
.Y(n_41)
);

FAx1_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_3),
.CI(n_7),
.CON(n_51),
.SN(n_51)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_1),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_37),
.B1(n_31),
.B2(n_38),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_26),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_37),
.B1(n_39),
.B2(n_4),
.Y(n_49)
);

AO21x1_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_50),
.B(n_56),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_18),
.B(n_19),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_21),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_20),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_59),
.B(n_61),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_63),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_64),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_30),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_71),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_70),
.B(n_68),
.Y(n_75)
);

AOI221xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_70),
.B1(n_75),
.B2(n_68),
.C(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_75),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_73),
.C(n_72),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_65),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_64),
.C(n_67),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_28),
.B(n_29),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_66),
.Y(n_83)
);


endmodule