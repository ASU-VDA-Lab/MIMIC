module fake_jpeg_3118_n_176 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_176);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_10),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_25),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_2),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_21),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_68),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_65),
.B(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_0),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_74),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_65),
.B(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_65),
.B(n_54),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_50),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_55),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_51),
.Y(n_90)
);

BUFx2_ASAP7_75t_SL g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_91),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_64),
.B1(n_58),
.B2(n_60),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_56),
.B1(n_2),
.B2(n_3),
.Y(n_117)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_46),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_57),
.B1(n_58),
.B2(n_67),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_97),
.B(n_56),
.C(n_52),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_45),
.B(n_56),
.C(n_57),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_62),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_0),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_56),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_103),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_78),
.B(n_67),
.C(n_45),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_40),
.B1(n_37),
.B2(n_35),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_97),
.A2(n_78),
.B1(n_80),
.B2(n_49),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_110),
.A2(n_97),
.B1(n_94),
.B2(n_87),
.Y(n_125)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_116),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_20),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_1),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_94),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_114),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_119),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_134),
.B1(n_137),
.B2(n_9),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_85),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_127),
.Y(n_145)
);

AO21x1_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_28),
.B(n_27),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_97),
.B1(n_89),
.B2(n_41),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_26),
.B1(n_19),
.B2(n_12),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_114),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_1),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_4),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_132),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_102),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_101),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_100),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_139),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_105),
.C(n_33),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_125),
.A2(n_105),
.B1(n_30),
.B2(n_29),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_134),
.B1(n_137),
.B2(n_129),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_146),
.B(n_147),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_8),
.B(n_9),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_136),
.B(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_149),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_10),
.C(n_11),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_11),
.C(n_12),
.Y(n_152)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_154),
.B(n_161),
.Y(n_166)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_144),
.A2(n_132),
.B1(n_131),
.B2(n_15),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_160),
.A2(n_145),
.A3(n_143),
.B1(n_155),
.B2(n_157),
.C1(n_161),
.C2(n_138),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_162),
.A2(n_164),
.B1(n_165),
.B2(n_13),
.Y(n_169)
);

NAND4xp25_ASAP7_75t_SL g164 ( 
.A(n_154),
.B(n_142),
.C(n_150),
.D(n_153),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_156),
.A2(n_141),
.A3(n_132),
.B1(n_139),
.B2(n_152),
.C1(n_151),
.C2(n_16),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_158),
.C(n_14),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_169),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_158),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_166),
.C(n_14),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_168),
.C(n_15),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_171),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_13),
.B(n_17),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);


endmodule