module real_jpeg_6949_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_1),
.Y(n_127)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_1),
.Y(n_129)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_1),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_1),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_1),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_1),
.Y(n_144)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_1),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_1),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_1),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_2),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_2),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_2),
.A2(n_243),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_2),
.A2(n_243),
.B1(n_411),
.B2(n_413),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_2),
.A2(n_243),
.B1(n_466),
.B2(n_471),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_3),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_4),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_4),
.A2(n_47),
.B1(n_159),
.B2(n_161),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_4),
.A2(n_47),
.B1(n_140),
.B2(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_4),
.A2(n_47),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_5),
.B(n_275),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_5),
.A2(n_274),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_5),
.B(n_194),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_5),
.B(n_161),
.C(n_384),
.Y(n_383)
);

OAI22xp33_ASAP7_75t_L g387 ( 
.A1(n_5),
.A2(n_388),
.B1(n_389),
.B2(n_391),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_5),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_5),
.B(n_98),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_5),
.A2(n_151),
.B1(n_432),
.B2(n_435),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_6),
.A2(n_265),
.B1(n_291),
.B2(n_293),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_6),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_6),
.A2(n_293),
.B1(n_355),
.B2(n_356),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_6),
.A2(n_293),
.B1(n_395),
.B2(n_398),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_6),
.A2(n_293),
.B1(n_416),
.B2(n_433),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_7),
.A2(n_296),
.B1(n_298),
.B2(n_299),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_7),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_7),
.A2(n_298),
.B1(n_329),
.B2(n_333),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_7),
.A2(n_298),
.B1(n_406),
.B2(n_407),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_7),
.A2(n_216),
.B1(n_298),
.B2(n_422),
.Y(n_421)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_9),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_9),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_9),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_9),
.Y(n_314)
);

INVx8_ASAP7_75t_L g349 ( 
.A(n_9),
.Y(n_349)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_9),
.Y(n_437)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_10),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_10),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_10),
.A2(n_67),
.B1(n_77),
.B2(n_115),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_10),
.A2(n_67),
.B1(n_133),
.B2(n_136),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_10),
.A2(n_67),
.B1(n_216),
.B2(n_221),
.Y(n_215)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_13),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_13),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_13),
.Y(n_142)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_13),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_13),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_14),
.A2(n_100),
.B1(n_101),
.B2(n_105),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_14),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_14),
.A2(n_100),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_14),
.A2(n_100),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_14),
.A2(n_100),
.B1(n_285),
.B2(n_288),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_17),
.A2(n_73),
.B1(n_76),
.B2(n_77),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_17),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_17),
.A2(n_76),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_17),
.A2(n_76),
.B1(n_233),
.B2(n_235),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_17),
.A2(n_76),
.B1(n_217),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_202),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_200),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_175),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_27),
.B(n_175),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_27),
.B(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_27),
.B(n_204),
.Y(n_501)
);

FAx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_107),
.CI(n_149),
.CON(n_27),
.SN(n_27)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_28),
.A2(n_29),
.B(n_70),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_70),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_51),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_30),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_41),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_31),
.A2(n_41),
.B(n_52),
.Y(n_110)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_31),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_31),
.A2(n_52),
.B1(n_62),
.B2(n_232),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_31),
.B(n_388),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_32)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_34),
.Y(n_161)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g153 ( 
.A(n_36),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_36),
.Y(n_160)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_36),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_38),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_38),
.Y(n_412)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_38),
.Y(n_416)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_40),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_41),
.A2(n_52),
.B(n_169),
.Y(n_321)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_42),
.Y(n_166)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_44),
.Y(n_397)
);

INVx6_ASAP7_75t_L g454 ( 
.A(n_44),
.Y(n_454)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_45),
.Y(n_470)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_46),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g390 ( 
.A(n_46),
.Y(n_390)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_46),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_80),
.B1(n_82),
.B2(n_85),
.Y(n_79)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_50),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_62),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_52),
.A2(n_164),
.B(n_169),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_52),
.A2(n_484),
.B(n_485),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_53),
.A2(n_165),
.B1(n_170),
.B2(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_53),
.A2(n_170),
.B1(n_387),
.B2(n_394),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_53),
.A2(n_170),
.B1(n_394),
.B2(n_405),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_53),
.A2(n_170),
.B1(n_405),
.B2(n_465),
.Y(n_464)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_61),
.Y(n_54)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_55),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_61),
.Y(n_399)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_63),
.B(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_66),
.Y(n_406)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_69),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_78),
.B1(n_98),
.B2(n_99),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_72),
.A2(n_79),
.B(n_191),
.Y(n_247)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_73),
.Y(n_256)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_75),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_75),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_99),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_78),
.B(n_114),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_78),
.A2(n_184),
.B(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_78),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_78),
.A2(n_98),
.B1(n_354),
.B2(n_463),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_87),
.Y(n_78)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_79),
.B(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_79),
.A2(n_308),
.B1(n_328),
.B2(n_336),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_79),
.A2(n_308),
.B1(n_328),
.B2(n_353),
.Y(n_352)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx6_ASAP7_75t_L g455 ( 
.A(n_82),
.Y(n_455)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_84),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_91),
.B1(n_94),
.B2(n_97),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_90),
.Y(n_264)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_96),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_114),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_SL g463 ( 
.A1(n_101),
.A2(n_388),
.B(n_456),
.Y(n_463)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_103),
.Y(n_355)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_104),
.Y(n_106)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_118),
.B2(n_148),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_116),
.B2(n_117),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_110),
.A2(n_117),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_111),
.B(n_117),
.C(n_118),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_113),
.A2(n_185),
.B(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_118),
.A2(n_148),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_125),
.B(n_130),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_119),
.B(n_132),
.Y(n_174)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_119),
.A2(n_138),
.B1(n_240),
.B2(n_295),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_119),
.A2(n_138),
.B1(n_323),
.B2(n_326),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_126),
.Y(n_244)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_128),
.Y(n_265)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_129),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_137),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_134),
.Y(n_297)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_136),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_172),
.B(n_174),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_137),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_137),
.A2(n_194),
.B1(n_290),
.B2(n_294),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_138),
.A2(n_240),
.B(n_245),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_145),
.Y(n_139)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_147),
.Y(n_272)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_162),
.B(n_171),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_150),
.A2(n_171),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_150),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_150),
.A2(n_163),
.B1(n_207),
.B2(n_366),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_156),
.B(n_158),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_151),
.B(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_151),
.A2(n_278),
.B1(n_283),
.B2(n_284),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_151),
.A2(n_284),
.B(n_313),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_151),
.A2(n_224),
.B(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_151),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_151),
.A2(n_421),
.B1(n_432),
.B2(n_435),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_151),
.A2(n_158),
.B(n_313),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_155),
.Y(n_426)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_163),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_172),
.B(n_194),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_192),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_191),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx8_ASAP7_75t_L g451 ( 
.A(n_186),
.Y(n_451)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_190),
.Y(n_332)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_190),
.Y(n_335)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_196),
.Y(n_292)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_197),
.Y(n_276)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_248),
.B(n_500),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_209),
.C(n_210),
.Y(n_204)
);

FAx1_ASAP7_75t_L g374 ( 
.A(n_205),
.B(n_209),
.CI(n_210),
.CON(n_374),
.SN(n_374)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_238),
.C(n_246),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_211),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_229),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_212),
.A2(n_229),
.B1(n_230),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_212),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_224),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_214),
.A2(n_279),
.B(n_345),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_215),
.Y(n_315)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_218),
.Y(n_434)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_219),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_220),
.Y(n_287)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_222),
.B(n_441),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_228),
.Y(n_283)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_238),
.A2(n_239),
.B1(n_246),
.B2(n_247),
.Y(n_368)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_375),
.B(n_494),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_360),
.C(n_372),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_338),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_251),
.A2(n_496),
.B(n_497),
.Y(n_495)
);

NOR2xp67_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_317),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_252),
.B(n_317),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_301),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_253),
.B(n_302),
.C(n_304),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_260),
.C(n_289),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_254),
.B(n_289),
.Y(n_319)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_255),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_259),
.B(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_260),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_277),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_261),
.B(n_277),
.Y(n_341)
);

OAI32xp33_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_265),
.A3(n_266),
.B1(n_270),
.B2(n_273),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g357 ( 
.A(n_264),
.Y(n_357)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVxp33_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_282),
.Y(n_422)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_290),
.Y(n_326)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_311),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_309),
.B2(n_310),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_306),
.B(n_310),
.C(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_311),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_316),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_316),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_320),
.C(n_337),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_320),
.B(n_337),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.C(n_327),
.Y(n_320)
);

FAx1_ASAP7_75t_L g340 ( 
.A(n_321),
.B(n_322),
.CI(n_327),
.CON(n_340),
.SN(n_340)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_333),
.B(n_388),
.Y(n_456)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_358),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_339),
.B(n_358),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.C(n_342),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_340),
.B(n_492),
.Y(n_491)
);

BUFx24_ASAP7_75t_SL g502 ( 
.A(n_340),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_341),
.B(n_342),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_350),
.C(n_352),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_343),
.A2(n_344),
.B1(n_350),
.B2(n_351),
.Y(n_479)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_346),
.B(n_388),
.Y(n_441)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx8_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_352),
.B(n_479),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

A2O1A1O1Ixp25_ASAP7_75t_L g494 ( 
.A1(n_360),
.A2(n_372),
.B(n_495),
.C(n_498),
.D(n_499),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_361),
.B(n_371),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_361),
.B(n_371),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_362),
.B(n_365),
.C(n_370),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_367),
.B1(n_369),
.B2(n_370),
.Y(n_364)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_365),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_367),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_373),
.B(n_374),
.Y(n_499)
);

BUFx24_ASAP7_75t_SL g504 ( 
.A(n_374),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_489),
.B(n_493),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_474),
.B(n_488),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_445),
.B(n_473),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_379),
.A2(n_417),
.B(n_444),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_400),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_380),
.B(n_400),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_386),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_381),
.B(n_386),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx3_ASAP7_75t_SL g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_390),
.Y(n_472)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_393),
.Y(n_407)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_409),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_403),
.B1(n_404),
.B2(n_408),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_402),
.B(n_408),
.C(n_409),
.Y(n_446)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_404),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_407),
.B(n_458),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_410),
.Y(n_424)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_428),
.B(n_443),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_427),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_427),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_420),
.A2(n_423),
.B1(n_424),
.B2(n_425),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_429),
.A2(n_438),
.B(n_442),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_430),
.B(n_431),
.Y(n_442)
);

INVx4_ASAP7_75t_SL g433 ( 
.A(n_434),
.Y(n_433)
);

INVx5_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_446),
.B(n_447),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_461),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_448),
.B(n_462),
.C(n_464),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_449),
.B(n_460),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_449),
.B(n_460),
.Y(n_482)
);

OAI32xp33_ASAP7_75t_L g449 ( 
.A1(n_450),
.A2(n_452),
.A3(n_455),
.B1(n_456),
.B2(n_457),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx6_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_464),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_465),
.Y(n_484)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_475),
.B(n_476),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_477),
.A2(n_478),
.B1(n_480),
.B2(n_481),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_477),
.B(n_483),
.C(n_486),
.Y(n_490)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_482),
.A2(n_483),
.B1(n_486),
.B2(n_487),
.Y(n_481)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_482),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_483),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_490),
.B(n_491),
.Y(n_493)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);


endmodule