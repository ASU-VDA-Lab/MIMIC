module fake_netlist_1_7889_n_1143 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_280, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1143);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1143;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_564;
wire n_353;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_476;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1125;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_1094;
wire n_652;
wire n_968;
wire n_303;
wire n_1060;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_529;
wire n_312;
wire n_1011;
wire n_1025;
wire n_1132;
wire n_880;
wire n_1101;
wire n_630;
wire n_511;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_624;
wire n_426;
wire n_725;
wire n_818;
wire n_769;
wire n_844;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_828;
wire n_767;
wire n_1063;
wire n_293;
wire n_1138;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_1046;
wire n_478;
wire n_482;
wire n_415;
wire n_394;
wire n_703;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_805;
wire n_729;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_666;
wire n_621;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_806;
wire n_881;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_955;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1069;
wire n_1123;
wire n_811;
wire n_1021;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_924;
wire n_912;
wire n_947;
wire n_1043;
wire n_582;
wire n_378;
wire n_1141;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_1127;
INVxp67_ASAP7_75t_SL g282 ( .A(n_33), .Y(n_282) );
INVxp33_ASAP7_75t_SL g283 ( .A(n_102), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_180), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g285 ( .A(n_68), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_24), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_230), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_252), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_114), .Y(n_289) );
INVxp67_ASAP7_75t_L g290 ( .A(n_121), .Y(n_290) );
INVxp33_ASAP7_75t_L g291 ( .A(n_247), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_213), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_38), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_246), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_234), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_222), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_229), .Y(n_297) );
BUFx10_ASAP7_75t_L g298 ( .A(n_96), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_163), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_211), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_47), .Y(n_301) );
INVxp67_ASAP7_75t_SL g302 ( .A(n_92), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_243), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_127), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_33), .Y(n_305) );
CKINVDCx16_ASAP7_75t_R g306 ( .A(n_195), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_227), .Y(n_307) );
CKINVDCx16_ASAP7_75t_R g308 ( .A(n_24), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_78), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_161), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_98), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_218), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_103), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_249), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_214), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_81), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_128), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_19), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_148), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_260), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_38), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_157), .Y(n_322) );
INVx1_ASAP7_75t_SL g323 ( .A(n_16), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_275), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_257), .Y(n_325) );
CKINVDCx16_ASAP7_75t_R g326 ( .A(n_199), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_82), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_154), .Y(n_328) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_190), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_122), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_65), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_273), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_80), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_35), .Y(n_334) );
CKINVDCx14_ASAP7_75t_R g335 ( .A(n_208), .Y(n_335) );
INVxp67_ASAP7_75t_SL g336 ( .A(n_185), .Y(n_336) );
BUFx10_ASAP7_75t_L g337 ( .A(n_113), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_54), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_110), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_75), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_248), .Y(n_341) );
INVxp67_ASAP7_75t_SL g342 ( .A(n_215), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_240), .B(n_94), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_60), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_244), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_149), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_158), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_203), .Y(n_348) );
INVxp67_ASAP7_75t_SL g349 ( .A(n_217), .Y(n_349) );
INVxp67_ASAP7_75t_SL g350 ( .A(n_196), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_16), .Y(n_351) );
CKINVDCx14_ASAP7_75t_R g352 ( .A(n_27), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_90), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_70), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_81), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_62), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_186), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_11), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_118), .B(n_133), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_97), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_104), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_174), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_166), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_83), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_151), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_124), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_202), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_209), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_116), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_225), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_132), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_120), .Y(n_372) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_223), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_216), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_241), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_144), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_176), .Y(n_377) );
INVx4_ASAP7_75t_R g378 ( .A(n_106), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_236), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_207), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_188), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_13), .Y(n_382) );
INVxp33_ASAP7_75t_SL g383 ( .A(n_267), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_239), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_75), .Y(n_385) );
BUFx10_ASAP7_75t_L g386 ( .A(n_32), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_156), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_238), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_274), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_46), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_268), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_183), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_175), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_95), .Y(n_394) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_210), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_187), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_242), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_77), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_44), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_263), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_181), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_8), .Y(n_402) );
INVxp33_ASAP7_75t_SL g403 ( .A(n_280), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_145), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_251), .Y(n_405) );
INVxp33_ASAP7_75t_SL g406 ( .A(n_85), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_172), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_30), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_93), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_264), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_129), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_269), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_12), .Y(n_413) );
CKINVDCx16_ASAP7_75t_R g414 ( .A(n_189), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_147), .Y(n_415) );
INVxp33_ASAP7_75t_SL g416 ( .A(n_219), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_9), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_134), .Y(n_418) );
BUFx3_ASAP7_75t_L g419 ( .A(n_224), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_13), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_245), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_212), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_165), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_26), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_155), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_142), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_91), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_109), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_87), .B(n_169), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_164), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_69), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_256), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_101), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_347), .B(n_0), .Y(n_434) );
NOR2xp33_ASAP7_75t_R g435 ( .A(n_335), .B(n_84), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_347), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_331), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_347), .B(n_0), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_322), .B(n_1), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_331), .Y(n_440) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_306), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_352), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_291), .B(n_1), .Y(n_443) );
INVx5_ASAP7_75t_L g444 ( .A(n_310), .Y(n_444) );
INVx3_ASAP7_75t_L g445 ( .A(n_298), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_326), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_338), .Y(n_447) );
XNOR2xp5_ASAP7_75t_L g448 ( .A(n_285), .B(n_2), .Y(n_448) );
BUFx2_ASAP7_75t_L g449 ( .A(n_352), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_310), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_298), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_338), .Y(n_452) );
OAI21x1_ASAP7_75t_L g453 ( .A1(n_363), .A2(n_88), .B(n_86), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_308), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_291), .B(n_2), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_358), .Y(n_456) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_310), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_310), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_358), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_287), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_288), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_292), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_315), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_294), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_387), .B(n_3), .Y(n_465) );
INVx6_ASAP7_75t_L g466 ( .A(n_298), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_295), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_315), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_337), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_432), .B(n_4), .Y(n_470) );
BUFx2_ASAP7_75t_L g471 ( .A(n_293), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_436), .Y(n_472) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_457), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_444), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_449), .B(n_414), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_445), .B(n_301), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_466), .B(n_290), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_434), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_445), .B(n_337), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_445), .B(n_284), .Y(n_480) );
NAND3xp33_ASAP7_75t_L g481 ( .A(n_460), .B(n_297), .C(n_296), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_471), .B(n_335), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_466), .B(n_369), .Y(n_483) );
CKINVDCx11_ASAP7_75t_R g484 ( .A(n_454), .Y(n_484) );
INVx4_ASAP7_75t_L g485 ( .A(n_434), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_436), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_466), .B(n_433), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_471), .B(n_305), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_436), .Y(n_489) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_457), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_445), .B(n_301), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_445), .B(n_284), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_436), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_444), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_460), .B(n_303), .C(n_300), .Y(n_495) );
AND2x6_ASAP7_75t_L g496 ( .A(n_434), .B(n_372), .Y(n_496) );
NOR2xp33_ASAP7_75t_SL g497 ( .A(n_441), .B(n_361), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_436), .Y(n_498) );
INVx4_ASAP7_75t_L g499 ( .A(n_434), .Y(n_499) );
NAND3x1_ASAP7_75t_L g500 ( .A(n_443), .B(n_318), .C(n_309), .Y(n_500) );
OAI22xp33_ASAP7_75t_L g501 ( .A1(n_442), .A2(n_285), .B1(n_344), .B2(n_334), .Y(n_501) );
INVx4_ASAP7_75t_L g502 ( .A(n_434), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_443), .B(n_386), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_444), .Y(n_504) );
INVx8_ASAP7_75t_L g505 ( .A(n_438), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_443), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_451), .B(n_299), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_438), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_444), .Y(n_509) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_457), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_466), .B(n_283), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_438), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_466), .B(n_283), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_438), .Y(n_514) );
INVx4_ASAP7_75t_L g515 ( .A(n_438), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_444), .Y(n_516) );
NOR2x2_ASAP7_75t_L g517 ( .A(n_497), .B(n_448), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_476), .B(n_466), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_506), .B(n_451), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_485), .B(n_455), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_506), .B(n_451), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_503), .B(n_451), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_503), .B(n_451), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_485), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_482), .B(n_455), .Y(n_525) );
INVx2_ASAP7_75t_SL g526 ( .A(n_488), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_500), .A2(n_455), .B1(n_469), .B2(n_470), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_491), .B(n_469), .Y(n_528) );
NOR2xp33_ASAP7_75t_R g529 ( .A(n_484), .B(n_446), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_485), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_488), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_500), .A2(n_469), .B1(n_470), .B2(n_439), .Y(n_532) );
INVx5_ASAP7_75t_L g533 ( .A(n_496), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_511), .B(n_469), .Y(n_534) );
INVx3_ASAP7_75t_L g535 ( .A(n_485), .Y(n_535) );
INVx3_ASAP7_75t_L g536 ( .A(n_499), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_472), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_513), .B(n_469), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_492), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_507), .B(n_439), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_475), .A2(n_465), .B1(n_388), .B2(n_462), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_472), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_499), .B(n_461), .Y(n_543) );
NOR2xp33_ASAP7_75t_R g544 ( .A(n_505), .B(n_334), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_499), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_505), .A2(n_465), .B1(n_464), .B2(n_462), .Y(n_546) );
INVx3_ASAP7_75t_L g547 ( .A(n_502), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_502), .Y(n_548) );
AND2x4_ASAP7_75t_L g549 ( .A(n_479), .B(n_464), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_502), .B(n_435), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_L g551 ( .A1(n_508), .A2(n_467), .B(n_321), .C(n_440), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_486), .Y(n_552) );
NAND3xp33_ASAP7_75t_L g553 ( .A(n_502), .B(n_316), .C(n_286), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_515), .B(n_467), .Y(n_554) );
BUFx3_ASAP7_75t_L g555 ( .A(n_505), .Y(n_555) );
INVx2_ASAP7_75t_SL g556 ( .A(n_505), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_515), .B(n_435), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_496), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_486), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_489), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_515), .B(n_304), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_477), .B(n_299), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_508), .B(n_386), .Y(n_563) );
BUFx2_ASAP7_75t_L g564 ( .A(n_496), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_483), .B(n_330), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_493), .Y(n_566) );
AND2x4_ASAP7_75t_SL g567 ( .A(n_478), .B(n_386), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_478), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_512), .B(n_307), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_478), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_512), .A2(n_514), .B1(n_496), .B2(n_495), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_514), .B(n_311), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_487), .B(n_496), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_496), .Y(n_574) );
A2O1A1Ixp33_ASAP7_75t_L g575 ( .A1(n_498), .A2(n_453), .B(n_440), .C(n_447), .Y(n_575) );
NOR2xp33_ASAP7_75t_R g576 ( .A(n_496), .B(n_344), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_480), .B(n_448), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_481), .B(n_330), .Y(n_578) );
BUFx4f_ASAP7_75t_L g579 ( .A(n_516), .Y(n_579) );
NOR2x2_ASAP7_75t_L g580 ( .A(n_501), .B(n_364), .Y(n_580) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_474), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_474), .B(n_371), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_494), .A2(n_424), .B1(n_327), .B2(n_340), .Y(n_583) );
BUFx12f_ASAP7_75t_L g584 ( .A(n_473), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_494), .B(n_383), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_504), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_504), .A2(n_383), .B1(n_406), .B2(n_403), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_509), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_509), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_473), .B(n_371), .Y(n_590) );
CKINVDCx8_ASAP7_75t_R g591 ( .A(n_473), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_510), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_510), .Y(n_593) );
INVx1_ASAP7_75t_SL g594 ( .A(n_510), .Y(n_594) );
NAND2xp33_ASAP7_75t_L g595 ( .A(n_473), .B(n_429), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_473), .Y(n_596) );
BUFx2_ASAP7_75t_L g597 ( .A(n_544), .Y(n_597) );
INVxp67_ASAP7_75t_L g598 ( .A(n_526), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_524), .Y(n_599) );
A2O1A1Ixp33_ASAP7_75t_L g600 ( .A1(n_539), .A2(n_453), .B(n_333), .C(n_354), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_555), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_530), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_525), .A2(n_406), .B1(n_416), .B2(n_403), .Y(n_603) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_591), .Y(n_604) );
BUFx3_ASAP7_75t_L g605 ( .A(n_588), .Y(n_605) );
INVx4_ASAP7_75t_L g606 ( .A(n_555), .Y(n_606) );
INVx3_ASAP7_75t_L g607 ( .A(n_535), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_539), .A2(n_364), .B1(n_402), .B2(n_282), .Y(n_608) );
O2A1O1Ixp33_ASAP7_75t_L g609 ( .A1(n_531), .A2(n_351), .B(n_356), .C(n_355), .Y(n_609) );
INVx2_ASAP7_75t_SL g610 ( .A(n_567), .Y(n_610) );
AND2x4_ASAP7_75t_L g611 ( .A(n_522), .B(n_382), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_540), .B(n_377), .Y(n_612) );
AND2x4_ASAP7_75t_L g613 ( .A(n_522), .B(n_385), .Y(n_613) );
INVxp67_ASAP7_75t_L g614 ( .A(n_563), .Y(n_614) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_529), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_546), .B(n_377), .Y(n_616) );
INVx2_ASAP7_75t_SL g617 ( .A(n_567), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_523), .B(n_381), .Y(n_618) );
OAI221xp5_ASAP7_75t_L g619 ( .A1(n_541), .A2(n_323), .B1(n_398), .B2(n_399), .C(n_390), .Y(n_619) );
BUFx12f_ASAP7_75t_L g620 ( .A(n_549), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g621 ( .A1(n_551), .A2(n_408), .B(n_417), .C(n_413), .Y(n_621) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_533), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_545), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_548), .Y(n_624) );
A2O1A1Ixp33_ASAP7_75t_L g625 ( .A1(n_518), .A2(n_453), .B(n_431), .C(n_420), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_577), .B(n_402), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_568), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_520), .A2(n_447), .B1(n_452), .B2(n_437), .Y(n_628) );
BUFx2_ASAP7_75t_L g629 ( .A(n_576), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_L g630 ( .A1(n_518), .A2(n_456), .B(n_459), .C(n_452), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_573), .A2(n_359), .B(n_329), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_554), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_543), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_527), .A2(n_459), .B1(n_456), .B2(n_336), .Y(n_634) );
AO21x2_ASAP7_75t_L g635 ( .A1(n_575), .A2(n_314), .B(n_312), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_570), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_535), .Y(n_637) );
A2O1A1Ixp33_ASAP7_75t_L g638 ( .A1(n_528), .A2(n_317), .B(n_320), .C(n_319), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_520), .B(n_381), .Y(n_639) );
INVx3_ASAP7_75t_L g640 ( .A(n_536), .Y(n_640) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_576), .Y(n_641) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_533), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_519), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_549), .B(n_393), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_521), .B(n_393), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_556), .B(n_394), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_536), .Y(n_647) );
BUFx5_ASAP7_75t_L g648 ( .A(n_584), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_537), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_532), .B(n_394), .Y(n_650) );
BUFx2_ASAP7_75t_L g651 ( .A(n_529), .Y(n_651) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_533), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_533), .B(n_410), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_547), .Y(n_654) );
INVx3_ASAP7_75t_L g655 ( .A(n_547), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_587), .B(n_410), .Y(n_656) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_564), .Y(n_657) );
OR2x6_ASAP7_75t_L g658 ( .A(n_558), .B(n_324), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_542), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_552), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_559), .Y(n_661) );
CKINVDCx6p67_ASAP7_75t_R g662 ( .A(n_582), .Y(n_662) );
INVx1_ASAP7_75t_SL g663 ( .A(n_586), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_571), .A2(n_342), .B1(n_349), .B2(n_302), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_571), .A2(n_332), .B1(n_339), .B2(n_328), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_583), .Y(n_666) );
OAI221xp5_ASAP7_75t_L g667 ( .A1(n_553), .A2(n_395), .B1(n_373), .B2(n_350), .C(n_341), .Y(n_667) );
BUFx2_ASAP7_75t_L g668 ( .A(n_517), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_561), .A2(n_346), .B(n_345), .Y(n_669) );
NOR2xp33_ASAP7_75t_R g670 ( .A(n_595), .B(n_411), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_578), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_569), .A2(n_360), .B1(n_365), .B2(n_348), .Y(n_672) );
BUFx12f_ASAP7_75t_L g673 ( .A(n_517), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_580), .Y(n_674) );
OAI21xp33_ASAP7_75t_L g675 ( .A1(n_585), .A2(n_367), .B(n_366), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_560), .Y(n_676) );
BUFx8_ASAP7_75t_SL g677 ( .A(n_580), .Y(n_677) );
INVx4_ASAP7_75t_L g678 ( .A(n_579), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_585), .B(n_425), .Y(n_679) );
OAI22xp33_ASAP7_75t_L g680 ( .A1(n_558), .A2(n_425), .B1(n_313), .B2(n_325), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_561), .A2(n_374), .B(n_368), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_562), .B(n_289), .Y(n_682) );
INVx5_ASAP7_75t_L g683 ( .A(n_581), .Y(n_683) );
AOI222xp33_ASAP7_75t_L g684 ( .A1(n_569), .A2(n_392), .B1(n_426), .B2(n_423), .C1(n_421), .C2(n_430), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_565), .B(n_353), .Y(n_685) );
INVx4_ASAP7_75t_L g686 ( .A(n_579), .Y(n_686) );
INVx2_ASAP7_75t_SL g687 ( .A(n_572), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_566), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_574), .A2(n_375), .B1(n_379), .B2(n_376), .Y(n_689) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_581), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_574), .A2(n_538), .B1(n_534), .B2(n_572), .Y(n_691) );
AND2x4_ASAP7_75t_L g692 ( .A(n_550), .B(n_384), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_557), .B(n_357), .Y(n_693) );
NAND2xp33_ASAP7_75t_L g694 ( .A(n_581), .B(n_396), .Y(n_694) );
BUFx12f_ASAP7_75t_L g695 ( .A(n_581), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_589), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_575), .A2(n_391), .B1(n_397), .B2(n_389), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_590), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_593), .B(n_401), .Y(n_699) );
BUFx6f_ASAP7_75t_L g700 ( .A(n_592), .Y(n_700) );
A2O1A1Ixp33_ASAP7_75t_L g701 ( .A1(n_594), .A2(n_405), .B(n_407), .C(n_404), .Y(n_701) );
OAI221xp5_ASAP7_75t_L g702 ( .A1(n_596), .A2(n_418), .B1(n_428), .B2(n_415), .C(n_412), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_525), .B(n_409), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_546), .A2(n_380), .B1(n_400), .B2(n_363), .Y(n_704) );
BUFx2_ASAP7_75t_L g705 ( .A(n_544), .Y(n_705) );
INVxp67_ASAP7_75t_L g706 ( .A(n_526), .Y(n_706) );
BUFx6f_ASAP7_75t_L g707 ( .A(n_591), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_554), .Y(n_708) );
BUFx3_ASAP7_75t_L g709 ( .A(n_588), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_525), .B(n_370), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_529), .Y(n_711) );
AND2x4_ASAP7_75t_L g712 ( .A(n_522), .B(n_372), .Y(n_712) );
INVx4_ASAP7_75t_L g713 ( .A(n_555), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_524), .Y(n_714) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_544), .Y(n_715) );
INVx4_ASAP7_75t_L g716 ( .A(n_555), .Y(n_716) );
OAI21x1_ASAP7_75t_L g717 ( .A1(n_697), .A2(n_400), .B(n_380), .Y(n_717) );
BUFx2_ASAP7_75t_L g718 ( .A(n_648), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_625), .A2(n_422), .B(n_343), .Y(n_719) );
AO21x2_ASAP7_75t_L g720 ( .A1(n_635), .A2(n_422), .B(n_450), .Y(n_720) );
OAI21x1_ASAP7_75t_L g721 ( .A1(n_698), .A2(n_458), .B(n_450), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_611), .Y(n_722) );
NAND2xp33_ASAP7_75t_R g723 ( .A(n_615), .B(n_4), .Y(n_723) );
OR2x2_ASAP7_75t_L g724 ( .A(n_608), .B(n_5), .Y(n_724) );
OA21x2_ASAP7_75t_L g725 ( .A1(n_600), .A2(n_463), .B(n_458), .Y(n_725) );
INVx4_ASAP7_75t_L g726 ( .A(n_648), .Y(n_726) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_604), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_633), .A2(n_419), .B1(n_463), .B2(n_427), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_660), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_630), .A2(n_463), .B(n_490), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_611), .Y(n_731) );
OAI21x1_ASAP7_75t_L g732 ( .A1(n_661), .A2(n_362), .B(n_315), .Y(n_732) );
NOR3xp33_ASAP7_75t_L g733 ( .A(n_619), .B(n_378), .C(n_5), .Y(n_733) );
NAND2x1p5_ASAP7_75t_L g734 ( .A(n_604), .B(n_315), .Y(n_734) );
INVxp67_ASAP7_75t_SL g735 ( .A(n_604), .Y(n_735) );
AO31x2_ASAP7_75t_L g736 ( .A1(n_704), .A2(n_457), .A3(n_468), .B(n_362), .Y(n_736) );
OAI21x1_ASAP7_75t_L g737 ( .A1(n_649), .A2(n_362), .B(n_457), .Y(n_737) );
BUFx3_ASAP7_75t_L g738 ( .A(n_648), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_635), .A2(n_510), .B(n_490), .Y(n_739) );
INVx4_ASAP7_75t_SL g740 ( .A(n_707), .Y(n_740) );
OAI21x1_ASAP7_75t_L g741 ( .A1(n_659), .A2(n_468), .B(n_457), .Y(n_741) );
NOR2x1_ASAP7_75t_SL g742 ( .A(n_658), .B(n_444), .Y(n_742) );
OAI22xp33_ASAP7_75t_L g743 ( .A1(n_668), .A2(n_444), .B1(n_468), .B2(n_8), .Y(n_743) );
OAI21x1_ASAP7_75t_L g744 ( .A1(n_676), .A2(n_468), .B(n_490), .Y(n_744) );
OAI21x1_ASAP7_75t_L g745 ( .A1(n_688), .A2(n_468), .B(n_490), .Y(n_745) );
BUFx5_ASAP7_75t_L g746 ( .A(n_695), .Y(n_746) );
BUFx8_ASAP7_75t_L g747 ( .A(n_651), .Y(n_747) );
O2A1O1Ixp33_ASAP7_75t_SL g748 ( .A1(n_638), .A2(n_99), .B(n_100), .C(n_89), .Y(n_748) );
AND2x2_ASAP7_75t_SL g749 ( .A(n_597), .B(n_705), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g750 ( .A1(n_691), .A2(n_510), .B(n_444), .Y(n_750) );
OAI21x1_ASAP7_75t_L g751 ( .A1(n_669), .A2(n_107), .B(n_105), .Y(n_751) );
NAND3xp33_ASAP7_75t_SL g752 ( .A(n_663), .B(n_6), .C(n_7), .Y(n_752) );
OR2x6_ASAP7_75t_L g753 ( .A(n_673), .B(n_610), .Y(n_753) );
OR2x2_ASAP7_75t_L g754 ( .A(n_608), .B(n_7), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_626), .B(n_9), .Y(n_755) );
OAI21x1_ASAP7_75t_L g756 ( .A1(n_681), .A2(n_111), .B(n_108), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_613), .Y(n_757) );
A2O1A1Ixp33_ASAP7_75t_L g758 ( .A1(n_675), .A2(n_10), .B(n_12), .C(n_14), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_675), .A2(n_115), .B(n_112), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_599), .Y(n_760) );
AO21x2_ASAP7_75t_L g761 ( .A1(n_701), .A2(n_119), .B(n_117), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_602), .Y(n_762) );
NOR2x1_ASAP7_75t_L g763 ( .A(n_711), .B(n_14), .Y(n_763) );
OAI21x1_ASAP7_75t_L g764 ( .A1(n_627), .A2(n_125), .B(n_123), .Y(n_764) );
INVx3_ASAP7_75t_L g765 ( .A(n_648), .Y(n_765) );
BUFx6f_ASAP7_75t_L g766 ( .A(n_707), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g767 ( .A(n_677), .Y(n_767) );
O2A1O1Ixp33_ASAP7_75t_L g768 ( .A1(n_634), .A2(n_15), .B(n_17), .C(n_18), .Y(n_768) );
NAND2x1p5_ASAP7_75t_L g769 ( .A(n_707), .B(n_15), .Y(n_769) );
AO21x2_ASAP7_75t_L g770 ( .A1(n_704), .A2(n_130), .B(n_126), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_631), .A2(n_135), .B(n_131), .Y(n_771) );
OAI21xp5_ASAP7_75t_L g772 ( .A1(n_643), .A2(n_20), .B(n_21), .Y(n_772) );
OAI21x1_ASAP7_75t_L g773 ( .A1(n_636), .A2(n_137), .B(n_136), .Y(n_773) );
BUFx2_ASAP7_75t_L g774 ( .A(n_605), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_709), .Y(n_775) );
INVx2_ASAP7_75t_SL g776 ( .A(n_617), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_674), .A2(n_22), .B1(n_23), .B2(n_25), .Y(n_777) );
OR2x6_ASAP7_75t_SL g778 ( .A(n_666), .B(n_25), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_665), .A2(n_26), .B1(n_27), .B2(n_28), .Y(n_779) );
BUFx2_ASAP7_75t_L g780 ( .A(n_620), .Y(n_780) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_690), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_692), .A2(n_28), .B1(n_29), .B2(n_30), .Y(n_782) );
NOR2x1_ASAP7_75t_SL g783 ( .A(n_658), .B(n_29), .Y(n_783) );
OAI21xp5_ASAP7_75t_L g784 ( .A1(n_664), .A2(n_31), .B(n_32), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_712), .Y(n_785) );
OAI21x1_ASAP7_75t_L g786 ( .A1(n_696), .A2(n_139), .B(n_138), .Y(n_786) );
BUFx6f_ASAP7_75t_L g787 ( .A(n_690), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_623), .Y(n_788) );
OR2x2_ASAP7_75t_L g789 ( .A(n_603), .B(n_34), .Y(n_789) );
NAND2x1p5_ASAP7_75t_L g790 ( .A(n_606), .B(n_34), .Y(n_790) );
BUFx2_ASAP7_75t_L g791 ( .A(n_715), .Y(n_791) );
INVx4_ASAP7_75t_L g792 ( .A(n_606), .Y(n_792) );
OAI21x1_ASAP7_75t_L g793 ( .A1(n_653), .A2(n_141), .B(n_140), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_624), .Y(n_794) );
NAND2xp5_ASAP7_75t_SL g795 ( .A(n_601), .B(n_35), .Y(n_795) );
INVx4_ASAP7_75t_L g796 ( .A(n_713), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_714), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_614), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_632), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_708), .Y(n_800) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_601), .Y(n_801) );
AO32x2_ASAP7_75t_L g802 ( .A1(n_689), .A2(n_36), .A3(n_37), .B1(n_39), .B2(n_40), .Y(n_802) );
AO21x2_ASAP7_75t_L g803 ( .A1(n_670), .A2(n_146), .B(n_143), .Y(n_803) );
OR2x2_ASAP7_75t_L g804 ( .A(n_603), .B(n_36), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_703), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_703), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g807 ( .A1(n_671), .A2(n_37), .B1(n_39), .B2(n_40), .Y(n_807) );
OR2x2_ASAP7_75t_L g808 ( .A(n_644), .B(n_41), .Y(n_808) );
AND2x4_ASAP7_75t_L g809 ( .A(n_678), .B(n_42), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_612), .B(n_42), .Y(n_810) );
BUFx3_ASAP7_75t_L g811 ( .A(n_713), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_639), .Y(n_812) );
NOR2x1_ASAP7_75t_SL g813 ( .A(n_658), .B(n_43), .Y(n_813) );
AND2x2_ASAP7_75t_L g814 ( .A(n_710), .B(n_43), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_598), .Y(n_815) );
A2O1A1Ixp33_ASAP7_75t_L g816 ( .A1(n_609), .A2(n_44), .B(n_45), .C(n_46), .Y(n_816) );
OAI21x1_ASAP7_75t_SL g817 ( .A1(n_646), .A2(n_45), .B(n_47), .Y(n_817) );
INVx5_ASAP7_75t_L g818 ( .A(n_716), .Y(n_818) );
AO21x2_ASAP7_75t_L g819 ( .A1(n_692), .A2(n_184), .B(n_281), .Y(n_819) );
OA21x2_ASAP7_75t_L g820 ( .A1(n_702), .A2(n_182), .B(n_279), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_644), .Y(n_821) );
OAI21x1_ASAP7_75t_L g822 ( .A1(n_689), .A2(n_179), .B(n_278), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_706), .B(n_48), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_628), .Y(n_824) );
BUFx6f_ASAP7_75t_L g825 ( .A(n_690), .Y(n_825) );
AOI22xp33_ASAP7_75t_SL g826 ( .A1(n_629), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_637), .Y(n_827) );
INVx4_ASAP7_75t_L g828 ( .A(n_678), .Y(n_828) );
OAI21x1_ASAP7_75t_L g829 ( .A1(n_607), .A2(n_192), .B(n_277), .Y(n_829) );
OAI21x1_ASAP7_75t_L g830 ( .A1(n_607), .A2(n_191), .B(n_276), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_647), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_654), .Y(n_832) );
OAI21x1_ASAP7_75t_L g833 ( .A1(n_640), .A2(n_178), .B(n_272), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_621), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_640), .Y(n_835) );
BUFx6f_ASAP7_75t_L g836 ( .A(n_622), .Y(n_836) );
OAI21x1_ASAP7_75t_L g837 ( .A1(n_655), .A2(n_177), .B(n_271), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_684), .A2(n_52), .B1(n_53), .B2(n_54), .Y(n_838) );
OAI21x1_ASAP7_75t_L g839 ( .A1(n_655), .A2(n_194), .B(n_270), .Y(n_839) );
OAI21x1_ASAP7_75t_L g840 ( .A1(n_699), .A2(n_193), .B(n_266), .Y(n_840) );
AOI221xp5_ASAP7_75t_L g841 ( .A1(n_667), .A2(n_55), .B1(n_56), .B2(n_57), .C(n_58), .Y(n_841) );
AND2x4_ASAP7_75t_L g842 ( .A(n_686), .B(n_55), .Y(n_842) );
INVx3_ASAP7_75t_L g843 ( .A(n_657), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_687), .Y(n_844) );
AO21x2_ASAP7_75t_L g845 ( .A1(n_739), .A2(n_679), .B(n_650), .Y(n_845) );
AOI21xp5_ASAP7_75t_L g846 ( .A1(n_739), .A2(n_646), .B(n_694), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_733), .A2(n_662), .B1(n_684), .B2(n_641), .Y(n_847) );
AOI221xp5_ASAP7_75t_L g848 ( .A1(n_805), .A2(n_656), .B1(n_616), .B2(n_672), .C(n_618), .Y(n_848) );
AOI22xp33_ASAP7_75t_SL g849 ( .A1(n_783), .A2(n_686), .B1(n_645), .B2(n_657), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_724), .B(n_682), .Y(n_850) );
OAI221xp5_ASAP7_75t_L g851 ( .A1(n_755), .A2(n_685), .B1(n_693), .B2(n_657), .C(n_683), .Y(n_851) );
OAI22xp33_ASAP7_75t_L g852 ( .A1(n_754), .A2(n_838), .B1(n_804), .B2(n_789), .Y(n_852) );
AND2x2_ASAP7_75t_L g853 ( .A(n_806), .B(n_56), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_733), .A2(n_680), .B1(n_652), .B2(n_642), .Y(n_854) );
AOI22xp33_ASAP7_75t_SL g855 ( .A1(n_813), .A2(n_683), .B1(n_642), .B2(n_652), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_838), .A2(n_683), .B1(n_652), .B2(n_642), .Y(n_856) );
OAI22xp33_ASAP7_75t_L g857 ( .A1(n_807), .A2(n_622), .B1(n_700), .B2(n_59), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_834), .B(n_622), .Y(n_858) );
AND2x4_ASAP7_75t_L g859 ( .A(n_726), .B(n_57), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_808), .A2(n_61), .B1(n_63), .B2(n_64), .Y(n_860) );
INVxp67_ASAP7_75t_L g861 ( .A(n_801), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_821), .A2(n_63), .B1(n_64), .B2(n_65), .Y(n_862) );
OAI211xp5_ASAP7_75t_L g863 ( .A1(n_807), .A2(n_66), .B(n_67), .C(n_68), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_790), .A2(n_71), .B1(n_72), .B2(n_73), .Y(n_864) );
OA21x2_ASAP7_75t_L g865 ( .A1(n_750), .A2(n_206), .B(n_265), .Y(n_865) );
OA21x2_ASAP7_75t_L g866 ( .A1(n_750), .A2(n_719), .B(n_732), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_760), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_798), .B(n_74), .Y(n_868) );
OAI221xp5_ASAP7_75t_L g869 ( .A1(n_823), .A2(n_76), .B1(n_77), .B2(n_78), .C(n_79), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_762), .Y(n_870) );
AO31x2_ASAP7_75t_L g871 ( .A1(n_730), .A2(n_150), .A3(n_152), .B(n_153), .Y(n_871) );
AOI21xp5_ASAP7_75t_L g872 ( .A1(n_730), .A2(n_159), .B(n_160), .Y(n_872) );
AOI221xp5_ASAP7_75t_L g873 ( .A1(n_768), .A2(n_162), .B1(n_167), .B2(n_168), .C(n_170), .Y(n_873) );
AOI21x1_ASAP7_75t_L g874 ( .A1(n_725), .A2(n_171), .B(n_173), .Y(n_874) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_818), .Y(n_875) );
BUFx2_ASAP7_75t_L g876 ( .A(n_746), .Y(n_876) );
OAI21x1_ASAP7_75t_L g877 ( .A1(n_744), .A2(n_197), .B(n_198), .Y(n_877) );
AOI221xp5_ASAP7_75t_L g878 ( .A1(n_784), .A2(n_841), .B1(n_779), .B2(n_743), .C(n_722), .Y(n_878) );
AND2x2_ASAP7_75t_L g879 ( .A(n_778), .B(n_200), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_790), .A2(n_201), .B1(n_204), .B2(n_205), .Y(n_880) );
AOI21xp33_ASAP7_75t_L g881 ( .A1(n_728), .A2(n_810), .B(n_824), .Y(n_881) );
OAI221xp5_ASAP7_75t_L g882 ( .A1(n_731), .A2(n_220), .B1(n_221), .B2(n_226), .C(n_228), .Y(n_882) );
HB1xp67_ASAP7_75t_L g883 ( .A(n_818), .Y(n_883) );
BUFx2_ASAP7_75t_L g884 ( .A(n_746), .Y(n_884) );
AOI222xp33_ASAP7_75t_L g885 ( .A1(n_784), .A2(n_231), .B1(n_232), .B2(n_233), .C1(n_235), .C2(n_237), .Y(n_885) );
AOI222xp33_ASAP7_75t_L g886 ( .A1(n_757), .A2(n_250), .B1(n_253), .B2(n_254), .C1(n_255), .C2(n_258), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_788), .Y(n_887) );
AOI22xp33_ASAP7_75t_SL g888 ( .A1(n_772), .A2(n_259), .B1(n_261), .B2(n_262), .Y(n_888) );
INVx2_ASAP7_75t_L g889 ( .A(n_794), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_814), .B(n_749), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_812), .B(n_799), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_815), .B(n_774), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_800), .B(n_785), .Y(n_893) );
HB1xp67_ASAP7_75t_L g894 ( .A(n_818), .Y(n_894) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_818), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_797), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_809), .A2(n_842), .B1(n_791), .B2(n_753), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_753), .A2(n_795), .B1(n_747), .B2(n_780), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_802), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_802), .Y(n_900) );
OR2x6_ASAP7_75t_L g901 ( .A(n_726), .B(n_753), .Y(n_901) );
OAI22xp33_ASAP7_75t_L g902 ( .A1(n_723), .A2(n_743), .B1(n_718), .B2(n_752), .Y(n_902) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_817), .A2(n_742), .B1(n_769), .B2(n_820), .Y(n_903) );
AND2x4_ASAP7_75t_L g904 ( .A(n_738), .B(n_765), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_747), .A2(n_826), .B1(n_782), .B2(n_763), .Y(n_905) );
INVx2_ASAP7_75t_SL g906 ( .A(n_746), .Y(n_906) );
INVx2_ASAP7_75t_L g907 ( .A(n_827), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_802), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_811), .B(n_746), .Y(n_909) );
AOI21xp5_ASAP7_75t_L g910 ( .A1(n_725), .A2(n_745), .B(n_720), .Y(n_910) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_826), .A2(n_769), .B1(n_796), .B2(n_792), .Y(n_911) );
INVx3_ASAP7_75t_L g912 ( .A(n_765), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_844), .Y(n_913) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_775), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_831), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_832), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_777), .A2(n_792), .B1(n_796), .B2(n_776), .Y(n_917) );
OAI21xp33_ASAP7_75t_L g918 ( .A1(n_816), .A2(n_758), .B(n_717), .Y(n_918) );
INVx2_ASAP7_75t_L g919 ( .A(n_736), .Y(n_919) );
AOI22xp33_ASAP7_75t_SL g920 ( .A1(n_820), .A2(n_770), .B1(n_819), .B2(n_803), .Y(n_920) );
INVx1_ASAP7_75t_SL g921 ( .A(n_727), .Y(n_921) );
NAND4xp25_ASAP7_75t_L g922 ( .A(n_828), .B(n_771), .C(n_759), .D(n_835), .Y(n_922) );
AND2x4_ASAP7_75t_L g923 ( .A(n_740), .B(n_766), .Y(n_923) );
AOI221xp5_ASAP7_75t_L g924 ( .A1(n_767), .A2(n_748), .B1(n_771), .B2(n_759), .C(n_735), .Y(n_924) );
AOI21xp5_ASAP7_75t_L g925 ( .A1(n_720), .A2(n_741), .B(n_737), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_736), .Y(n_926) );
OAI22xp33_ASAP7_75t_L g927 ( .A1(n_734), .A2(n_843), .B1(n_836), .B2(n_825), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_819), .A2(n_761), .B1(n_803), .B2(n_740), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_740), .B(n_836), .Y(n_929) );
OAI21xp33_ASAP7_75t_L g930 ( .A1(n_822), .A2(n_840), .B(n_721), .Y(n_930) );
A2O1A1Ixp33_ASAP7_75t_L g931 ( .A1(n_751), .A2(n_756), .B(n_793), .C(n_837), .Y(n_931) );
AOI211xp5_ASAP7_75t_L g932 ( .A1(n_829), .A2(n_839), .B(n_833), .C(n_830), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_781), .B(n_825), .Y(n_933) );
AO21x2_ASAP7_75t_L g934 ( .A1(n_764), .A2(n_773), .B(n_786), .Y(n_934) );
NAND3xp33_ASAP7_75t_L g935 ( .A(n_781), .B(n_787), .C(n_825), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_781), .Y(n_936) );
AO21x2_ASAP7_75t_L g937 ( .A1(n_787), .A2(n_739), .B(n_750), .Y(n_937) );
INVx2_ASAP7_75t_L g938 ( .A(n_729), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_733), .A2(n_674), .B1(n_673), .B2(n_668), .Y(n_939) );
OAI21x1_ASAP7_75t_SL g940 ( .A1(n_742), .A2(n_813), .B(n_783), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_724), .B(n_503), .Y(n_941) );
OAI22xp33_ASAP7_75t_L g942 ( .A1(n_724), .A2(n_608), .B1(n_497), .B2(n_754), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_724), .B(n_503), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_942), .B(n_941), .Y(n_944) );
HB1xp67_ASAP7_75t_L g945 ( .A(n_875), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_899), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_943), .B(n_852), .Y(n_947) );
OR2x2_ASAP7_75t_L g948 ( .A(n_861), .B(n_921), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_900), .Y(n_949) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_875), .Y(n_950) );
AND2x2_ASAP7_75t_L g951 ( .A(n_938), .B(n_867), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_908), .Y(n_952) );
INVx2_ASAP7_75t_SL g953 ( .A(n_883), .Y(n_953) );
INVx3_ASAP7_75t_L g954 ( .A(n_923), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_858), .Y(n_955) );
BUFx3_ASAP7_75t_L g956 ( .A(n_876), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_926), .Y(n_957) );
BUFx3_ASAP7_75t_L g958 ( .A(n_884), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_870), .B(n_887), .Y(n_959) );
HB1xp67_ASAP7_75t_L g960 ( .A(n_894), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_850), .B(n_939), .Y(n_961) );
BUFx2_ASAP7_75t_SL g962 ( .A(n_859), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_889), .B(n_896), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_919), .Y(n_964) );
AND2x2_ASAP7_75t_L g965 ( .A(n_907), .B(n_915), .Y(n_965) );
INVx2_ASAP7_75t_L g966 ( .A(n_937), .Y(n_966) );
INVx2_ASAP7_75t_L g967 ( .A(n_937), .Y(n_967) );
HB1xp67_ASAP7_75t_L g968 ( .A(n_895), .Y(n_968) );
AND2x4_ASAP7_75t_L g969 ( .A(n_895), .B(n_923), .Y(n_969) );
HB1xp67_ASAP7_75t_L g970 ( .A(n_909), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_891), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_871), .Y(n_972) );
INVx2_ASAP7_75t_L g973 ( .A(n_866), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_916), .B(n_853), .Y(n_974) );
BUFx5_ASAP7_75t_L g975 ( .A(n_936), .Y(n_975) );
OA21x2_ASAP7_75t_L g976 ( .A1(n_910), .A2(n_925), .B(n_924), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_845), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_845), .Y(n_978) );
INVx2_ASAP7_75t_L g979 ( .A(n_865), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_893), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_861), .Y(n_981) );
OAI22xp5_ASAP7_75t_L g982 ( .A1(n_905), .A2(n_897), .B1(n_854), .B2(n_847), .Y(n_982) );
INVx4_ASAP7_75t_SL g983 ( .A(n_901), .Y(n_983) );
INVx2_ASAP7_75t_L g984 ( .A(n_865), .Y(n_984) );
OAI222xp33_ASAP7_75t_L g985 ( .A1(n_902), .A2(n_901), .B1(n_911), .B2(n_879), .C1(n_864), .C2(n_849), .Y(n_985) );
NAND2x1_ASAP7_75t_L g986 ( .A(n_940), .B(n_928), .Y(n_986) );
BUFx6f_ASAP7_75t_L g987 ( .A(n_933), .Y(n_987) );
NAND2xp5_ASAP7_75t_SL g988 ( .A(n_855), .B(n_849), .Y(n_988) );
AND2x4_ASAP7_75t_L g989 ( .A(n_912), .B(n_935), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_874), .Y(n_990) );
INVx3_ASAP7_75t_L g991 ( .A(n_901), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_890), .B(n_848), .Y(n_992) );
INVx3_ASAP7_75t_L g993 ( .A(n_904), .Y(n_993) );
INVx2_ASAP7_75t_L g994 ( .A(n_877), .Y(n_994) );
HB1xp67_ASAP7_75t_L g995 ( .A(n_906), .Y(n_995) );
INVx2_ASAP7_75t_L g996 ( .A(n_934), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_878), .B(n_881), .Y(n_997) );
HB1xp67_ASAP7_75t_L g998 ( .A(n_892), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_868), .B(n_898), .Y(n_999) );
INVx2_ASAP7_75t_L g1000 ( .A(n_913), .Y(n_1000) );
INVx2_ASAP7_75t_L g1001 ( .A(n_929), .Y(n_1001) );
INVx2_ASAP7_75t_L g1002 ( .A(n_856), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_885), .B(n_863), .Y(n_1003) );
AO21x2_ASAP7_75t_L g1004 ( .A1(n_910), .A2(n_925), .B(n_930), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_863), .B(n_855), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_846), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_862), .B(n_888), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_917), .B(n_860), .Y(n_1008) );
HB1xp67_ASAP7_75t_L g1009 ( .A(n_914), .Y(n_1009) );
NOR2x1_ASAP7_75t_L g1010 ( .A(n_922), .B(n_927), .Y(n_1010) );
NOR2xp33_ASAP7_75t_L g1011 ( .A(n_869), .B(n_857), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_888), .B(n_873), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_846), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_903), .Y(n_1014) );
INVx2_ASAP7_75t_L g1015 ( .A(n_880), .Y(n_1015) );
INVx2_ASAP7_75t_L g1016 ( .A(n_882), .Y(n_1016) );
BUFx2_ASAP7_75t_L g1017 ( .A(n_931), .Y(n_1017) );
BUFx3_ASAP7_75t_L g1018 ( .A(n_851), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_886), .B(n_920), .Y(n_1019) );
INVx2_ASAP7_75t_L g1020 ( .A(n_932), .Y(n_1020) );
NOR2x1_ASAP7_75t_SL g1021 ( .A(n_872), .B(n_918), .Y(n_1021) );
HB1xp67_ASAP7_75t_L g1022 ( .A(n_945), .Y(n_1022) );
HB1xp67_ASAP7_75t_L g1023 ( .A(n_950), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_957), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_946), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_946), .Y(n_1026) );
AND2x4_ASAP7_75t_L g1027 ( .A(n_983), .B(n_991), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_949), .Y(n_1028) );
INVx2_ASAP7_75t_L g1029 ( .A(n_973), .Y(n_1029) );
AOI221xp5_ASAP7_75t_L g1030 ( .A1(n_982), .A2(n_947), .B1(n_944), .B2(n_992), .C(n_985), .Y(n_1030) );
AND2x4_ASAP7_75t_L g1031 ( .A(n_983), .B(n_991), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_949), .B(n_952), .Y(n_1032) );
OR2x2_ASAP7_75t_L g1033 ( .A(n_953), .B(n_960), .Y(n_1033) );
OAI321xp33_ASAP7_75t_L g1034 ( .A1(n_988), .A2(n_1003), .A3(n_1005), .B1(n_1019), .B2(n_997), .C(n_1012), .Y(n_1034) );
INVx1_ASAP7_75t_SL g1035 ( .A(n_1009), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_964), .Y(n_1036) );
AND2x4_ASAP7_75t_L g1037 ( .A(n_983), .B(n_991), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_951), .B(n_959), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1000), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_964), .Y(n_1040) );
INVxp67_ASAP7_75t_L g1041 ( .A(n_968), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_955), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_963), .B(n_965), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_965), .B(n_955), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g1045 ( .A1(n_1003), .A2(n_1011), .B1(n_1019), .B2(n_1012), .Y(n_1045) );
INVx8_ASAP7_75t_L g1046 ( .A(n_969), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_974), .B(n_1014), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_981), .Y(n_1048) );
NOR2xp33_ASAP7_75t_L g1049 ( .A(n_998), .B(n_999), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_977), .Y(n_1050) );
BUFx6f_ASAP7_75t_L g1051 ( .A(n_987), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_971), .B(n_980), .Y(n_1052) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_970), .Y(n_1053) );
AND2x4_ASAP7_75t_L g1054 ( .A(n_956), .B(n_958), .Y(n_1054) );
AOI22xp5_ASAP7_75t_L g1055 ( .A1(n_1008), .A2(n_961), .B1(n_1007), .B2(n_962), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_1020), .B(n_1001), .Y(n_1056) );
HB1xp67_ASAP7_75t_L g1057 ( .A(n_948), .Y(n_1057) );
BUFx6f_ASAP7_75t_L g1058 ( .A(n_987), .Y(n_1058) );
INVx5_ASAP7_75t_L g1059 ( .A(n_969), .Y(n_1059) );
INVx4_ASAP7_75t_L g1060 ( .A(n_956), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_978), .Y(n_1061) );
AO21x2_ASAP7_75t_L g1062 ( .A1(n_990), .A2(n_972), .B(n_1006), .Y(n_1062) );
AND2x4_ASAP7_75t_L g1063 ( .A(n_969), .B(n_989), .Y(n_1063) );
INVx2_ASAP7_75t_L g1064 ( .A(n_1029), .Y(n_1064) );
NOR2xp33_ASAP7_75t_L g1065 ( .A(n_1035), .B(n_993), .Y(n_1065) );
AND2x4_ASAP7_75t_L g1066 ( .A(n_1063), .B(n_966), .Y(n_1066) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_1057), .B(n_966), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1047), .B(n_967), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_1030), .A2(n_1018), .B1(n_1016), .B2(n_1015), .Y(n_1069) );
NAND4xp25_ASAP7_75t_L g1070 ( .A(n_1045), .B(n_1018), .C(n_1010), .D(n_1017), .Y(n_1070) );
INVx2_ASAP7_75t_SL g1071 ( .A(n_1060), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1024), .Y(n_1072) );
NOR2xp33_ASAP7_75t_L g1073 ( .A(n_1049), .B(n_993), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1048), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_1038), .B(n_993), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1022), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1023), .Y(n_1077) );
HB1xp67_ASAP7_75t_L g1078 ( .A(n_1053), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1047), .B(n_967), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1032), .B(n_1017), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1032), .B(n_1006), .Y(n_1081) );
NOR2xp33_ASAP7_75t_SL g1082 ( .A(n_1060), .B(n_995), .Y(n_1082) );
AND2x4_ASAP7_75t_L g1083 ( .A(n_1063), .B(n_1013), .Y(n_1083) );
OR2x2_ASAP7_75t_L g1084 ( .A(n_1043), .B(n_976), .Y(n_1084) );
AND2x4_ASAP7_75t_L g1085 ( .A(n_1063), .B(n_986), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1025), .Y(n_1086) );
INVx2_ASAP7_75t_SL g1087 ( .A(n_1060), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1025), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_1026), .B(n_996), .Y(n_1089) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_1033), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1026), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_1044), .B(n_975), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1039), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1028), .B(n_1004), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1028), .Y(n_1095) );
XOR2xp5_ASAP7_75t_L g1096 ( .A(n_1070), .B(n_1055), .Y(n_1096) );
NOR2xp33_ASAP7_75t_L g1097 ( .A(n_1078), .B(n_1034), .Y(n_1097) );
OR2x6_ASAP7_75t_L g1098 ( .A(n_1085), .B(n_1046), .Y(n_1098) );
NOR2xp33_ASAP7_75t_L g1099 ( .A(n_1076), .B(n_1041), .Y(n_1099) );
INVx2_ASAP7_75t_L g1100 ( .A(n_1064), .Y(n_1100) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1064), .Y(n_1101) );
NAND2xp5_ASAP7_75t_SL g1102 ( .A(n_1082), .B(n_1054), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1090), .Y(n_1103) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_1084), .B(n_1061), .Y(n_1104) );
OR2x2_ASAP7_75t_L g1105 ( .A(n_1084), .B(n_1061), .Y(n_1105) );
NOR2xp33_ASAP7_75t_L g1106 ( .A(n_1077), .B(n_1052), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1072), .Y(n_1107) );
INVx1_ASAP7_75t_SL g1108 ( .A(n_1071), .Y(n_1108) );
OR2x2_ASAP7_75t_L g1109 ( .A(n_1067), .B(n_1050), .Y(n_1109) );
INVx1_ASAP7_75t_SL g1110 ( .A(n_1087), .Y(n_1110) );
OAI21xp5_ASAP7_75t_L g1111 ( .A1(n_1069), .A2(n_1016), .B(n_1042), .Y(n_1111) );
AOI22xp5_ASAP7_75t_L g1112 ( .A1(n_1073), .A2(n_1031), .B1(n_1037), .B2(n_1027), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1086), .Y(n_1113) );
AOI221x1_ASAP7_75t_L g1114 ( .A1(n_1097), .A2(n_1065), .B1(n_1074), .B2(n_1091), .C(n_1088), .Y(n_1114) );
INVxp67_ASAP7_75t_L g1115 ( .A(n_1108), .Y(n_1115) );
OAI22xp5_ASAP7_75t_L g1116 ( .A1(n_1096), .A2(n_1059), .B1(n_1092), .B2(n_1075), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1103), .B(n_1081), .Y(n_1117) );
INVx2_ASAP7_75t_L g1118 ( .A(n_1100), .Y(n_1118) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1100), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1113), .Y(n_1120) );
OAI321xp33_ASAP7_75t_L g1121 ( .A1(n_1102), .A2(n_1111), .A3(n_1112), .B1(n_1098), .B2(n_1104), .C(n_1105), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_1099), .A2(n_1083), .B1(n_1080), .B2(n_1085), .Y(n_1122) );
AOI22xp5_ASAP7_75t_L g1123 ( .A1(n_1106), .A2(n_1083), .B1(n_1066), .B2(n_1079), .Y(n_1123) );
AOI21xp5_ASAP7_75t_L g1124 ( .A1(n_1121), .A2(n_1098), .B(n_1110), .Y(n_1124) );
INVx2_ASAP7_75t_L g1125 ( .A(n_1118), .Y(n_1125) );
INVx2_ASAP7_75t_L g1126 ( .A(n_1118), .Y(n_1126) );
NOR2xp33_ASAP7_75t_L g1127 ( .A(n_1115), .B(n_1109), .Y(n_1127) );
XNOR2xp5_ASAP7_75t_L g1128 ( .A(n_1123), .B(n_1098), .Y(n_1128) );
AOI22xp5_ASAP7_75t_L g1129 ( .A1(n_1128), .A2(n_1122), .B1(n_1116), .B2(n_1117), .Y(n_1129) );
OAI211xp5_ASAP7_75t_SL g1130 ( .A1(n_1124), .A2(n_1120), .B(n_1109), .C(n_1107), .Y(n_1130) );
AOI22xp5_ASAP7_75t_L g1131 ( .A1(n_1127), .A2(n_1079), .B1(n_1068), .B2(n_1066), .Y(n_1131) );
A2O1A1Ixp33_ASAP7_75t_L g1132 ( .A1(n_1129), .A2(n_1125), .B(n_1126), .C(n_1027), .Y(n_1132) );
AOI221xp5_ASAP7_75t_L g1133 ( .A1(n_1130), .A2(n_1119), .B1(n_1095), .B2(n_1093), .C(n_1094), .Y(n_1133) );
NAND4xp75_ASAP7_75t_L g1134 ( .A(n_1133), .B(n_1114), .C(n_1131), .D(n_1056), .Y(n_1134) );
AOI21xp5_ASAP7_75t_L g1135 ( .A1(n_1132), .A2(n_1036), .B(n_1040), .Y(n_1135) );
NOR3xp33_ASAP7_75t_L g1136 ( .A(n_1134), .B(n_954), .C(n_1002), .Y(n_1136) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1135), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1137), .Y(n_1138) );
OAI22xp5_ASAP7_75t_SL g1139 ( .A1(n_1138), .A2(n_1136), .B1(n_989), .B2(n_984), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_1139), .B(n_1101), .Y(n_1140) );
OAI21xp5_ASAP7_75t_SL g1141 ( .A1(n_1140), .A2(n_1089), .B(n_994), .Y(n_1141) );
OAI22xp5_ASAP7_75t_SL g1142 ( .A1(n_1141), .A2(n_979), .B1(n_1051), .B2(n_1058), .Y(n_1142) );
AOI21xp5_ASAP7_75t_L g1143 ( .A1(n_1142), .A2(n_1021), .B(n_1062), .Y(n_1143) );
endmodule