module fake_jpeg_509_n_177 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_20),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_66),
.Y(n_71)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_68),
.Y(n_73)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_62),
.B(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_78),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_63),
.A2(n_52),
.B1(n_46),
.B2(n_50),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_75),
.A2(n_65),
.B1(n_46),
.B2(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_68),
.B(n_48),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_50),
.B1(n_59),
.B2(n_51),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_61),
.B1(n_53),
.B2(n_45),
.Y(n_97)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_80),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_81),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_79),
.A2(n_75),
.B1(n_68),
.B2(n_65),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_55),
.B1(n_60),
.B2(n_57),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_57),
.B1(n_55),
.B2(n_47),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_49),
.B1(n_47),
.B2(n_59),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_97),
.B1(n_70),
.B2(n_80),
.Y(n_98)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_96),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_94),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_49),
.B(n_53),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_73),
.B(n_45),
.C(n_4),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_1),
.B(n_2),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_73),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_2),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_102),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_61),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_106),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_72),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_115),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_72),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_40),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_113),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_80),
.B1(n_45),
.B2(n_5),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_36),
.B1(n_35),
.B2(n_34),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_39),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_45),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_87),
.C(n_37),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_3),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_3),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_32),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_86),
.B1(n_87),
.B2(n_6),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_118),
.B1(n_126),
.B2(n_129),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_106),
.A2(n_86),
.B1(n_87),
.B2(n_6),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_125),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_100),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_132),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_111),
.C(n_103),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_112),
.A2(n_4),
.B(n_5),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_12),
.B(n_13),
.Y(n_146)
);

XOR2x2_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_33),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_30),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_99),
.B1(n_109),
.B2(n_107),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_104),
.B1(n_10),
.B2(n_11),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_7),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_133),
.B(n_14),
.Y(n_148)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_130),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_138),
.B(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_146),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_119),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_128),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_14),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_129),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_153),
.A2(n_146),
.B(n_136),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_125),
.C(n_120),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_156),
.C(n_159),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_121),
.A3(n_120),
.B1(n_127),
.B2(n_122),
.C1(n_19),
.C2(n_20),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_15),
.C(n_16),
.Y(n_159)
);

INVxp67_ASAP7_75t_SL g160 ( 
.A(n_151),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_165),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_158),
.A2(n_147),
.B(n_144),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_162),
.C(n_164),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_141),
.B1(n_137),
.B2(n_145),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_137),
.B1(n_139),
.B2(n_17),
.Y(n_165)
);

AOI321xp33_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_154),
.A3(n_153),
.B1(n_159),
.B2(n_155),
.C(n_21),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_166),
.A2(n_160),
.B1(n_16),
.B2(n_17),
.Y(n_170)
);

NOR2xp67_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_168),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_169),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_15),
.B(n_18),
.C(n_22),
.Y(n_174)
);

OAI21x1_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_18),
.B(n_22),
.Y(n_175)
);

OAI21x1_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_23),
.B(n_24),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_23),
.Y(n_177)
);


endmodule