module fake_jpeg_7331_n_119 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_119);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_119;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_30),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_20),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_27),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_22),
.Y(n_44)
);

OA22x2_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_25),
.B1(n_12),
.B2(n_21),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_47),
.B1(n_13),
.B2(n_29),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_41),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_44),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_1),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_22),
.B1(n_23),
.B2(n_14),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_13),
.B1(n_16),
.B2(n_33),
.Y(n_49)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_58),
.B1(n_47),
.B2(n_46),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_39),
.C(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_54),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_46),
.B1(n_37),
.B2(n_29),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_24),
.C(n_20),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_57),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_33),
.B1(n_24),
.B2(n_16),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_37),
.B1(n_59),
.B2(n_33),
.Y(n_72)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_67),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

AND2x6_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_54),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_69),
.B(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_68),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_48),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_74),
.B1(n_66),
.B2(n_71),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_37),
.B1(n_59),
.B2(n_29),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_42),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_80),
.C(n_64),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_69),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_48),
.C(n_24),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_84),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

BUFx24_ASAP7_75t_SL g85 ( 
.A(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_80),
.C(n_73),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_88),
.B(n_89),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_90),
.A2(n_91),
.B(n_78),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_70),
.B(n_65),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_97),
.B(n_82),
.Y(n_101)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_81),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_95),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_97),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_74),
.B(n_76),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_98),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_61),
.B1(n_17),
.B2(n_4),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_106),
.Y(n_110)
);

OAI221xp5_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.C(n_94),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_93),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_2),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_100),
.B1(n_3),
.B2(n_5),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_112),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_114),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_116),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_110),
.B1(n_111),
.B2(n_107),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_8),
.B(n_9),
.C(n_114),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_8),
.Y(n_119)
);


endmodule