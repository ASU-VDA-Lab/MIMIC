module real_jpeg_2202_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_197;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_244;
wire n_128;
wire n_179;
wire n_167;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_2),
.A2(n_38),
.B1(n_55),
.B2(n_57),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_2),
.A2(n_38),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_38),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_46),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_3),
.A2(n_46),
.B1(n_55),
.B2(n_57),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_3),
.A2(n_46),
.B1(n_65),
.B2(n_66),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_46),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_3),
.B(n_55),
.C(n_70),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_3),
.B(n_72),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_3),
.B(n_36),
.C(n_52),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_3),
.B(n_26),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_3),
.B(n_40),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_3),
.B(n_25),
.C(n_41),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_3),
.B(n_50),
.Y(n_209)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_5),
.A2(n_28),
.B1(n_35),
.B2(n_36),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_5),
.A2(n_28),
.B1(n_55),
.B2(n_57),
.Y(n_245)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_10),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_233),
.B1(n_254),
.B2(n_255),
.Y(n_13)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_14),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_123),
.B(n_232),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_101),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_17),
.B(n_101),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_77),
.C(n_88),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_18),
.B(n_77),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_47),
.B2(n_48),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_19),
.B(n_49),
.C(n_76),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_21),
.A2(n_32),
.B1(n_33),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_21),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_22),
.B(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_23),
.B(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_23),
.A2(n_26),
.B1(n_93),
.B2(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_26),
.Y(n_23)
);

AO22x1_ASAP7_75t_L g40 ( 
.A1(n_24),
.A2(n_25),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_25),
.B(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_27),
.A2(n_29),
.B(n_92),
.Y(n_91)
);

OA21x2_ASAP7_75t_L g154 ( 
.A1(n_29),
.A2(n_92),
.B(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_30),
.B(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_32),
.A2(n_33),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_32),
.A2(n_33),
.B1(n_182),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_33),
.B(n_177),
.C(n_182),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_33),
.B(n_134),
.C(n_209),
.Y(n_214)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_34),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_36),
.B1(n_41),
.B2(n_42),
.Y(n_43)
);

AOI22x1_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_36),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_36),
.B(n_202),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_39),
.A2(n_44),
.B(n_45),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_39),
.B(n_44),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_40),
.A2(n_86),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_44),
.A2(n_83),
.B(n_84),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_62),
.B1(n_75),
.B2(n_76),
.Y(n_48)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_49),
.B(n_97),
.C(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_49),
.A2(n_75),
.B1(n_145),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_49),
.A2(n_75),
.B1(n_94),
.B2(n_95),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_49),
.B(n_94),
.C(n_216),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_54),
.B(n_58),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_50),
.A2(n_54),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_59),
.B(n_60),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_51),
.A2(n_244),
.B(n_246),
.Y(n_243)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_55),
.Y(n_57)
);

AO22x1_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_57),
.B1(n_70),
.B2(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_55),
.B(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_58),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_62),
.A2(n_76),
.B1(n_118),
.B2(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_62),
.B(n_118),
.C(n_129),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_69),
.B1(n_72),
.B2(n_74),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OA21x2_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_70),
.B(n_71),
.C(n_72),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_70),
.Y(n_71)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_66),
.B(n_132),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_74),
.Y(n_100)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_82),
.B2(n_87),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_82),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_87),
.B1(n_109),
.B2(n_112),
.Y(n_108)
);

INVxp33_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_80),
.B(n_93),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_87),
.A2(n_105),
.B(n_112),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_88),
.B(n_230),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.C(n_97),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_89),
.A2(n_90),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_91),
.A2(n_94),
.B1(n_95),
.B2(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_91),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_94),
.A2(n_95),
.B1(n_201),
.B2(n_203),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_94),
.B(n_203),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_97),
.A2(n_98),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_97),
.A2(n_98),
.B1(n_239),
.B2(n_248),
.Y(n_238)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_99),
.B(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_122),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_113),
.B2(n_114),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_104),
.B(n_113),
.C(n_122),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_109),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_118),
.B(n_121),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_118),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g241 ( 
.A(n_117),
.B(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_153),
.C(n_154),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_118),
.A2(n_137),
.B1(n_178),
.B2(n_181),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_121),
.A2(n_238),
.B1(n_249),
.B2(n_250),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_121),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_227),
.B(n_231),
.Y(n_123)
);

OAI211xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_156),
.B(n_170),
.C(n_226),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_146),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_146),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_138),
.B2(n_139),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_141),
.C(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_136),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_133),
.A2(n_134),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_134),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_134),
.B(n_197),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.C(n_152),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_152),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_154),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_SL g170 ( 
.A(n_157),
.B(n_171),
.C(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_158),
.B(n_159),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_160),
.B(n_162),
.C(n_168),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_167),
.B2(n_168),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_188),
.B(n_225),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_174),
.B(n_176),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_178),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_200),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_219),
.B(n_224),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_213),
.B(n_218),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_205),
.B(n_212),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_199),
.B(n_204),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_196),
.B(n_198),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_201),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_211),
.Y(n_212)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_209),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_215),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_223),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_229),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_233),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_253),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_252),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_252),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_251),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_243),
.B2(n_247),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_243),
.Y(n_247)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);


endmodule