module fake_jpeg_20541_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_2),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_68),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_2),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_70),
.Y(n_75)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_72),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_72),
.A2(n_51),
.B1(n_60),
.B2(n_48),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_77),
.B1(n_79),
.B2(n_81),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_41),
.B1(n_47),
.B2(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_50),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_64),
.B1(n_57),
.B2(n_62),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_49),
.B1(n_58),
.B2(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_89),
.Y(n_103)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_86),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_73),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_77),
.B(n_63),
.Y(n_89)
);

NOR2x1_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_44),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_94),
.B1(n_4),
.B2(n_5),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_93),
.B(n_59),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_73),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_98),
.B(n_104),
.Y(n_113)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_59),
.A3(n_55),
.B1(n_45),
.B2(n_6),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_27),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_28),
.B1(n_36),
.B2(n_35),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_106),
.B1(n_107),
.B2(n_39),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_3),
.Y(n_104)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_90),
.A2(n_7),
.B1(n_13),
.B2(n_15),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_18),
.B1(n_21),
.B2(n_25),
.Y(n_107)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_108),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_121),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_122),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_118),
.B(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_116),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_109),
.B1(n_120),
.B2(n_99),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_103),
.B(n_119),
.C(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_129),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_30),
.B(n_31),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_34),
.Y(n_132)
);


endmodule