module fake_jpeg_26062_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_3),
.B(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_32),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_0),
.C(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_35),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_20),
.Y(n_34)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_14),
.B(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_27),
.B1(n_16),
.B2(n_21),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_43),
.B1(n_34),
.B2(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_15),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_27),
.B1(n_16),
.B2(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_30),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_28),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_57),
.B1(n_60),
.B2(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_56),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

AND2x6_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_10),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_SL g71 ( 
.A(n_54),
.B(n_40),
.C(n_24),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_59),
.Y(n_80)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_34),
.B1(n_47),
.B2(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_17),
.B1(n_13),
.B2(n_22),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_62),
.Y(n_70)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_28),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_65),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_28),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_79),
.B1(n_48),
.B2(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_71),
.B(n_82),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_28),
.C(n_40),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_58),
.C(n_66),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_78),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_79),
.B1(n_60),
.B2(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_38),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_30),
.B1(n_24),
.B2(n_8),
.Y(n_79)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_22),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_80),
.B1(n_71),
.B2(n_72),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_88),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_92),
.B1(n_79),
.B2(n_82),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_70),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_63),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_95),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_53),
.B1(n_54),
.B2(n_64),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_65),
.B(n_62),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_74),
.B(n_75),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_24),
.C(n_26),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_96),
.B(n_102),
.Y(n_108)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_103),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_74),
.B(n_69),
.Y(n_101)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_22),
.B1(n_17),
.B2(n_13),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_13),
.B1(n_17),
.B2(n_26),
.Y(n_104)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_25),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_19),
.Y(n_113)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_87),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_88),
.C(n_85),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_24),
.C(n_25),
.Y(n_119)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_95),
.C(n_97),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_116),
.C(n_119),
.Y(n_121)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_96),
.A3(n_102),
.B1(n_86),
.B2(n_100),
.C1(n_106),
.C2(n_103),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_112),
.B(n_109),
.Y(n_124)
);

AOI321xp33_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_87),
.A3(n_104),
.B1(n_106),
.B2(n_14),
.C(n_23),
.Y(n_118)
);

AOI31xp67_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_23),
.A3(n_19),
.B(n_24),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_112),
.B(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_123),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_120),
.B(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_125),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_121),
.A2(n_111),
.B1(n_107),
.B2(n_109),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_107),
.C(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_9),
.Y(n_132)
);

AOI322xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_6),
.C2(n_8),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_131),
.B(n_129),
.Y(n_134)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

OAI31xp33_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_127),
.A3(n_130),
.B(n_12),
.Y(n_135)
);

AOI221xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_4),
.B1(n_6),
.B2(n_133),
.C(n_120),
.Y(n_136)
);


endmodule