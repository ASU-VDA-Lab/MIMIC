module fake_jpeg_2750_n_575 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_575);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_575;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_5),
.B(n_12),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_53),
.B(n_60),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_58),
.B(n_61),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_24),
.B(n_18),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_63),
.B(n_68),
.Y(n_159)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_64),
.Y(n_158)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_65),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_21),
.B(n_17),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_79),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_0),
.B(n_1),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_71),
.B(n_37),
.C(n_36),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_24),
.B(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_72),
.B(n_77),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_73),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_17),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_80),
.Y(n_171)
);

BUFx4f_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_40),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_93),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_30),
.B(n_16),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_84),
.B(n_94),
.Y(n_155)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_28),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_30),
.B(n_15),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_91),
.B(n_95),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_40),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_34),
.B(n_14),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_34),
.B(n_13),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_35),
.B(n_14),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_101),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_40),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_29),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_19),
.Y(n_106)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_35),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_54),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_122),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_75),
.A2(n_23),
.B1(n_32),
.B2(n_29),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_123),
.A2(n_137),
.B1(n_162),
.B2(n_20),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_55),
.A2(n_23),
.B1(n_32),
.B2(n_29),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_124),
.A2(n_127),
.B1(n_136),
.B2(n_74),
.Y(n_198)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_87),
.A2(n_32),
.B1(n_38),
.B2(n_19),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_101),
.B(n_38),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_131),
.B(n_132),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_62),
.A2(n_19),
.B1(n_27),
.B2(n_45),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_80),
.A2(n_51),
.B1(n_45),
.B2(n_22),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_56),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_149),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_64),
.B(n_51),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_164),
.Y(n_183)
);

AND2x4_ASAP7_75t_L g152 ( 
.A(n_71),
.B(n_25),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_152),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_57),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_69),
.B(n_49),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_156),
.B(n_165),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_66),
.A2(n_39),
.B1(n_37),
.B2(n_36),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_92),
.B(n_49),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_85),
.B(n_39),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_20),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_172),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_173),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_176),
.Y(n_238)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_178),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_135),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_179),
.B(n_187),
.Y(n_249)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_120),
.Y(n_180)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_180),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_181),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_182),
.Y(n_260)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_186),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_116),
.B(n_88),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_114),
.B(n_90),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_188),
.B(n_197),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_189),
.B(n_194),
.Y(n_252)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_120),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g236 ( 
.A(n_190),
.Y(n_236)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_191),
.Y(n_270)
);

BUFx8_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_193),
.Y(n_271)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_195),
.Y(n_273)
);

INVx2_ASAP7_75t_R g196 ( 
.A(n_125),
.Y(n_196)
);

NAND2xp33_ASAP7_75t_SL g245 ( 
.A(n_196),
.B(n_148),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_119),
.Y(n_197)
);

OA22x2_ASAP7_75t_L g283 ( 
.A1(n_198),
.A2(n_46),
.B1(n_31),
.B2(n_118),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_150),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_199),
.B(n_203),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_142),
.Y(n_200)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_138),
.A2(n_67),
.B1(n_78),
.B2(n_104),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_201),
.A2(n_215),
.B1(n_220),
.B2(n_148),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_152),
.A2(n_99),
.B1(n_143),
.B2(n_146),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_202),
.A2(n_213),
.B1(n_225),
.B2(n_227),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_117),
.Y(n_203)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_204),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_111),
.B(n_14),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_205),
.B(n_221),
.Y(n_272)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_130),
.Y(n_207)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

CKINVDCx12_ASAP7_75t_R g208 ( 
.A(n_134),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_208),
.Y(n_254)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_209),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_210),
.Y(n_265)
);

CKINVDCx6p67_ASAP7_75t_R g212 ( 
.A(n_134),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_212),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_152),
.A2(n_81),
.B1(n_102),
.B2(n_59),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_130),
.Y(n_214)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_159),
.A2(n_89),
.B1(n_83),
.B2(n_81),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_134),
.Y(n_216)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_216),
.Y(n_269)
);

AND2x2_ASAP7_75t_SL g217 ( 
.A(n_138),
.B(n_59),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_217),
.B(n_139),
.Y(n_281)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_142),
.Y(n_219)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_219),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_160),
.A2(n_25),
.B1(n_31),
.B2(n_13),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_109),
.B(n_13),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_139),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_222),
.B(n_223),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_155),
.B(n_11),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_113),
.B(n_1),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_224),
.B(n_230),
.Y(n_276)
);

INVx11_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_226),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_143),
.A2(n_54),
.B1(n_86),
.B2(n_46),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_151),
.Y(n_228)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_228),
.Y(n_280)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_121),
.Y(n_229)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_229),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_167),
.B(n_1),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_121),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_231),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_112),
.B(n_1),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_232),
.B(n_233),
.Y(n_284)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_170),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_237),
.B(n_241),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_158),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_183),
.B(n_146),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_244),
.B(n_251),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_L g293 ( 
.A1(n_245),
.A2(n_277),
.B(n_261),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_247),
.B(n_264),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_184),
.A2(n_127),
.B(n_136),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_248),
.A2(n_180),
.B(n_214),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_183),
.B(n_137),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_177),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_185),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_198),
.A2(n_123),
.B1(n_157),
.B2(n_108),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_258),
.A2(n_283),
.B1(n_285),
.B2(n_227),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_108),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_261),
.B(n_263),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_157),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_189),
.B(n_151),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_206),
.B(n_115),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_282),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_202),
.A2(n_124),
.B1(n_147),
.B2(n_161),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_213),
.A2(n_140),
.B1(n_129),
.B2(n_161),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_175),
.A2(n_118),
.B1(n_147),
.B2(n_161),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_287),
.Y(n_326)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_243),
.Y(n_288)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_288),
.Y(n_341)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_289),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_290),
.Y(n_340)
);

CKINVDCx12_ASAP7_75t_R g291 ( 
.A(n_254),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_291),
.Y(n_352)
);

BUFx12_ASAP7_75t_L g292 ( 
.A(n_236),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_292),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g370 ( 
.A(n_293),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g377 ( 
.A(n_295),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_267),
.B(n_175),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_297),
.B(n_302),
.Y(n_345)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_298),
.Y(n_375)
);

AND2x6_ASAP7_75t_L g299 ( 
.A(n_252),
.B(n_212),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_299),
.B(n_327),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_196),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_300),
.A2(n_325),
.B(n_329),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_248),
.A2(n_218),
.B(n_212),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_301),
.A2(n_283),
.B(n_259),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_249),
.B(n_174),
.Y(n_302)
);

O2A1O1Ixp33_ASAP7_75t_L g303 ( 
.A1(n_251),
.A2(n_192),
.B(n_181),
.C(n_190),
.Y(n_303)
);

O2A1O1Ixp33_ASAP7_75t_L g372 ( 
.A1(n_303),
.A2(n_317),
.B(n_273),
.C(n_260),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_262),
.B(n_200),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_304),
.B(n_313),
.Y(n_351)
);

INVx13_ASAP7_75t_L g305 ( 
.A(n_254),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_305),
.Y(n_348)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_250),
.Y(n_307)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_307),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_252),
.A2(n_210),
.B1(n_226),
.B2(n_140),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_308),
.A2(n_335),
.B1(n_285),
.B2(n_255),
.Y(n_357)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_270),
.Y(n_309)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_309),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_243),
.Y(n_310)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_310),
.Y(n_359)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_270),
.Y(n_311)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_311),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_272),
.B(n_219),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_238),
.Y(n_314)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_314),
.Y(n_367)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_286),
.Y(n_315)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_315),
.Y(n_378)
);

INVx13_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_316),
.Y(n_344)
);

O2A1O1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_244),
.A2(n_192),
.B(n_225),
.C(n_228),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_238),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_318),
.B(n_319),
.Y(n_354)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_235),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_240),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_320),
.B(n_321),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_277),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_246),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_322),
.Y(n_337)
);

INVx13_ASAP7_75t_L g323 ( 
.A(n_253),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_323),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_245),
.B(n_216),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_324),
.A2(n_275),
.B(n_256),
.Y(n_362)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_266),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_268),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_328),
.B(n_330),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_258),
.A2(n_178),
.B1(n_207),
.B2(n_195),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_241),
.B(n_274),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_253),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_332),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_284),
.B(n_182),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_242),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_334),
.B(n_336),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_252),
.A2(n_129),
.B1(n_193),
.B2(n_204),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_234),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_294),
.B(n_281),
.C(n_264),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_343),
.B(n_355),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_301),
.A2(n_239),
.B(n_282),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_353),
.A2(n_363),
.B(n_373),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_294),
.B(n_237),
.C(n_269),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_312),
.B(n_276),
.Y(n_356)
);

XNOR2x1_ASAP7_75t_L g381 ( 
.A(n_356),
.B(n_374),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_357),
.B(n_366),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_362),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_294),
.A2(n_247),
.B1(n_283),
.B2(n_278),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_364),
.A2(n_369),
.B1(n_324),
.B2(n_326),
.Y(n_402)
);

OA21x2_ASAP7_75t_L g366 ( 
.A1(n_296),
.A2(n_283),
.B(n_256),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_321),
.A2(n_265),
.B1(n_186),
.B2(n_271),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_368),
.A2(n_346),
.B1(n_378),
.B2(n_347),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_296),
.A2(n_279),
.B1(n_271),
.B2(n_273),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_372),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_296),
.A2(n_259),
.B(n_260),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_312),
.B(n_279),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_300),
.A2(n_172),
.B1(n_176),
.B2(n_173),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_326),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_306),
.B(n_182),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_379),
.B(n_289),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_337),
.B(n_331),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_380),
.B(n_389),
.Y(n_434)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_346),
.Y(n_382)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_382),
.Y(n_422)
);

INVx13_ASAP7_75t_L g383 ( 
.A(n_352),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_383),
.Y(n_446)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_384),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_366),
.A2(n_325),
.B1(n_308),
.B2(n_299),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_385),
.A2(n_388),
.B1(n_414),
.B2(n_370),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_358),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_386),
.B(n_392),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_365),
.Y(n_387)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_387),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_366),
.A2(n_333),
.B1(n_335),
.B2(n_306),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_377),
.B(n_319),
.Y(n_389)
);

INVx13_ASAP7_75t_L g391 ( 
.A(n_348),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g420 ( 
.A(n_391),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_354),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_356),
.B(n_336),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_393),
.B(n_395),
.Y(n_425)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_394),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_365),
.B(n_333),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_378),
.Y(n_396)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_396),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_342),
.B(n_300),
.Y(n_397)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_397),
.Y(n_447)
);

INVx13_ASAP7_75t_L g400 ( 
.A(n_344),
.Y(n_400)
);

OAI21xp33_ASAP7_75t_SL g448 ( 
.A1(n_400),
.A2(n_401),
.B(n_407),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_342),
.B(n_374),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_402),
.A2(n_340),
.B1(n_357),
.B2(n_369),
.Y(n_432)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_350),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_405),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_345),
.B(n_327),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_404),
.B(n_408),
.Y(n_417)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_349),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_362),
.B(n_303),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_406),
.A2(n_411),
.B(n_415),
.Y(n_423)
);

AND2x2_ASAP7_75t_SL g407 ( 
.A(n_343),
.B(n_317),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_351),
.B(n_355),
.Y(n_408)
);

AOI21x1_ASAP7_75t_SL g430 ( 
.A1(n_409),
.A2(n_353),
.B(n_339),
.Y(n_430)
);

INVx13_ASAP7_75t_L g410 ( 
.A(n_344),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_413),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_338),
.B(n_364),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_412),
.B(n_379),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_375),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_363),
.A2(n_315),
.B1(n_318),
.B2(n_314),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_386),
.B(n_338),
.Y(n_419)
);

NAND3xp33_ASAP7_75t_L g454 ( 
.A(n_419),
.B(n_427),
.C(n_431),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_421),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_423),
.B(n_372),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_426),
.A2(n_406),
.B1(n_414),
.B2(n_409),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_387),
.B(n_307),
.Y(n_427)
);

A2O1A1Ixp33_ASAP7_75t_SL g464 ( 
.A1(n_430),
.A2(n_399),
.B(n_406),
.C(n_390),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_392),
.B(n_361),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_432),
.A2(n_433),
.B1(n_385),
.B2(n_398),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_399),
.A2(n_340),
.B1(n_368),
.B2(n_339),
.Y(n_433)
);

XNOR2x1_ASAP7_75t_L g435 ( 
.A(n_381),
.B(n_376),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_SL g461 ( 
.A(n_435),
.B(n_402),
.C(n_399),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_405),
.B(n_361),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_437),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_416),
.B(n_373),
.C(n_350),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_438),
.B(n_441),
.C(n_449),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_395),
.B(n_309),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g467 ( 
.A(n_439),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_371),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_440),
.B(n_443),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_381),
.B(n_360),
.C(n_371),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_407),
.B(n_401),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_411),
.B(n_397),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_445),
.B(n_450),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_407),
.B(n_360),
.C(n_367),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_411),
.B(n_311),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_428),
.Y(n_453)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_453),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_413),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_455),
.B(n_457),
.Y(n_492)
);

FAx1_ASAP7_75t_SL g457 ( 
.A(n_448),
.B(n_390),
.CI(n_398),
.CON(n_457),
.SN(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_428),
.B(n_384),
.Y(n_458)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_458),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_459),
.A2(n_477),
.B1(n_423),
.B2(n_447),
.Y(n_485)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_418),
.Y(n_460)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_460),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_461),
.B(n_410),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_425),
.B(n_367),
.Y(n_462)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_462),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_425),
.B(n_396),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_463),
.B(n_475),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_464),
.A2(n_469),
.B(n_433),
.Y(n_487)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_436),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_465),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_438),
.B(n_388),
.C(n_403),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_466),
.B(n_476),
.C(n_478),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_420),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_468),
.A2(n_472),
.B1(n_473),
.B2(n_410),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_415),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_443),
.B(n_409),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_471),
.B(n_426),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_446),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_440),
.B(n_394),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_441),
.B(n_382),
.C(n_375),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_422),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_449),
.B(n_328),
.C(n_298),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_479),
.A2(n_432),
.B1(n_429),
.B2(n_446),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_456),
.B(n_421),
.C(n_435),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_481),
.B(n_483),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_456),
.B(n_429),
.C(n_447),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_484),
.B(n_496),
.Y(n_517)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_485),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_430),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_486),
.B(n_495),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_487),
.A2(n_479),
.B(n_469),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_488),
.B(n_464),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_417),
.C(n_442),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_490),
.B(n_491),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_476),
.B(n_444),
.C(n_442),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_466),
.B(n_444),
.C(n_422),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_494),
.B(n_499),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_474),
.B(n_341),
.Y(n_495)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_498),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_341),
.C(n_359),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_454),
.A2(n_359),
.B1(n_400),
.B2(n_334),
.Y(n_501)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_501),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_467),
.A2(n_400),
.B1(n_383),
.B2(n_288),
.Y(n_503)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_503),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_500),
.B(n_452),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_507),
.B(n_513),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_480),
.B(n_471),
.C(n_461),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_509),
.B(n_512),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_480),
.B(n_458),
.C(n_451),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_453),
.C(n_473),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_514),
.A2(n_517),
.B(n_504),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_483),
.B(n_457),
.C(n_464),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_515),
.B(n_518),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_491),
.B(n_457),
.C(n_464),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_502),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_520),
.A2(n_482),
.B1(n_489),
.B2(n_493),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_490),
.B(n_383),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_521),
.B(n_316),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_522),
.A2(n_292),
.B(n_242),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_499),
.C(n_495),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_523),
.B(n_529),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_511),
.Y(n_524)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_524),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_525),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_484),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_526),
.B(n_528),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_515),
.A2(n_492),
.B(n_481),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_527),
.A2(n_231),
.B(n_229),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_508),
.B(n_486),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_516),
.A2(n_482),
.B1(n_497),
.B2(n_496),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_512),
.B(n_310),
.C(n_391),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_533),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_510),
.A2(n_514),
.B1(n_519),
.B2(n_522),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_534),
.B(n_535),
.Y(n_548)
);

BUFx24_ASAP7_75t_SL g535 ( 
.A(n_505),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_513),
.A2(n_391),
.B1(n_305),
.B2(n_323),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_536),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_537),
.A2(n_539),
.B(n_509),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_538),
.B(n_233),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_530),
.A2(n_517),
.B(n_518),
.Y(n_540)
);

AOI21xp33_ASAP7_75t_SL g554 ( 
.A1(n_540),
.A2(n_532),
.B(n_531),
.Y(n_554)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_541),
.Y(n_559)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_542),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_523),
.B(n_292),
.C(n_233),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_547),
.B(n_528),
.Y(n_555)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_551),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_533),
.B(n_2),
.Y(n_552)
);

NOR2x1_ASAP7_75t_L g557 ( 
.A(n_552),
.B(n_524),
.Y(n_557)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_554),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_555),
.B(n_556),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_544),
.B(n_526),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_557),
.B(n_25),
.C(n_46),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_543),
.A2(n_539),
.B1(n_25),
.B2(n_31),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_558),
.B(n_545),
.C(n_541),
.Y(n_561)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_561),
.Y(n_568)
);

AOI322xp5_ASAP7_75t_L g563 ( 
.A1(n_559),
.A2(n_548),
.A3(n_546),
.B1(n_549),
.B2(n_544),
.C1(n_550),
.C2(n_547),
.Y(n_563)
);

O2A1O1Ixp33_ASAP7_75t_SL g567 ( 
.A1(n_563),
.A2(n_553),
.B(n_25),
.C(n_4),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_564),
.B(n_560),
.C(n_555),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_566),
.B(n_565),
.Y(n_569)
);

AOI322xp5_ASAP7_75t_L g570 ( 
.A1(n_567),
.A2(n_568),
.A3(n_562),
.B1(n_5),
.B2(n_7),
.C1(n_2),
.C2(n_9),
.Y(n_570)
);

NAND2x1p5_ASAP7_75t_SL g571 ( 
.A(n_569),
.B(n_570),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g572 ( 
.A1(n_571),
.A2(n_3),
.B(n_7),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_572),
.B(n_8),
.C(n_9),
.Y(n_573)
);

NOR2xp67_ASAP7_75t_L g574 ( 
.A(n_573),
.B(n_8),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_SL g575 ( 
.A1(n_574),
.A2(n_8),
.B(n_9),
.Y(n_575)
);


endmodule