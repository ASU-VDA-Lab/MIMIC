module real_jpeg_10435_n_12 (n_5, n_4, n_8, n_0, n_278, n_1, n_11, n_2, n_6, n_277, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_278;
input n_1;
input n_11;
input n_2;
input n_6;
input n_277;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_262;
wire n_19;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_130;
wire n_144;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_167;
wire n_244;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_1),
.A2(n_86),
.B1(n_87),
.B2(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_1),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_1),
.A2(n_8),
.B(n_86),
.Y(n_143)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_4),
.A2(n_40),
.B(n_44),
.C(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_40),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_4),
.A2(n_8),
.B(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_SL g73 ( 
.A(n_5),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_7),
.A2(n_29),
.B1(n_40),
.B2(n_42),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_7),
.A2(n_29),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_7),
.A2(n_29),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_8),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_8),
.B(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_8),
.A2(n_35),
.B1(n_86),
.B2(n_87),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_8),
.A2(n_73),
.B(n_87),
.C(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_8),
.B(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_8),
.A2(n_35),
.B1(n_133),
.B2(n_134),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_156),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_9),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_9),
.A2(n_40),
.B1(n_42),
.B2(n_156),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_9),
.A2(n_86),
.B1(n_87),
.B2(n_156),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_9),
.A2(n_133),
.B1(n_134),
.B2(n_156),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_10),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_11),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_11),
.A2(n_40),
.B1(n_42),
.B2(n_174),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_11),
.A2(n_86),
.B1(n_87),
.B2(n_174),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_263),
.Y(n_12)
);

OAI321xp33_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_231),
.A3(n_256),
.B1(n_261),
.B2(n_262),
.C(n_277),
.Y(n_13)
);

AOI321xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_185),
.A3(n_205),
.B1(n_225),
.B2(n_230),
.C(n_278),
.Y(n_14)
);

NOR3xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_148),
.C(n_182),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_120),
.B(n_147),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_101),
.B(n_119),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_79),
.B(n_100),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_64),
.B(n_78),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_54),
.B(n_63),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.Y(n_21)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_22),
.B(n_36),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_22),
.A2(n_56),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_22),
.B(n_105),
.C(n_111),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_30),
.B(n_31),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_24),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_25),
.B(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_30),
.B(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_30),
.A2(n_98),
.B1(n_155),
.B2(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_31),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_32),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_35),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_33),
.A2(n_154),
.B(n_157),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_34),
.B(n_97),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_42),
.B(n_45),
.C(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_44),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_SL g95 ( 
.A1(n_35),
.A2(n_40),
.B(n_74),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_35),
.A2(n_114),
.B(n_133),
.C(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_37),
.B(n_51),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_37),
.A2(n_53),
.B1(n_84),
.B2(n_92),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_37),
.B(n_84),
.C(n_99),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_37),
.A2(n_53),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B(n_46),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_39),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_76)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_40),
.A2(n_42),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_44),
.B(n_48),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_44),
.A2(n_201),
.B(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_44),
.A2(n_48),
.B1(n_201),
.B2(n_212),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_46),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_47),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_53),
.B(n_153),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B(n_62),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_60),
.B(n_61),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_61),
.A2(n_67),
.B1(n_68),
.B2(n_77),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_69),
.C(n_76),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_61),
.A2(n_77),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_61),
.B(n_141),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_66),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_85),
.B(n_88),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_71),
.A2(n_85),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_71),
.B(n_106),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_71),
.A2(n_106),
.B1(n_238),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_73),
.B(n_87),
.C(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_72),
.A2(n_237),
.B(n_239),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_73),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_87),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_75),
.A2(n_76),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_75),
.A2(n_76),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_75),
.B(n_171),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_104),
.C(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_80),
.B(n_81),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_93),
.B2(n_99),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_84),
.A2(n_92),
.B1(n_126),
.B2(n_129),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_84),
.B(n_126),
.C(n_131),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_84),
.A2(n_92),
.B1(n_161),
.B2(n_162),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_84),
.B(n_161),
.C(n_195),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_86),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_88),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_89),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_93),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_97),
.B(n_173),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_103),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_116),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_108),
.B1(n_109),
.B2(n_115),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_105),
.A2(n_115),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_105),
.B(n_161),
.C(n_164),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_132),
.B(n_135),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_114),
.B(n_133),
.C(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_113),
.A2(n_136),
.B1(n_137),
.B2(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_113),
.B(n_137),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_113),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_133),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_115),
.A2(n_211),
.B(n_213),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_115),
.B(n_211),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_117),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_122),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_139),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_123),
.B(n_140),
.C(n_146),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_130),
.B2(n_131),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_126),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_128),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_130),
.A2(n_131),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_130),
.A2(n_131),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_130),
.A2(n_131),
.B1(n_248),
.B2(n_254),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_130),
.B(n_240),
.C(n_243),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_130),
.B(n_254),
.C(n_255),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_131),
.B(n_176),
.C(n_178),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_132),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_133),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_135),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_136),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_140),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_144),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g226 ( 
.A1(n_149),
.A2(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_165),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_150),
.B(n_165),
.Y(n_228)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_158),
.CI(n_159),
.CON(n_150),
.SN(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_161),
.A2(n_162),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_161),
.B(n_241),
.C(n_252),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_181),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_175),
.C(n_181),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_180),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_184),
.Y(n_227)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_186),
.A2(n_226),
.B(n_229),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_187),
.B(n_188),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_204),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_196),
.B2(n_197),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_197),
.C(n_204),
.Y(n_206)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_192),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_203),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_199),
.B1(n_217),
.B2(n_220),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_200),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_199),
.A2(n_215),
.B(n_217),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_200),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_207),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_223),
.B2(n_224),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_214),
.B1(n_221),
.B2(n_222),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_210),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_222),
.C(n_224),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_212),
.B(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_233),
.C(n_244),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_213),
.B(n_233),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_214),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_217),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_223),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_246),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_246),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_240),
.B1(n_241),
.B2(n_243),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_236),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_240),
.A2(n_241),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_244),
.A2(n_245),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_255),
.Y(n_246)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_257),
.B(n_258),
.Y(n_261)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_259),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_274),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_273),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_273),
.Y(n_274)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_266),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_269),
.CI(n_272),
.CON(n_266),
.SN(n_266)
);


endmodule