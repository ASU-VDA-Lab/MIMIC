module real_aes_16717_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_891;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
AND2x4_ASAP7_75t_L g884 ( .A(n_0), .B(n_885), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_1), .A2(n_32), .B1(n_135), .B2(n_185), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_2), .A2(n_93), .B1(n_519), .B2(n_520), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_2), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_3), .A2(n_10), .B1(n_545), .B2(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g885 ( .A(n_4), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_5), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_6), .A2(n_11), .B1(n_565), .B2(n_566), .Y(n_564) );
OR2x2_ASAP7_75t_L g114 ( .A(n_7), .B(n_28), .Y(n_114) );
BUFx2_ASAP7_75t_L g888 ( .A(n_7), .Y(n_888) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_8), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_9), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_12), .B(n_150), .Y(n_149) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_13), .A2(n_99), .B1(n_229), .B2(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_14), .A2(n_29), .B1(n_576), .B2(n_577), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_15), .B(n_150), .Y(n_592) );
OAI21x1_ASAP7_75t_L g130 ( .A1(n_16), .A2(n_45), .B(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_17), .B(n_244), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_18), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_19), .A2(n_37), .B1(n_205), .B2(n_234), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_20), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_21), .A2(n_42), .B1(n_205), .B2(n_545), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_22), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_23), .B(n_576), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_24), .B(n_179), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_25), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_26), .B(n_128), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_27), .Y(n_228) );
HB1xp67_ASAP7_75t_L g890 ( .A(n_28), .Y(n_890) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_30), .A2(n_82), .B1(n_135), .B2(n_620), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_31), .A2(n_36), .B1(n_135), .B2(n_568), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g864 ( .A(n_33), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_34), .A2(n_49), .B1(n_545), .B2(n_547), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_35), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_38), .B(n_150), .Y(n_218) );
INVx2_ASAP7_75t_L g107 ( .A(n_39), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_40), .B(n_222), .Y(n_239) );
INVx1_ASAP7_75t_L g112 ( .A(n_41), .Y(n_112) );
BUFx3_ASAP7_75t_L g515 ( .A(n_41), .Y(n_515) );
OAI22x1_ASAP7_75t_SL g503 ( .A1(n_43), .A2(n_504), .B1(n_505), .B2(n_508), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_43), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_44), .B(n_168), .Y(n_246) );
AND2x2_ASAP7_75t_L g207 ( .A(n_46), .B(n_168), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_47), .B(n_165), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_48), .A2(n_78), .B1(n_506), .B2(n_507), .Y(n_505) );
INVxp67_ASAP7_75t_L g506 ( .A(n_48), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_50), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_51), .B(n_234), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_52), .A2(n_69), .B1(n_234), .B2(n_547), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_53), .A2(n_72), .B1(n_135), .B2(n_568), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_54), .B(n_184), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_55), .A2(n_139), .B(n_148), .C(n_198), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_56), .A2(n_95), .B1(n_545), .B2(n_566), .Y(n_601) );
INVx1_ASAP7_75t_L g131 ( .A(n_57), .Y(n_131) );
AND2x4_ASAP7_75t_L g153 ( .A(n_58), .B(n_154), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_59), .A2(n_60), .B1(n_205), .B2(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_61), .B(n_128), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_62), .B(n_168), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_63), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_64), .B(n_205), .Y(n_221) );
CKINVDCx16_ASAP7_75t_R g873 ( .A(n_65), .Y(n_873) );
INVx1_ASAP7_75t_L g154 ( .A(n_66), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_67), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_68), .B(n_128), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_70), .B(n_135), .Y(n_177) );
NAND3xp33_ASAP7_75t_L g240 ( .A(n_71), .B(n_185), .C(n_222), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_73), .B(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g141 ( .A(n_74), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_75), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_76), .B(n_150), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_77), .B(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g507 ( .A(n_78), .Y(n_507) );
XNOR2x1_ASAP7_75t_L g528 ( .A(n_78), .B(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_79), .A2(n_96), .B1(n_148), .B2(n_205), .Y(n_621) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_80), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g641 ( .A(n_81), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_83), .A2(n_89), .B1(n_179), .B2(n_267), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_84), .A2(n_103), .B1(n_877), .B2(n_891), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_85), .B(n_150), .Y(n_230) );
NAND2xp33_ASAP7_75t_SL g166 ( .A(n_86), .B(n_138), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_87), .B(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_88), .B(n_128), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_90), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_91), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g527 ( .A(n_91), .Y(n_527) );
NAND2xp33_ASAP7_75t_L g595 ( .A(n_92), .B(n_150), .Y(n_595) );
INVx1_ASAP7_75t_L g520 ( .A(n_93), .Y(n_520) );
NAND2xp33_ASAP7_75t_L g137 ( .A(n_94), .B(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_97), .B(n_168), .Y(n_188) );
NAND3xp33_ASAP7_75t_L g162 ( .A(n_98), .B(n_138), .C(n_161), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_100), .B(n_135), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_101), .B(n_179), .Y(n_182) );
AO21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_115), .B(n_509), .Y(n_103) );
NOR2xp33_ASAP7_75t_SL g104 ( .A(n_105), .B(n_108), .Y(n_104) );
BUFx8_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g512 ( .A(n_107), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_107), .B(n_869), .Y(n_868) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
CKINVDCx8_ASAP7_75t_R g876 ( .A(n_109), .Y(n_876) );
AND2x6_ASAP7_75t_SL g109 ( .A(n_110), .B(n_113), .Y(n_109) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
HB1xp67_ASAP7_75t_L g881 ( .A(n_112), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_113), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NOR2x1_ASAP7_75t_L g871 ( .A(n_114), .B(n_515), .Y(n_871) );
INVxp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
XNOR2x1_ASAP7_75t_L g116 ( .A(n_117), .B(n_503), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g529 ( .A(n_118), .Y(n_529) );
NAND4xp75_ASAP7_75t_L g118 ( .A(n_119), .B(n_349), .C(n_422), .D(n_481), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_305), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_275), .Y(n_120) );
OAI221xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_208), .B1(n_247), .B2(n_252), .C(n_256), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI21xp33_ASAP7_75t_SL g256 ( .A1(n_123), .A2(n_257), .B(n_261), .Y(n_256) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_171), .Y(n_123) );
AND2x2_ASAP7_75t_L g302 ( .A(n_124), .B(n_259), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_124), .B(n_313), .Y(n_375) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_155), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx2_ASAP7_75t_L g258 ( .A(n_126), .Y(n_258) );
INVx4_ASAP7_75t_L g281 ( .A(n_126), .Y(n_281) );
AND2x2_ASAP7_75t_L g309 ( .A(n_126), .B(n_172), .Y(n_309) );
OR2x2_ASAP7_75t_L g471 ( .A(n_126), .B(n_255), .Y(n_471) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_132), .Y(n_126) );
INVx2_ASAP7_75t_L g639 ( .A(n_128), .Y(n_639) );
INVx4_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x4_ASAP7_75t_SL g151 ( .A(n_129), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_SL g157 ( .A(n_129), .Y(n_157) );
INVx2_ASAP7_75t_L g213 ( .A(n_129), .Y(n_213) );
BUFx3_ASAP7_75t_L g580 ( .A(n_129), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_129), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_SL g588 ( .A(n_129), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_129), .B(n_604), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_129), .B(n_641), .Y(n_640) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g170 ( .A(n_130), .Y(n_170) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_142), .B(n_151), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_137), .B(n_139), .Y(n_133) );
OAI22xp33_ASAP7_75t_L g203 ( .A1(n_135), .A2(n_204), .B1(n_205), .B2(n_206), .Y(n_203) );
INVx1_ASAP7_75t_L g547 ( .A(n_135), .Y(n_547) );
INVx1_ASAP7_75t_L g566 ( .A(n_135), .Y(n_566) );
INVx4_ASAP7_75t_L g568 ( .A(n_135), .Y(n_568) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_136), .Y(n_138) );
INVx1_ASAP7_75t_L g148 ( .A(n_136), .Y(n_148) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_136), .Y(n_150) );
INVx1_ASAP7_75t_L g165 ( .A(n_136), .Y(n_165) );
INVx1_ASAP7_75t_L g180 ( .A(n_136), .Y(n_180) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_136), .Y(n_185) );
INVx2_ASAP7_75t_L g200 ( .A(n_136), .Y(n_200) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_136), .Y(n_205) );
INVx1_ASAP7_75t_L g217 ( .A(n_136), .Y(n_217) );
INVx1_ASAP7_75t_L g270 ( .A(n_136), .Y(n_270) );
INVx2_ASAP7_75t_L g234 ( .A(n_138), .Y(n_234) );
INVx1_ASAP7_75t_L g576 ( .A(n_138), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_139), .A2(n_164), .B(n_166), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_139), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_139), .A2(n_216), .B(n_218), .Y(n_215) );
BUFx4f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g146 ( .A(n_141), .Y(n_146) );
INVx1_ASAP7_75t_L g161 ( .A(n_141), .Y(n_161) );
BUFx8_ASAP7_75t_L g222 ( .A(n_141), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_145), .B1(n_147), .B2(n_149), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_144), .A2(n_232), .B(n_233), .Y(n_231) );
INVx2_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx3_ASAP7_75t_L g187 ( .A(n_146), .Y(n_187) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_150), .A2(n_160), .B(n_162), .Y(n_159) );
INVx1_ASAP7_75t_L g244 ( .A(n_150), .Y(n_244) );
INVx3_ASAP7_75t_L g545 ( .A(n_150), .Y(n_545) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_152), .A2(n_159), .B(n_163), .Y(n_158) );
OAI21x1_ASAP7_75t_L g175 ( .A1(n_152), .A2(n_176), .B(n_181), .Y(n_175) );
OAI21x1_ASAP7_75t_L g214 ( .A1(n_152), .A2(n_215), .B(n_219), .Y(n_214) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_152), .A2(n_227), .B(n_231), .Y(n_226) );
OAI21x1_ASAP7_75t_L g237 ( .A1(n_152), .A2(n_238), .B(n_241), .Y(n_237) );
BUFx10_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx10_ASAP7_75t_L g195 ( .A(n_153), .Y(n_195) );
INVx1_ASAP7_75t_L g557 ( .A(n_153), .Y(n_557) );
INVx2_ASAP7_75t_L g284 ( .A(n_155), .Y(n_284) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_155), .Y(n_310) );
INVx1_ASAP7_75t_L g320 ( .A(n_155), .Y(n_320) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g255 ( .A(n_156), .Y(n_255) );
AND2x2_ASAP7_75t_L g411 ( .A(n_156), .B(n_190), .Y(n_411) );
OAI21x1_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_167), .Y(n_156) );
INVx1_ASAP7_75t_L g245 ( .A(n_161), .Y(n_245) );
INVx1_ASAP7_75t_SL g569 ( .A(n_161), .Y(n_569) );
INVx1_ASAP7_75t_L g622 ( .A(n_161), .Y(n_622) );
INVx1_ASAP7_75t_L g577 ( .A(n_165), .Y(n_577) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g174 ( .A(n_169), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_169), .B(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_169), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g193 ( .A(n_170), .Y(n_193) );
INVx2_ASAP7_75t_L g273 ( .A(n_170), .Y(n_273) );
INVx2_ASAP7_75t_L g368 ( .A(n_171), .Y(n_368) );
AND2x2_ASAP7_75t_L g372 ( .A(n_171), .B(n_284), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_171), .B(n_403), .Y(n_501) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_189), .Y(n_171) );
INVx2_ASAP7_75t_L g335 ( .A(n_172), .Y(n_335) );
AND2x2_ASAP7_75t_L g429 ( .A(n_172), .B(n_295), .Y(n_429) );
AND2x2_ASAP7_75t_L g480 ( .A(n_172), .B(n_281), .Y(n_480) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g254 ( .A(n_173), .Y(n_254) );
OAI21x1_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_188), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_174), .A2(n_226), .B(n_235), .Y(n_225) );
OAI21x1_ASAP7_75t_L g251 ( .A1(n_174), .A2(n_226), .B(n_235), .Y(n_251) );
OAI21xp33_ASAP7_75t_SL g260 ( .A1(n_174), .A2(n_175), .B(n_188), .Y(n_260) );
INVx1_ASAP7_75t_L g565 ( .A(n_179), .Y(n_565) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_186), .Y(n_181) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g202 ( .A(n_187), .Y(n_202) );
AND2x2_ASAP7_75t_L g259 ( .A(n_189), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g283 ( .A(n_190), .Y(n_283) );
AOI21x1_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_196), .B(n_207), .Y(n_190) );
NOR2xp67_ASAP7_75t_SL g191 ( .A(n_192), .B(n_194), .Y(n_191) );
INVx2_ASAP7_75t_L g548 ( .A(n_192), .Y(n_548) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AO31x2_ASAP7_75t_L g264 ( .A1(n_193), .A2(n_195), .A3(n_265), .B(n_271), .Y(n_264) );
NOR2xp33_ASAP7_75t_SL g571 ( .A(n_193), .B(n_572), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_193), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g542 ( .A(n_194), .Y(n_542) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AO31x2_ASAP7_75t_L g562 ( .A1(n_195), .A2(n_563), .A3(n_570), .B(n_571), .Y(n_562) );
AO31x2_ASAP7_75t_L g573 ( .A1(n_195), .A2(n_574), .A3(n_580), .B(n_581), .Y(n_573) );
AO31x2_ASAP7_75t_L g635 ( .A1(n_195), .A2(n_636), .A3(n_639), .B(n_640), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_201), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
INVx2_ASAP7_75t_SL g620 ( .A(n_200), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_202), .A2(n_266), .B1(n_268), .B2(n_269), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_202), .A2(n_268), .B1(n_544), .B2(n_546), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_202), .A2(n_268), .B1(n_554), .B2(n_555), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_202), .A2(n_268), .B1(n_575), .B2(n_578), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_202), .A2(n_268), .B1(n_637), .B2(n_638), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_205), .A2(n_239), .B(n_240), .Y(n_238) );
INVx2_ASAP7_75t_L g267 ( .A(n_205), .Y(n_267) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_224), .Y(n_209) );
INVx2_ASAP7_75t_L g248 ( .A(n_210), .Y(n_248) );
AND2x2_ASAP7_75t_L g412 ( .A(n_210), .B(n_262), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_210), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_210), .B(n_433), .Y(n_442) );
OR2x2_ASAP7_75t_L g465 ( .A(n_210), .B(n_324), .Y(n_465) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NOR2xp67_ASAP7_75t_L g348 ( .A(n_211), .B(n_291), .Y(n_348) );
AND2x2_ASAP7_75t_L g454 ( .A(n_211), .B(n_263), .Y(n_454) );
BUFx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g288 ( .A(n_212), .Y(n_288) );
OAI21x1_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_223), .Y(n_212) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_213), .A2(n_237), .B(n_246), .Y(n_236) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_213), .A2(n_237), .B(n_246), .Y(n_263) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_213), .A2(n_214), .B(n_223), .Y(n_300) );
INVx2_ASAP7_75t_L g229 ( .A(n_217), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_222), .Y(n_219) );
O2A1O1Ixp5_ASAP7_75t_L g227 ( .A1(n_222), .A2(n_228), .B(n_229), .C(n_230), .Y(n_227) );
INVx6_ASAP7_75t_L g268 ( .A(n_222), .Y(n_268) );
O2A1O1Ixp5_ASAP7_75t_L g590 ( .A1(n_222), .A2(n_568), .B(n_591), .C(n_592), .Y(n_590) );
AND2x2_ASAP7_75t_L g341 ( .A(n_224), .B(n_286), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_224), .B(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_224), .B(n_397), .Y(n_405) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_236), .Y(n_224) );
AND2x2_ASAP7_75t_L g317 ( .A(n_225), .B(n_263), .Y(n_317) );
INVx1_ASAP7_75t_L g461 ( .A(n_225), .Y(n_461) );
AND2x2_ASAP7_75t_L g249 ( .A(n_236), .B(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g324 ( .A(n_236), .B(n_264), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_236), .B(n_264), .Y(n_382) );
AOI21x1_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_245), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_248), .B(n_365), .Y(n_364) );
AND2x4_ASAP7_75t_L g487 ( .A(n_248), .B(n_290), .Y(n_487) );
AND2x2_ASAP7_75t_L g417 ( .A(n_249), .B(n_418), .Y(n_417) );
INVxp67_ASAP7_75t_SL g274 ( .A(n_250), .Y(n_274) );
AND2x2_ASAP7_75t_L g298 ( .A(n_250), .B(n_299), .Y(n_298) );
BUFx3_ASAP7_75t_L g304 ( .A(n_250), .Y(n_304) );
INVxp67_ASAP7_75t_SL g340 ( .A(n_250), .Y(n_340) );
INVx1_ASAP7_75t_L g365 ( .A(n_250), .Y(n_365) );
AND2x2_ASAP7_75t_L g371 ( .A(n_250), .B(n_263), .Y(n_371) );
INVx1_ASAP7_75t_L g452 ( .A(n_250), .Y(n_452) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g294 ( .A(n_253), .B(n_295), .Y(n_294) );
AOI32xp33_ASAP7_75t_SL g426 ( .A1(n_253), .A2(n_318), .A3(n_427), .B1(n_429), .B2(n_430), .Y(n_426) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g279 ( .A(n_254), .Y(n_279) );
OR2x2_ASAP7_75t_L g328 ( .A(n_254), .B(n_284), .Y(n_328) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_255), .Y(n_332) );
INVxp67_ASAP7_75t_L g358 ( .A(n_255), .Y(n_358) );
OR2x2_ASAP7_75t_L g460 ( .A(n_255), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
OR3x2_ASAP7_75t_L g325 ( .A(n_258), .B(n_326), .C(n_328), .Y(n_325) );
INVx1_ASAP7_75t_L g431 ( .A(n_258), .Y(n_431) );
AND2x2_ASAP7_75t_L g359 ( .A(n_259), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g415 ( .A(n_259), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_259), .B(n_310), .Y(n_421) );
BUFx2_ASAP7_75t_L g314 ( .A(n_260), .Y(n_314) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_274), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_262), .B(n_298), .Y(n_297) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_262), .Y(n_494) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g291 ( .A(n_263), .Y(n_291) );
INVx1_ASAP7_75t_L g433 ( .A(n_263), .Y(n_433) );
INVx1_ASAP7_75t_L g292 ( .A(n_264), .Y(n_292) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_264), .Y(n_338) );
OR2x2_ASAP7_75t_L g379 ( .A(n_264), .B(n_300), .Y(n_379) );
AND2x2_ASAP7_75t_L g397 ( .A(n_264), .B(n_300), .Y(n_397) );
AND2x2_ASAP7_75t_L g418 ( .A(n_264), .B(n_288), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_268), .A2(n_564), .B1(n_567), .B2(n_569), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_268), .A2(n_594), .B(n_595), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_268), .A2(n_569), .B1(n_601), .B2(n_602), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_268), .A2(n_619), .B1(n_621), .B2(n_622), .Y(n_618) );
INVx1_ASAP7_75t_L g579 ( .A(n_270), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
BUFx2_ASAP7_75t_L g570 ( .A(n_273), .Y(n_570) );
BUFx2_ASAP7_75t_L g486 ( .A(n_274), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_293), .C(n_301), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_285), .Y(n_276) );
INVx3_ASAP7_75t_L g408 ( .A(n_277), .Y(n_408) );
AND2x4_ASAP7_75t_L g277 ( .A(n_278), .B(n_282), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g438 ( .A(n_279), .B(n_394), .Y(n_438) );
INVx1_ASAP7_75t_L g360 ( .A(n_280), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_280), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g445 ( .A(n_280), .B(n_284), .Y(n_445) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g319 ( .A(n_281), .B(n_320), .Y(n_319) );
NAND2x1_ASAP7_75t_L g334 ( .A(n_281), .B(n_335), .Y(n_334) );
BUFx2_ASAP7_75t_L g403 ( .A(n_281), .Y(n_403) );
NAND2xp33_ASAP7_75t_R g386 ( .A(n_282), .B(n_309), .Y(n_386) );
AND2x2_ASAP7_75t_L g402 ( .A(n_282), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g468 ( .A(n_282), .Y(n_468) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx2_ASAP7_75t_L g295 ( .A(n_283), .Y(n_295) );
INVx1_ASAP7_75t_L g327 ( .A(n_283), .Y(n_327) );
INVx2_ASAP7_75t_L g394 ( .A(n_283), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_284), .B(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_286), .B(n_289), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g316 ( .A(n_287), .B(n_317), .Y(n_316) );
BUFx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g303 ( .A(n_290), .B(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_L g474 ( .A(n_290), .B(n_365), .Y(n_474) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AND2x2_ASAP7_75t_L g355 ( .A(n_292), .B(n_300), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g322 ( .A(n_298), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g425 ( .A(n_299), .Y(n_425) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g483 ( .A(n_302), .Y(n_483) );
INVx1_ASAP7_75t_L g311 ( .A(n_303), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_304), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g381 ( .A(n_304), .B(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g428 ( .A(n_304), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_304), .B(n_378), .Y(n_477) );
NOR3xp33_ASAP7_75t_L g305 ( .A(n_306), .B(n_312), .C(n_329), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_307), .B(n_311), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
AND2x2_ASAP7_75t_L g343 ( .A(n_309), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g436 ( .A(n_309), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_315), .B1(n_321), .B2(n_325), .Y(n_312) );
NAND3x2_ASAP7_75t_L g455 ( .A(n_313), .B(n_456), .C(n_457), .Y(n_455) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
NAND2x1_ASAP7_75t_L g395 ( .A(n_317), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g367 ( .A(n_319), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g439 ( .A(n_319), .Y(n_439) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g491 ( .A(n_323), .B(n_424), .Y(n_491) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g353 ( .A(n_324), .Y(n_353) );
NOR2x1p5_ASAP7_75t_SL g400 ( .A(n_326), .B(n_328), .Y(n_400) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g344 ( .A(n_327), .Y(n_344) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_327), .Y(n_446) );
OAI22xp33_ASAP7_75t_SL g329 ( .A1(n_330), .A2(n_336), .B1(n_342), .B2(n_345), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g489 ( .A(n_332), .B(n_436), .Y(n_489) );
INVxp67_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
OR2x6_ASAP7_75t_L g409 ( .A(n_334), .B(n_410), .Y(n_409) );
NOR2xp33_ASAP7_75t_SL g336 ( .A(n_337), .B(n_341), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g391 ( .A(n_338), .Y(n_391) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_343), .A2(n_459), .B1(n_464), .B2(n_466), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_343), .A2(n_437), .B1(n_494), .B2(n_495), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_343), .B(n_491), .Y(n_498) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR2x1_ASAP7_75t_L g349 ( .A(n_350), .B(n_383), .Y(n_349) );
NAND3xp33_ASAP7_75t_SL g350 ( .A(n_351), .B(n_361), .C(n_373), .Y(n_350) );
AO21x1_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B(n_356), .Y(n_351) );
INVx1_ASAP7_75t_L g453 ( .A(n_352), .Y(n_453) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
AOI32xp33_ASAP7_75t_L g473 ( .A1(n_357), .A2(n_474), .A3(n_475), .B1(n_476), .B2(n_478), .Y(n_473) );
BUFx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx2_ASAP7_75t_L g456 ( .A(n_360), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_366), .B1(n_369), .B2(n_372), .Y(n_361) );
INVxp67_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g389 ( .A(n_365), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_365), .B(n_397), .Y(n_398) );
AOI22xp33_ASAP7_75t_SL g373 ( .A1(n_366), .A2(n_374), .B1(n_376), .B2(n_380), .Y(n_373) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g470 ( .A(n_368), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI322xp33_ASAP7_75t_L g482 ( .A1(n_370), .A2(n_463), .A3(n_483), .B1(n_484), .B2(n_488), .C1(n_489), .C2(n_490), .Y(n_482) );
INVx2_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g502 ( .A(n_371), .B(n_391), .Y(n_502) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g463 ( .A(n_379), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_380), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g420 ( .A(n_382), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_406), .Y(n_383) );
AOI211xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .B(n_392), .C(n_401), .Y(n_384) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI22xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .B1(n_398), .B2(n_399), .Y(n_392) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_397), .B(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_397), .B(n_433), .Y(n_496) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_404), .Y(n_401) );
INVxp67_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_412), .B(n_413), .Y(n_406) );
NAND2x1_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
NOR2x1_ASAP7_75t_SL g435 ( .A(n_410), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g457 ( .A(n_410), .Y(n_457) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g472 ( .A(n_412), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .B1(n_419), .B2(n_421), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g475 ( .A(n_415), .Y(n_475) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NOR3x1_ASAP7_75t_L g422 ( .A(n_423), .B(n_447), .C(n_469), .Y(n_422) );
OAI211xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B(n_434), .C(n_443), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g441 ( .A(n_428), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_429), .B(n_431), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI21xp5_ASAP7_75t_SL g434 ( .A1(n_435), .A2(n_437), .B(n_440), .Y(n_434) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVxp67_ASAP7_75t_L g488 ( .A(n_438), .Y(n_488) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_455), .B(n_458), .Y(n_447) );
NOR3xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_453), .C(n_454), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_467), .B(n_468), .Y(n_466) );
OAI21xp5_ASAP7_75t_SL g469 ( .A1(n_470), .A2(n_472), .B(n_473), .Y(n_469) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NOR3xp33_ASAP7_75t_L g481 ( .A(n_482), .B(n_492), .C(n_497), .Y(n_481) );
NAND2x1p5_ASAP7_75t_L g484 ( .A(n_485), .B(n_487), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp33_ASAP7_75t_SL g497 ( .A(n_498), .B(n_499), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OAI21x1_ASAP7_75t_SL g509 ( .A1(n_510), .A2(n_516), .B(n_862), .Y(n_509) );
INVx4_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x6_ASAP7_75t_SL g511 ( .A(n_512), .B(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
XNOR2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_521), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AOI21x1_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_528), .B(n_530), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
INVx8_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx12f_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
BUFx8_ASAP7_75t_SL g532 ( .A(n_526), .Y(n_532) );
AND2x2_ASAP7_75t_L g870 ( .A(n_526), .B(n_871), .Y(n_870) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx2_ASAP7_75t_L g883 ( .A(n_527), .Y(n_883) );
NOR2x1_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
AND3x4_ASAP7_75t_L g533 ( .A(n_534), .B(n_759), .C(n_837), .Y(n_533) );
NOR2x1_ASAP7_75t_L g534 ( .A(n_535), .B(n_702), .Y(n_534) );
NAND3xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_649), .C(n_672), .Y(n_535) );
AOI221x1_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_583), .B1(n_605), .B2(n_614), .C(n_625), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_560), .Y(n_537) );
AND2x4_ASAP7_75t_L g739 ( .A(n_538), .B(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_551), .Y(n_539) );
INVx2_ASAP7_75t_L g698 ( .A(n_540), .Y(n_698) );
INVx1_ASAP7_75t_L g725 ( .A(n_540), .Y(n_725) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g608 ( .A(n_541), .Y(n_608) );
AND2x4_ASAP7_75t_L g676 ( .A(n_541), .B(n_609), .Y(n_676) );
AO31x2_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .A3(n_548), .B(n_549), .Y(n_541) );
AO31x2_ASAP7_75t_L g599 ( .A1(n_542), .A2(n_570), .A3(n_600), .B(n_603), .Y(n_599) );
AO31x2_ASAP7_75t_L g552 ( .A1(n_548), .A2(n_553), .A3(n_556), .B(n_558), .Y(n_552) );
INVx1_ASAP7_75t_L g758 ( .A(n_551), .Y(n_758) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g609 ( .A(n_552), .Y(n_609) );
AND2x4_ASAP7_75t_L g647 ( .A(n_552), .B(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g667 ( .A(n_552), .B(n_573), .Y(n_667) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_552), .Y(n_719) );
INVx1_ASAP7_75t_L g812 ( .A(n_552), .Y(n_812) );
AND2x2_ASAP7_75t_L g858 ( .A(n_552), .B(n_562), .Y(n_858) );
AO31x2_ASAP7_75t_L g617 ( .A1(n_556), .A2(n_580), .A3(n_618), .B(n_623), .Y(n_617) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_SL g596 ( .A(n_557), .Y(n_596) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_561), .B(n_724), .Y(n_723) );
NAND2x1_ASAP7_75t_L g728 ( .A(n_561), .B(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g852 ( .A(n_561), .B(n_750), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_561), .B(n_806), .Y(n_856) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_573), .Y(n_561) );
INVx4_ASAP7_75t_SL g611 ( .A(n_562), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_562), .B(n_613), .Y(n_660) );
BUFx2_ASAP7_75t_L g744 ( .A(n_562), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_562), .B(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g613 ( .A(n_573), .Y(n_613) );
INVx2_ASAP7_75t_L g648 ( .A(n_573), .Y(n_648) );
AND2x2_ASAP7_75t_L g650 ( .A(n_573), .B(n_608), .Y(n_650) );
INVx1_ASAP7_75t_L g675 ( .A(n_573), .Y(n_675) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_573), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_573), .B(n_758), .Y(n_789) );
INVxp67_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVxp67_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g833 ( .A(n_585), .B(n_834), .Y(n_833) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_598), .Y(n_585) );
AND2x4_ASAP7_75t_L g629 ( .A(n_586), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g690 ( .A(n_586), .B(n_634), .Y(n_690) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx2_ASAP7_75t_L g776 ( .A(n_587), .Y(n_776) );
OAI21x1_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B(n_597), .Y(n_587) );
OAI21x1_ASAP7_75t_L g663 ( .A1(n_588), .A2(n_589), .B(n_597), .Y(n_663) );
OAI21x1_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_593), .B(n_596), .Y(n_589) );
AND2x4_ASAP7_75t_L g688 ( .A(n_598), .B(n_617), .Y(n_688) );
INVx3_ASAP7_75t_L g711 ( .A(n_598), .Y(n_711) );
INVx2_ASAP7_75t_L g732 ( .A(n_598), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_598), .B(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_598), .B(n_633), .Y(n_826) );
INVx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g616 ( .A(n_599), .B(n_617), .Y(n_616) );
BUFx2_ASAP7_75t_L g628 ( .A(n_599), .Y(n_628) );
AND2x2_ASAP7_75t_L g705 ( .A(n_599), .B(n_630), .Y(n_705) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_610), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx3_ASAP7_75t_L g683 ( .A(n_608), .Y(n_683) );
AND2x2_ASAP7_75t_L g718 ( .A(n_608), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g787 ( .A(n_608), .B(n_611), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_609), .B(n_611), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g749 ( .A(n_610), .B(n_750), .Y(n_749) );
AND2x4_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx2_ASAP7_75t_L g646 ( .A(n_611), .Y(n_646) );
AND2x2_ASAP7_75t_L g674 ( .A(n_611), .B(n_675), .Y(n_674) );
OR2x2_ASAP7_75t_L g692 ( .A(n_611), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g734 ( .A(n_611), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_611), .B(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g795 ( .A(n_611), .Y(n_795) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_616), .B(n_662), .Y(n_661) );
AND2x4_ASAP7_75t_SL g669 ( .A(n_616), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g748 ( .A(n_616), .B(n_632), .Y(n_748) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_616), .Y(n_783) );
INVx2_ASAP7_75t_L g800 ( .A(n_616), .Y(n_800) );
INVx2_ASAP7_75t_L g630 ( .A(n_617), .Y(n_630) );
OR2x2_ASAP7_75t_L g680 ( .A(n_617), .B(n_671), .Y(n_680) );
INVx1_ASAP7_75t_L g701 ( .A(n_617), .Y(n_701) );
BUFx2_ASAP7_75t_L g716 ( .A(n_617), .Y(n_716) );
OR2x2_ASAP7_75t_L g785 ( .A(n_617), .B(n_635), .Y(n_785) );
AOI21xp5_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_631), .B(n_643), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_L g751 ( .A1(n_626), .A2(n_707), .B(n_752), .C(n_755), .Y(n_751) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g651 ( .A(n_627), .B(n_652), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_627), .A2(n_685), .B1(n_851), .B2(n_852), .Y(n_850) );
AND2x4_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx1_ASAP7_75t_L g642 ( .A(n_629), .Y(n_642) );
AND2x4_ASAP7_75t_L g770 ( .A(n_629), .B(n_679), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_629), .B(n_825), .Y(n_824) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_642), .Y(n_631) );
INVx1_ASAP7_75t_L g652 ( .A(n_632), .Y(n_652) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x4_ASAP7_75t_L g670 ( .A(n_633), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_634), .B(n_663), .Y(n_713) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g662 ( .A(n_635), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g679 ( .A(n_635), .Y(n_679) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_635), .Y(n_754) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
AND2x2_ASAP7_75t_L g665 ( .A(n_645), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_646), .B(n_725), .Y(n_764) );
INVx2_ASAP7_75t_L g656 ( .A(n_647), .Y(n_656) );
AND2x2_ASAP7_75t_L g733 ( .A(n_647), .B(n_734), .Y(n_733) );
NAND2x1p5_ASAP7_75t_L g778 ( .A(n_647), .B(n_697), .Y(n_778) );
AND2x2_ASAP7_75t_L g815 ( .A(n_647), .B(n_787), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B(n_653), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_661), .B1(n_664), .B2(n_668), .Y(n_653) );
NOR2x1_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g859 ( .A(n_656), .Y(n_859) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g699 ( .A(n_662), .Y(n_699) );
AND2x2_ASAP7_75t_L g726 ( .A(n_662), .B(n_711), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_662), .B(n_705), .Y(n_796) );
AND2x4_ASAP7_75t_L g842 ( .A(n_662), .B(n_688), .Y(n_842) );
INVx1_ASAP7_75t_L g671 ( .A(n_663), .Y(n_671) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x4_ASAP7_75t_L g848 ( .A(n_666), .B(n_744), .Y(n_848) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OR2x2_ASAP7_75t_L g781 ( .A(n_667), .B(n_782), .Y(n_781) );
OR2x2_ASAP7_75t_L g809 ( .A(n_667), .B(n_683), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_668), .B(n_841), .Y(n_840) );
INVx3_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g790 ( .A(n_670), .B(n_791), .Y(n_790) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_677), .B1(n_681), .B2(n_685), .C(n_691), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
INVx1_ASAP7_75t_L g707 ( .A(n_674), .Y(n_707) );
AND2x2_ASAP7_75t_L g831 ( .A(n_674), .B(n_697), .Y(n_831) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_675), .Y(n_695) );
INVx3_ASAP7_75t_L g693 ( .A(n_676), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_676), .B(n_743), .Y(n_742) );
AND2x4_ASAP7_75t_L g765 ( .A(n_676), .B(n_766), .Y(n_765) );
NOR2xp67_ASAP7_75t_SL g677 ( .A(n_678), .B(n_680), .Y(n_677) );
AND2x2_ASAP7_75t_L g704 ( .A(n_678), .B(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_678), .B(n_711), .Y(n_773) );
AOI322xp5_ASAP7_75t_L g779 ( .A1(n_678), .A2(n_765), .A3(n_780), .B1(n_783), .B2(n_784), .C1(n_786), .C2(n_790), .Y(n_779) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g721 ( .A(n_679), .B(n_688), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_680), .B(n_732), .Y(n_731) );
NOR2x1_ASAP7_75t_L g829 ( .A(n_680), .B(n_830), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_681), .A2(n_823), .B1(n_827), .B2(n_831), .Y(n_822) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OR2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx4_ASAP7_75t_L g806 ( .A(n_683), .Y(n_806) );
OR2x2_ASAP7_75t_L g836 ( .A(n_683), .B(n_811), .Y(n_836) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_689), .Y(n_686) );
INVx2_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g849 ( .A(n_688), .Y(n_849) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_689), .B(n_715), .Y(n_736) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI211x1_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_694), .B(n_699), .C(n_700), .Y(n_691) );
INVx2_ASAP7_75t_L g729 ( .A(n_693), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g756 ( .A(n_697), .Y(n_756) );
NAND2x1_ASAP7_75t_L g847 ( .A(n_697), .B(n_848), .Y(n_847) );
INVx3_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g753 ( .A(n_698), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g818 ( .A(n_700), .Y(n_818) );
BUFx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_720), .C(n_735), .Y(n_702) );
OAI211xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_706), .B(n_708), .C(n_718), .Y(n_703) );
INVx1_ASAP7_75t_L g717 ( .A(n_704), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_705), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g775 ( .A(n_705), .B(n_776), .Y(n_775) );
NAND2xp33_ASAP7_75t_L g798 ( .A(n_705), .B(n_746), .Y(n_798) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_717), .Y(n_708) );
INVx1_ASAP7_75t_L g844 ( .A(n_709), .Y(n_844) );
NAND2x1p5_ASAP7_75t_L g709 ( .A(n_710), .B(n_714), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx2_ASAP7_75t_L g791 ( .A(n_711), .Y(n_791) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g746 ( .A(n_713), .Y(n_746) );
INVxp67_ASAP7_75t_SL g821 ( .A(n_713), .Y(n_821) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g750 ( .A(n_719), .Y(n_750) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B1(n_726), .B2(n_727), .C(n_730), .Y(n_720) );
INVxp67_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g782 ( .A(n_725), .Y(n_782) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .Y(n_730) );
INVx1_ASAP7_75t_L g768 ( .A(n_732), .Y(n_768) );
NOR2x1p5_ASAP7_75t_L g784 ( .A(n_732), .B(n_785), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_733), .A2(n_772), .B(n_774), .Y(n_771) );
INVx1_ASAP7_75t_L g740 ( .A(n_734), .Y(n_740) );
AOI211xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B(n_741), .C(n_751), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_745), .B1(n_747), .B2(n_749), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g830 ( .A(n_754), .Y(n_830) );
OR2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
NOR3xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_792), .C(n_813), .Y(n_759) );
NAND3xp33_ASAP7_75t_SL g760 ( .A(n_761), .B(n_771), .C(n_779), .Y(n_760) );
OAI21xp33_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_765), .B(n_767), .Y(n_761) );
INVxp67_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
AND2x2_ASAP7_75t_L g861 ( .A(n_768), .B(n_829), .Y(n_861) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OAI21xp5_ASAP7_75t_L g807 ( .A1(n_770), .A2(n_808), .B(n_810), .Y(n_807) );
INVxp67_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_777), .Y(n_774) );
OR2x2_ASAP7_75t_L g799 ( .A(n_776), .B(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g834 ( .A(n_785), .Y(n_834) );
AND2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_788), .Y(n_851) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
OR2x2_ASAP7_75t_L g794 ( .A(n_789), .B(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g804 ( .A(n_789), .Y(n_804) );
OAI221xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_796), .B1(n_797), .B2(n_801), .C(n_807), .Y(n_792) );
OAI21xp5_ASAP7_75t_L g838 ( .A1(n_793), .A2(n_839), .B(n_843), .Y(n_838) );
BUFx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
AOI32xp33_ASAP7_75t_L g832 ( .A1(n_795), .A2(n_806), .A3(n_833), .B1(n_834), .B2(n_835), .Y(n_832) );
AND2x2_ASAP7_75t_SL g797 ( .A(n_798), .B(n_799), .Y(n_797) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_808), .B(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OAI211xp5_ASAP7_75t_SL g813 ( .A1(n_814), .A2(n_816), .B(n_822), .C(n_832), .Y(n_813) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
AND2x4_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .Y(n_817) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
NOR3xp33_ASAP7_75t_L g837 ( .A(n_838), .B(n_845), .C(n_853), .Y(n_837) );
INVxp33_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
OAI21xp33_ASAP7_75t_SL g845 ( .A1(n_846), .A2(n_849), .B(n_850), .Y(n_845) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
AOI21xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_857), .B(n_860), .Y(n_853) );
INVxp67_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
NOR2xp33_ASAP7_75t_SL g857 ( .A(n_858), .B(n_859), .Y(n_857) );
INVx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
NOR2xp33_ASAP7_75t_SL g862 ( .A(n_863), .B(n_872), .Y(n_862) );
NOR2xp33_ASAP7_75t_L g863 ( .A(n_864), .B(n_865), .Y(n_863) );
BUFx6f_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
BUFx10_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
NOR2xp33_ASAP7_75t_SL g872 ( .A(n_873), .B(n_874), .Y(n_872) );
INVx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
CKINVDCx10_ASAP7_75t_R g877 ( .A(n_878), .Y(n_877) );
CKINVDCx11_ASAP7_75t_R g894 ( .A(n_878), .Y(n_894) );
OR2x6_ASAP7_75t_L g878 ( .A(n_879), .B(n_886), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
NOR2x1p5_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_883), .B(n_884), .Y(n_882) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_888), .B(n_889), .Y(n_887) );
INVxp33_ASAP7_75t_SL g889 ( .A(n_890), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g891 ( .A(n_892), .Y(n_891) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_893), .Y(n_892) );
CKINVDCx20_ASAP7_75t_R g893 ( .A(n_894), .Y(n_893) );
endmodule