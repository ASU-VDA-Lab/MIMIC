module fake_jpeg_23568_n_334 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_47),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_9),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_52),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_59),
.B(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_27),
.B1(n_22),
.B2(n_24),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_75),
.B1(n_78),
.B2(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_19),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_11),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_70),
.Y(n_109)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_72),
.Y(n_113)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_73),
.Y(n_116)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_20),
.B1(n_36),
.B2(n_34),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx4f_ASAP7_75t_SL g99 ( 
.A(n_76),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_20),
.B1(n_36),
.B2(n_33),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_19),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_79),
.B(n_86),
.Y(n_115)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_43),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_38),
.C(n_37),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_28),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_20),
.B1(n_34),
.B2(n_17),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_41),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_44),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_52),
.C(n_44),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_37),
.B1(n_35),
.B2(n_18),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_94),
.A2(n_98),
.B1(n_110),
.B2(n_61),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_9),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_71),
.A2(n_34),
.B1(n_17),
.B2(n_33),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_41),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_101),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_41),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_46),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_102),
.B(n_104),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_75),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_17),
.B1(n_33),
.B2(n_35),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_106),
.A2(n_118),
.B1(n_83),
.B2(n_61),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_18),
.B1(n_25),
.B2(n_21),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_120),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_57),
.B(n_46),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_62),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_69),
.B(n_21),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_117),
.B(n_83),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_65),
.A2(n_25),
.B1(n_22),
.B2(n_26),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_58),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_123),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_124),
.B(n_128),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_127),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_149),
.C(n_108),
.Y(n_165)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_130),
.Y(n_166)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_134),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_90),
.B(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_133),
.B(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_93),
.A2(n_67),
.B1(n_58),
.B2(n_65),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_135),
.A2(n_156),
.B1(n_103),
.B2(n_107),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_13),
.Y(n_178)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_0),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_153),
.B(n_116),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_96),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_144),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_101),
.A2(n_65),
.B1(n_67),
.B2(n_80),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_111),
.B1(n_120),
.B2(n_121),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_143),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_148),
.A2(n_27),
.B1(n_31),
.B2(n_26),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_91),
.B(n_104),
.C(n_109),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_151),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_91),
.B(n_0),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_89),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_122),
.B(n_108),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_160),
.A2(n_167),
.B(n_24),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_161),
.A2(n_183),
.B1(n_188),
.B2(n_191),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_157),
.A2(n_51),
.B1(n_87),
.B2(n_73),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_162),
.A2(n_164),
.B1(n_176),
.B2(n_184),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_145),
.A2(n_87),
.B1(n_60),
.B2(n_72),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_159),
.C(n_66),
.Y(n_204)
);

O2A1O1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_99),
.B(n_62),
.C(n_48),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_178),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_145),
.B(n_92),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_173),
.B(n_12),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_149),
.A2(n_113),
.B1(n_95),
.B2(n_119),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_126),
.A2(n_119),
.B1(n_46),
.B2(n_48),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_156),
.A2(n_128),
.B1(n_140),
.B2(n_136),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_187),
.B(n_189),
.Y(n_224)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_192),
.B1(n_29),
.B2(n_26),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_140),
.A2(n_31),
.B1(n_29),
.B2(n_27),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_153),
.A2(n_31),
.B1(n_29),
.B2(n_27),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_66),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_152),
.B(n_147),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_194),
.A2(n_199),
.B(n_211),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_136),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_198),
.Y(n_231)
);

NOR2x1_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_159),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_L g246 ( 
.A(n_197),
.B(n_185),
.C(n_13),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_137),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_201),
.Y(n_226)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_203),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_150),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_214),
.C(n_220),
.Y(n_236)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_210),
.Y(n_240)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_144),
.Y(n_208)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_127),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_130),
.B(n_129),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_222),
.B(n_210),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_132),
.C(n_146),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_160),
.B(n_31),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_216),
.A2(n_186),
.B1(n_189),
.B2(n_185),
.Y(n_230)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_179),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_219),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_29),
.C(n_26),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_191),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_233),
.C(n_237),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_230),
.A2(n_244),
.B1(n_247),
.B2(n_217),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_174),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_232),
.A2(n_238),
.B(n_171),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_187),
.C(n_192),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_177),
.C(n_168),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_245),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_224),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_242),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_211),
.A2(n_168),
.B1(n_177),
.B2(n_180),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_243),
.A2(n_217),
.B1(n_220),
.B2(n_215),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_203),
.A2(n_181),
.B1(n_186),
.B2(n_179),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_246),
.A2(n_235),
.B1(n_248),
.B2(n_241),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_213),
.A2(n_171),
.B1(n_180),
.B2(n_24),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_213),
.B1(n_222),
.B2(n_216),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_250),
.A2(n_252),
.B1(n_261),
.B2(n_230),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_251),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_197),
.B1(n_194),
.B2(n_214),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_198),
.Y(n_254)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_259),
.Y(n_276)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_195),
.C(n_202),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_233),
.C(n_1),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_263),
.A2(n_266),
.B(n_268),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_24),
.B1(n_22),
.B2(n_0),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_264),
.A2(n_240),
.B1(n_249),
.B2(n_234),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_227),
.Y(n_281)
);

AOI21xp33_ASAP7_75t_L g266 ( 
.A1(n_231),
.A2(n_7),
.B(n_2),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_250),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_234),
.A2(n_1),
.B(n_2),
.Y(n_268)
);

OA21x2_ASAP7_75t_L g269 ( 
.A1(n_232),
.A2(n_1),
.B(n_3),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_10),
.B(n_3),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_267),
.B1(n_258),
.B2(n_260),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_259),
.A2(n_232),
.B1(n_236),
.B2(n_237),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_252),
.B1(n_284),
.B2(n_261),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_256),
.B(n_251),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_277),
.Y(n_297)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_257),
.B(n_225),
.Y(n_277)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_279),
.Y(n_296)
);

AO21x1_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_282),
.B(n_269),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_227),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_254),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_268),
.C(n_263),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_5),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_287),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_5),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_257),
.Y(n_288)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_276),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_289),
.B(n_292),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_290),
.A2(n_293),
.B1(n_275),
.B2(n_286),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_300),
.C(n_278),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_295),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_279),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_298),
.A2(n_270),
.B(n_280),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_262),
.C(n_283),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_287),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_306),
.Y(n_317)
);

OAI21xp33_ASAP7_75t_SL g315 ( 
.A1(n_303),
.A2(n_282),
.B(n_265),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_305),
.B(n_299),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_280),
.C(n_270),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_295),
.B1(n_292),
.B2(n_269),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_297),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_264),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_278),
.C(n_271),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_311),
.A2(n_285),
.B(n_299),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_310),
.A2(n_294),
.B1(n_296),
.B2(n_298),
.Y(n_312)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_312),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_316),
.C(n_302),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_314),
.A2(n_307),
.B1(n_309),
.B2(n_313),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_318),
.B(n_319),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_311),
.B(n_306),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_321),
.B(n_322),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_317),
.A2(n_305),
.B(n_7),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_7),
.Y(n_325)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_325),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_8),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_327),
.A2(n_324),
.B(n_8),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_329),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_326),
.Y(n_331)
);

AOI221xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_8),
.B1(n_10),
.B2(n_15),
.C(n_16),
.Y(n_332)
);

XNOR2x2_ASAP7_75t_SL g333 ( 
.A(n_332),
.B(n_16),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_1),
.Y(n_334)
);


endmodule