module fake_aes_7845_n_879 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_879);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_879;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_163;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_769;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_844;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_482;
wire n_394;
wire n_235;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_876;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_225;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_836;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g103 ( .A(n_67), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_69), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_61), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_26), .Y(n_106) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_101), .Y(n_107) );
BUFx2_ASAP7_75t_L g108 ( .A(n_97), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_10), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_77), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_25), .Y(n_111) );
INVx1_ASAP7_75t_SL g112 ( .A(n_23), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_87), .Y(n_113) );
BUFx10_ASAP7_75t_L g114 ( .A(n_62), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_96), .Y(n_115) );
INVx2_ASAP7_75t_SL g116 ( .A(n_12), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_38), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_7), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_90), .Y(n_119) );
INVxp67_ASAP7_75t_L g120 ( .A(n_16), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_52), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_36), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_2), .Y(n_123) );
BUFx10_ASAP7_75t_L g124 ( .A(n_49), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_95), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_98), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_41), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_81), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_76), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_60), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_9), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_46), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_93), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_89), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_58), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_15), .Y(n_137) );
CKINVDCx16_ASAP7_75t_R g138 ( .A(n_39), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_78), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_2), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_30), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_92), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_27), .Y(n_143) );
BUFx3_ASAP7_75t_L g144 ( .A(n_51), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_26), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_21), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_140), .Y(n_147) );
INVx5_ASAP7_75t_L g148 ( .A(n_104), .Y(n_148) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_120), .Y(n_149) );
INVx5_ASAP7_75t_L g150 ( .A(n_104), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_108), .B(n_0), .Y(n_151) );
INVxp67_ASAP7_75t_L g152 ( .A(n_108), .Y(n_152) );
INVx4_ASAP7_75t_L g153 ( .A(n_111), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_104), .Y(n_154) );
INVx5_ASAP7_75t_L g155 ( .A(n_136), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_138), .B(n_0), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_138), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_140), .Y(n_158) );
INVx5_ASAP7_75t_L g159 ( .A(n_136), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_144), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_140), .Y(n_161) );
XOR2xp5_ASAP7_75t_L g162 ( .A(n_106), .B(n_1), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_144), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_144), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_116), .B(n_1), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_116), .B(n_3), .Y(n_166) );
BUFx12f_ASAP7_75t_L g167 ( .A(n_114), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_136), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_103), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_152), .A2(n_116), .B1(n_120), .B2(n_143), .Y(n_170) );
AO22x2_ASAP7_75t_L g171 ( .A1(n_162), .A2(n_129), .B1(n_119), .B2(n_126), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_152), .B(n_114), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_149), .B(n_114), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_166), .A2(n_123), .B1(n_122), .B2(n_117), .Y(n_174) );
AO22x2_ASAP7_75t_L g175 ( .A1(n_162), .A2(n_129), .B1(n_119), .B2(n_126), .Y(n_175) );
OAI22xp33_ASAP7_75t_SL g176 ( .A1(n_157), .A2(n_112), .B1(n_141), .B2(n_145), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_167), .B(n_114), .Y(n_177) );
OAI22xp33_ASAP7_75t_SL g178 ( .A1(n_157), .A2(n_112), .B1(n_145), .B2(n_109), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_166), .A2(n_146), .B1(n_132), .B2(n_109), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_148), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_167), .B(n_107), .Y(n_182) );
NAND3x1_ASAP7_75t_L g183 ( .A(n_156), .B(n_146), .C(n_132), .Y(n_183) );
AO22x2_ASAP7_75t_L g184 ( .A1(n_162), .A2(n_166), .B1(n_156), .B2(n_165), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_149), .B(n_124), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_153), .Y(n_186) );
OAI22xp33_ASAP7_75t_SL g187 ( .A1(n_165), .A2(n_103), .B1(n_130), .B2(n_135), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_167), .B(n_124), .Y(n_188) );
OR2x2_ASAP7_75t_L g189 ( .A(n_156), .B(n_111), .Y(n_189) );
AO22x2_ASAP7_75t_L g190 ( .A1(n_166), .A2(n_130), .B1(n_131), .B2(n_134), .Y(n_190) );
OAI22xp33_ASAP7_75t_SL g191 ( .A1(n_165), .A2(n_131), .B1(n_135), .B2(n_134), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_156), .A2(n_105), .B1(n_139), .B2(n_137), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_167), .B(n_124), .Y(n_193) );
AO22x2_ASAP7_75t_L g194 ( .A1(n_166), .A2(n_124), .B1(n_4), .B2(n_5), .Y(n_194) );
OAI22xp33_ASAP7_75t_SL g195 ( .A1(n_151), .A2(n_142), .B1(n_133), .B2(n_128), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_148), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_166), .B(n_111), .Y(n_197) );
OAI22xp33_ASAP7_75t_L g198 ( .A1(n_151), .A2(n_111), .B1(n_118), .B2(n_121), .Y(n_198) );
OA22x2_ASAP7_75t_L g199 ( .A1(n_166), .A2(n_127), .B1(n_125), .B2(n_115), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_169), .B(n_111), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_148), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_169), .A2(n_118), .B1(n_111), .B2(n_113), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_169), .A2(n_118), .B1(n_110), .B2(n_5), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_169), .B(n_118), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_147), .B(n_118), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_147), .B(n_118), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_147), .B(n_3), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_154), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_158), .B(n_4), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_154), .Y(n_210) );
AO22x2_ASAP7_75t_L g211 ( .A1(n_154), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_158), .B(n_6), .Y(n_212) );
AO22x2_ASAP7_75t_L g213 ( .A1(n_154), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_158), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_161), .B(n_11), .Y(n_215) );
AO22x2_ASAP7_75t_L g216 ( .A1(n_161), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_197), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_197), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_208), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_208), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_208), .Y(n_221) );
OR2x2_ASAP7_75t_L g222 ( .A(n_192), .B(n_161), .Y(n_222) );
XOR2xp5_ASAP7_75t_L g223 ( .A(n_184), .B(n_14), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_172), .B(n_148), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_210), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_210), .Y(n_226) );
NOR2x1p5_ASAP7_75t_L g227 ( .A(n_173), .B(n_153), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_210), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_173), .B(n_148), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_200), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_200), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_185), .B(n_148), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_188), .B(n_148), .Y(n_233) );
XOR2xp5_ASAP7_75t_L g234 ( .A(n_184), .B(n_16), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_204), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_181), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_204), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_185), .B(n_17), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_172), .B(n_148), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_181), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_182), .B(n_148), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_207), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_207), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_196), .Y(n_244) );
XOR2xp5_ASAP7_75t_L g245 ( .A(n_184), .B(n_17), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_201), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_209), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_189), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_209), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_177), .B(n_148), .Y(n_250) );
NOR2xp67_ASAP7_75t_L g251 ( .A(n_170), .B(n_148), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_188), .B(n_150), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_193), .B(n_150), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_212), .Y(n_254) );
NAND2xp33_ASAP7_75t_SL g255 ( .A(n_193), .B(n_160), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_212), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_215), .Y(n_257) );
OR2x2_ASAP7_75t_L g258 ( .A(n_189), .B(n_18), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_201), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_174), .Y(n_260) );
INVxp67_ASAP7_75t_SL g261 ( .A(n_190), .Y(n_261) );
OR2x2_ASAP7_75t_L g262 ( .A(n_180), .B(n_18), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_215), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_205), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g265 ( .A1(n_179), .A2(n_153), .B(n_150), .Y(n_265) );
INVx2_ASAP7_75t_SL g266 ( .A(n_190), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_205), .B(n_150), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_190), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_190), .B(n_150), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_184), .B(n_150), .Y(n_270) );
NOR2xp33_ASAP7_75t_SL g271 ( .A(n_176), .B(n_150), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_206), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_206), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_194), .B(n_150), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_196), .Y(n_275) );
INVxp67_ASAP7_75t_SL g276 ( .A(n_183), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_187), .B(n_150), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_194), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_248), .B(n_183), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_267), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_248), .B(n_191), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_242), .B(n_178), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_244), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_239), .B(n_195), .Y(n_284) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_274), .A2(n_199), .B(n_203), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_242), .B(n_199), .Y(n_286) );
BUFx4f_ASAP7_75t_L g287 ( .A(n_266), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_266), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_270), .B(n_171), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_267), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_268), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_270), .B(n_171), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_268), .B(n_171), .Y(n_293) );
OAI21xp33_ASAP7_75t_L g294 ( .A1(n_243), .A2(n_194), .B(n_199), .Y(n_294) );
BUFx8_ASAP7_75t_L g295 ( .A(n_269), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_261), .B(n_171), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_239), .B(n_175), .Y(n_297) );
AND2x2_ASAP7_75t_SL g298 ( .A(n_278), .B(n_214), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_239), .B(n_175), .Y(n_299) );
INVxp67_ASAP7_75t_L g300 ( .A(n_258), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_267), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_267), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_219), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_244), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_269), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_244), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_223), .B(n_175), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_239), .B(n_175), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_219), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_244), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_223), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_243), .B(n_194), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_232), .B(n_211), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_277), .A2(n_186), .B(n_179), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_258), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_217), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_247), .B(n_249), .Y(n_317) );
BUFx3_ASAP7_75t_L g318 ( .A(n_217), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_247), .B(n_198), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_220), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_234), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_232), .B(n_211), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_234), .A2(n_213), .B1(n_211), .B2(n_216), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_249), .B(n_150), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_254), .B(n_211), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_220), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_236), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_254), .B(n_150), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_236), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_291), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_325), .B(n_256), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_297), .B(n_245), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_303), .Y(n_333) );
INVx4_ASAP7_75t_L g334 ( .A(n_287), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_291), .Y(n_335) );
BUFx2_ASAP7_75t_SL g336 ( .A(n_291), .Y(n_336) );
OR2x6_ASAP7_75t_L g337 ( .A(n_293), .B(n_274), .Y(n_337) );
NOR2xp33_ASAP7_75t_SL g338 ( .A(n_287), .B(n_256), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_327), .Y(n_339) );
NAND2x1p5_ASAP7_75t_L g340 ( .A(n_291), .B(n_257), .Y(n_340) );
INVx2_ASAP7_75t_SL g341 ( .A(n_287), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_325), .B(n_257), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_316), .B(n_218), .Y(n_343) );
BUFx8_ASAP7_75t_L g344 ( .A(n_293), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_297), .B(n_245), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_297), .B(n_263), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_295), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_327), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_297), .B(n_263), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_307), .B(n_315), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_300), .B(n_276), .Y(n_351) );
NOR2xp33_ASAP7_75t_SL g352 ( .A(n_287), .B(n_251), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_325), .B(n_218), .Y(n_353) );
INVx3_ASAP7_75t_L g354 ( .A(n_287), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_327), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_325), .B(n_230), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_295), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_307), .B(n_238), .Y(n_358) );
AND2x2_ASAP7_75t_SL g359 ( .A(n_287), .B(n_238), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_327), .Y(n_360) );
INVxp67_ASAP7_75t_L g361 ( .A(n_288), .Y(n_361) );
INVxp67_ASAP7_75t_SL g362 ( .A(n_339), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_339), .Y(n_363) );
BUFx4f_ASAP7_75t_SL g364 ( .A(n_357), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_357), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_357), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_339), .Y(n_367) );
INVx2_ASAP7_75t_SL g368 ( .A(n_339), .Y(n_368) );
BUFx12f_ASAP7_75t_L g369 ( .A(n_347), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_347), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_339), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_357), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_348), .Y(n_373) );
BUFx2_ASAP7_75t_L g374 ( .A(n_357), .Y(n_374) );
BUFx8_ASAP7_75t_SL g375 ( .A(n_337), .Y(n_375) );
BUFx8_ASAP7_75t_L g376 ( .A(n_348), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_335), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_348), .B(n_293), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_348), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_344), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_348), .Y(n_381) );
INVx5_ASAP7_75t_L g382 ( .A(n_334), .Y(n_382) );
BUFx2_ASAP7_75t_SL g383 ( .A(n_355), .Y(n_383) );
BUFx3_ASAP7_75t_L g384 ( .A(n_344), .Y(n_384) );
INVx2_ASAP7_75t_SL g385 ( .A(n_355), .Y(n_385) );
INVxp67_ASAP7_75t_SL g386 ( .A(n_355), .Y(n_386) );
BUFx8_ASAP7_75t_L g387 ( .A(n_355), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_333), .B(n_293), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_344), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_355), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_367), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_376), .A2(n_323), .B1(n_307), .B2(n_298), .Y(n_392) );
AOI22xp33_ASAP7_75t_SL g393 ( .A1(n_364), .A2(n_311), .B1(n_307), .B2(n_321), .Y(n_393) );
CKINVDCx11_ASAP7_75t_R g394 ( .A(n_370), .Y(n_394) );
AOI22x1_ASAP7_75t_SL g395 ( .A1(n_389), .A2(n_321), .B1(n_260), .B2(n_311), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_362), .Y(n_396) );
BUFx3_ASAP7_75t_L g397 ( .A(n_376), .Y(n_397) );
BUFx10_ASAP7_75t_L g398 ( .A(n_371), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_367), .Y(n_399) );
BUFx12f_ASAP7_75t_L g400 ( .A(n_376), .Y(n_400) );
BUFx4f_ASAP7_75t_SL g401 ( .A(n_376), .Y(n_401) );
AOI22xp33_ASAP7_75t_SL g402 ( .A1(n_364), .A2(n_311), .B1(n_345), .B2(n_332), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_367), .Y(n_403) );
NAND2x1p5_ASAP7_75t_L g404 ( .A(n_382), .B(n_334), .Y(n_404) );
BUFx10_ASAP7_75t_L g405 ( .A(n_371), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_362), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_376), .A2(n_298), .B1(n_332), .B2(n_345), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_370), .Y(n_408) );
INVx5_ASAP7_75t_L g409 ( .A(n_382), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_364), .A2(n_345), .B1(n_332), .B2(n_359), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_388), .B(n_332), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_383), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_362), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_363), .B(n_360), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_369), .Y(n_415) );
AOI22xp33_ASAP7_75t_SL g416 ( .A1(n_376), .A2(n_345), .B1(n_359), .B2(n_344), .Y(n_416) );
BUFx4f_ASAP7_75t_L g417 ( .A(n_369), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_376), .A2(n_298), .B1(n_344), .B2(n_359), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_386), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_369), .Y(n_420) );
NAND2x1p5_ASAP7_75t_L g421 ( .A(n_382), .B(n_334), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_363), .Y(n_422) );
INVx8_ASAP7_75t_L g423 ( .A(n_382), .Y(n_423) );
INVx1_ASAP7_75t_SL g424 ( .A(n_383), .Y(n_424) );
CKINVDCx11_ASAP7_75t_R g425 ( .A(n_389), .Y(n_425) );
INVx6_ASAP7_75t_L g426 ( .A(n_376), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_367), .Y(n_427) );
OAI21xp5_ASAP7_75t_L g428 ( .A1(n_386), .A2(n_323), .B(n_294), .Y(n_428) );
INVx6_ASAP7_75t_L g429 ( .A(n_387), .Y(n_429) );
INVx8_ASAP7_75t_L g430 ( .A(n_382), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_367), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_383), .A2(n_323), .B1(n_359), .B2(n_358), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_387), .A2(n_298), .B1(n_344), .B2(n_359), .Y(n_433) );
BUFx2_ASAP7_75t_SL g434 ( .A(n_380), .Y(n_434) );
NOR2xp67_ASAP7_75t_L g435 ( .A(n_400), .B(n_363), .Y(n_435) );
OAI22xp5_ASAP7_75t_SL g436 ( .A1(n_408), .A2(n_384), .B1(n_380), .B2(n_369), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_414), .B(n_386), .Y(n_437) );
OAI21xp5_ASAP7_75t_SL g438 ( .A1(n_416), .A2(n_372), .B(n_366), .Y(n_438) );
BUFx2_ASAP7_75t_L g439 ( .A(n_400), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_392), .A2(n_298), .B1(n_387), .B2(n_300), .Y(n_440) );
OAI21xp33_ASAP7_75t_L g441 ( .A1(n_392), .A2(n_294), .B(n_213), .Y(n_441) );
BUFx2_ASAP7_75t_L g442 ( .A(n_400), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_396), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_398), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_401), .A2(n_387), .B1(n_380), .B2(n_384), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_410), .A2(n_387), .B1(n_380), .B2(n_384), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_418), .A2(n_358), .B1(n_380), .B2(n_384), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_397), .A2(n_387), .B1(n_384), .B2(n_344), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_394), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_396), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_425), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_433), .A2(n_358), .B1(n_374), .B2(n_366), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_397), .A2(n_387), .B1(n_374), .B2(n_372), .Y(n_453) );
AOI222xp33_ASAP7_75t_L g454 ( .A1(n_407), .A2(n_308), .B1(n_299), .B2(n_292), .C1(n_289), .C2(n_294), .Y(n_454) );
AOI22xp33_ASAP7_75t_SL g455 ( .A1(n_426), .A2(n_387), .B1(n_366), .B2(n_374), .Y(n_455) );
INVx4_ASAP7_75t_SL g456 ( .A(n_426), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_406), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_414), .B(n_371), .Y(n_458) );
BUFx2_ASAP7_75t_L g459 ( .A(n_397), .Y(n_459) );
AOI22xp33_ASAP7_75t_SL g460 ( .A1(n_426), .A2(n_372), .B1(n_366), .B2(n_374), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_432), .A2(n_372), .B1(n_365), .B2(n_292), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_402), .A2(n_365), .B1(n_289), .B2(n_292), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_426), .A2(n_358), .B1(n_383), .B2(n_382), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_406), .B(n_371), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_413), .B(n_373), .Y(n_465) );
OAI21xp33_ASAP7_75t_L g466 ( .A1(n_393), .A2(n_213), .B(n_216), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_413), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_419), .B(n_373), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_429), .A2(n_365), .B1(n_289), .B2(n_292), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_429), .A2(n_423), .B1(n_430), .B2(n_434), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_429), .A2(n_382), .B1(n_365), .B2(n_315), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_429), .A2(n_365), .B1(n_289), .B2(n_308), .Y(n_472) );
AOI22xp33_ASAP7_75t_SL g473 ( .A1(n_434), .A2(n_382), .B1(n_369), .B2(n_296), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_423), .A2(n_308), .B1(n_299), .B2(n_296), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_391), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_419), .B(n_373), .Y(n_476) );
OAI222xp33_ASAP7_75t_L g477 ( .A1(n_409), .A2(n_350), .B1(n_382), .B2(n_296), .C1(n_385), .C2(n_368), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_395), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_391), .B(n_373), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_423), .A2(n_299), .B1(n_308), .B2(n_296), .Y(n_480) );
OAI21xp33_ASAP7_75t_L g481 ( .A1(n_422), .A2(n_213), .B(n_216), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_398), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_391), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_411), .B(n_350), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_409), .B(n_350), .Y(n_485) );
AOI22xp33_ASAP7_75t_SL g486 ( .A1(n_423), .A2(n_382), .B1(n_295), .B2(n_299), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_398), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_399), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_423), .A2(n_295), .B1(n_284), .B2(n_350), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_395), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_399), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_412), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_409), .B(n_378), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_417), .A2(n_382), .B1(n_385), .B2(n_368), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_430), .A2(n_295), .B1(n_284), .B2(n_375), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_398), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_399), .B(n_368), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_417), .A2(n_382), .B1(n_385), .B2(n_368), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_430), .A2(n_295), .B1(n_375), .B2(n_337), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_430), .A2(n_295), .B1(n_337), .B2(n_382), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_417), .A2(n_368), .B1(n_385), .B2(n_379), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_405), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g503 ( .A1(n_430), .A2(n_216), .B1(n_385), .B2(n_381), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_415), .B(n_271), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_409), .A2(n_381), .B1(n_313), .B2(n_322), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_409), .A2(n_337), .B1(n_346), .B2(n_349), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_409), .B(n_378), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_447), .A2(n_417), .B1(n_428), .B2(n_337), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_440), .A2(n_441), .B1(n_452), .B2(n_466), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_458), .B(n_405), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_443), .Y(n_511) );
OAI221xp5_ASAP7_75t_L g512 ( .A1(n_503), .A2(n_222), .B1(n_282), .B2(n_262), .C(n_351), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_443), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_458), .B(n_405), .Y(n_514) );
AOI222xp33_ASAP7_75t_L g515 ( .A1(n_441), .A2(n_351), .B1(n_282), .B2(n_346), .C1(n_349), .C2(n_286), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_440), .A2(n_337), .B1(n_313), .B2(n_322), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_466), .A2(n_337), .B1(n_313), .B2(n_322), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_461), .A2(n_337), .B1(n_313), .B2(n_322), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_437), .B(n_403), .Y(n_519) );
OAI22xp33_ASAP7_75t_L g520 ( .A1(n_438), .A2(n_421), .B1(n_404), .B2(n_424), .Y(n_520) );
NOR2xp67_ASAP7_75t_L g521 ( .A(n_435), .B(n_403), .Y(n_521) );
OAI221xp5_ASAP7_75t_L g522 ( .A1(n_478), .A2(n_222), .B1(n_262), .B2(n_286), .C(n_281), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_446), .A2(n_337), .B1(n_378), .B2(n_421), .Y(n_523) );
OAI222xp33_ASAP7_75t_L g524 ( .A1(n_439), .A2(n_442), .B1(n_455), .B2(n_459), .C1(n_460), .C2(n_463), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_442), .A2(n_378), .B1(n_404), .B2(n_343), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_464), .B(n_379), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_481), .A2(n_343), .B1(n_346), .B2(n_349), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_481), .A2(n_343), .B1(n_346), .B2(n_349), .Y(n_528) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_450), .A2(n_427), .B(n_403), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_459), .A2(n_420), .B1(n_381), .B2(n_367), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_436), .A2(n_343), .B1(n_312), .B2(n_331), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_486), .A2(n_343), .B1(n_352), .B2(n_342), .Y(n_532) );
AOI22xp33_ASAP7_75t_SL g533 ( .A1(n_444), .A2(n_367), .B1(n_379), .B2(n_390), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_500), .A2(n_312), .B1(n_390), .B2(n_331), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_475), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_450), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_462), .A2(n_343), .B1(n_312), .B2(n_331), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_457), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_471), .A2(n_343), .B1(n_342), .B2(n_388), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_454), .A2(n_352), .B1(n_342), .B2(n_388), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_473), .A2(n_390), .B1(n_356), .B2(n_427), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_505), .A2(n_356), .B1(n_353), .B2(n_333), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_437), .B(n_497), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_478), .A2(n_356), .B1(n_353), .B2(n_333), .Y(n_544) );
OAI221xp5_ASAP7_75t_L g545 ( .A1(n_489), .A2(n_286), .B1(n_281), .B2(n_279), .C(n_317), .Y(n_545) );
OAI22xp33_ASAP7_75t_L g546 ( .A1(n_435), .A2(n_338), .B1(n_352), .B2(n_390), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_490), .A2(n_353), .B1(n_305), .B2(n_318), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_464), .B(n_390), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_448), .A2(n_305), .B1(n_318), .B2(n_316), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_445), .A2(n_427), .B1(n_431), .B2(n_360), .Y(n_550) );
OAI222xp33_ASAP7_75t_L g551 ( .A1(n_453), .A2(n_431), .B1(n_377), .B2(n_279), .C1(n_340), .C2(n_360), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_457), .B(n_431), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_485), .A2(n_318), .B1(n_316), .B2(n_367), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_506), .A2(n_318), .B1(n_316), .B2(n_367), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_499), .A2(n_360), .B1(n_367), .B2(n_361), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_469), .A2(n_367), .B1(n_377), .B2(n_285), .Y(n_556) );
OAI221xp5_ASAP7_75t_SL g557 ( .A1(n_495), .A2(n_279), .B1(n_317), .B2(n_319), .C(n_328), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_470), .A2(n_360), .B1(n_367), .B2(n_361), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_472), .A2(n_377), .B1(n_285), .B2(n_340), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_467), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_465), .B(n_377), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_493), .A2(n_377), .B1(n_285), .B2(n_340), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_444), .B(n_377), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_494), .A2(n_361), .B1(n_340), .B2(n_317), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_507), .A2(n_285), .B1(n_340), .B2(n_302), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_456), .B(n_338), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_465), .B(n_19), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_468), .B(n_19), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_504), .A2(n_340), .B1(n_301), .B2(n_302), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_484), .A2(n_301), .B1(n_302), .B2(n_314), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_482), .A2(n_301), .B1(n_302), .B2(n_314), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g572 ( .A1(n_467), .A2(n_255), .B1(n_224), .B2(n_290), .C(n_280), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_498), .A2(n_338), .B1(n_280), .B2(n_290), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_482), .A2(n_334), .B1(n_336), .B2(n_328), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_468), .A2(n_290), .B1(n_280), .B2(n_168), .C(n_233), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_487), .A2(n_301), .B1(n_314), .B2(n_334), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_487), .A2(n_334), .B1(n_241), .B2(n_336), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_496), .A2(n_330), .B1(n_168), .B2(n_319), .Y(n_578) );
CKINVDCx14_ASAP7_75t_R g579 ( .A(n_449), .Y(n_579) );
OAI21xp5_ASAP7_75t_SL g580 ( .A1(n_477), .A2(n_354), .B(n_341), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_502), .A2(n_330), .B1(n_168), .B2(n_320), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_476), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_502), .A2(n_330), .B1(n_168), .B2(n_320), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_474), .A2(n_330), .B1(n_168), .B2(n_320), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_476), .B(n_168), .C(n_159), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_501), .A2(n_328), .B1(n_341), .B2(n_324), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_479), .Y(n_587) );
NAND3xp33_ASAP7_75t_L g588 ( .A(n_451), .B(n_168), .C(n_159), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_480), .A2(n_330), .B1(n_168), .B2(n_309), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_451), .A2(n_168), .B1(n_273), .B2(n_272), .C(n_264), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_456), .A2(n_492), .B1(n_479), .B2(n_488), .Y(n_591) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_492), .A2(n_354), .B1(n_341), .B2(n_335), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_456), .A2(n_330), .B1(n_168), .B2(n_309), .Y(n_593) );
AOI22xp33_ASAP7_75t_SL g594 ( .A1(n_456), .A2(n_354), .B1(n_341), .B2(n_335), .Y(n_594) );
OAI221xp5_ASAP7_75t_L g595 ( .A1(n_475), .A2(n_324), .B1(n_202), .B2(n_264), .C(n_272), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_483), .A2(n_303), .B1(n_326), .B2(n_309), .Y(n_596) );
OAI221xp5_ASAP7_75t_SL g597 ( .A1(n_491), .A2(n_229), .B1(n_253), .B2(n_273), .C(n_252), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_483), .B(n_160), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_488), .A2(n_303), .B1(n_326), .B2(n_354), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g600 ( .A1(n_439), .A2(n_354), .B1(n_335), .B2(n_252), .Y(n_600) );
AOI22xp33_ASAP7_75t_SL g601 ( .A1(n_439), .A2(n_354), .B1(n_335), .B2(n_155), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_458), .B(n_20), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_440), .A2(n_227), .B1(n_329), .B2(n_235), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_443), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_543), .B(n_160), .Y(n_605) );
OAI221xp5_ASAP7_75t_L g606 ( .A1(n_544), .A2(n_153), .B1(n_164), .B2(n_160), .C(n_163), .Y(n_606) );
NOR2xp33_ASAP7_75t_SL g607 ( .A(n_524), .B(n_335), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_582), .B(n_20), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_582), .B(n_21), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_587), .B(n_22), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_587), .B(n_22), .Y(n_611) );
OAI21xp33_ASAP7_75t_L g612 ( .A1(n_509), .A2(n_160), .B(n_163), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_519), .B(n_160), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_520), .B(n_335), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_515), .A2(n_250), .B1(n_237), .B2(n_235), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_519), .B(n_160), .Y(n_616) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_521), .Y(n_617) );
OAI221xp5_ASAP7_75t_L g618 ( .A1(n_522), .A2(n_153), .B1(n_163), .B2(n_160), .C(n_164), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_511), .B(n_23), .Y(n_619) );
NOR3xp33_ASAP7_75t_L g620 ( .A(n_588), .B(n_153), .C(n_237), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_521), .B(n_335), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g622 ( .A(n_588), .B(n_585), .C(n_600), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_511), .B(n_24), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_508), .A2(n_163), .B1(n_164), .B2(n_335), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g625 ( .A1(n_512), .A2(n_163), .B1(n_164), .B2(n_231), .C(n_230), .Y(n_625) );
OAI21xp5_ASAP7_75t_SL g626 ( .A1(n_579), .A2(n_164), .B(n_163), .Y(n_626) );
NOR2xp67_ASAP7_75t_L g627 ( .A(n_585), .B(n_25), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_513), .B(n_27), .Y(n_628) );
OAI21xp33_ASAP7_75t_L g629 ( .A1(n_530), .A2(n_163), .B(n_164), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_533), .B(n_335), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_527), .A2(n_163), .B1(n_164), .B2(n_155), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_513), .B(n_28), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_536), .B(n_28), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_536), .B(n_29), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_528), .A2(n_329), .B1(n_155), .B2(n_159), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_538), .B(n_164), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_538), .B(n_29), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_517), .A2(n_164), .B1(n_159), .B2(n_155), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_560), .B(n_30), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_560), .B(n_31), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_604), .B(n_31), .Y(n_641) );
OAI221xp5_ASAP7_75t_SL g642 ( .A1(n_532), .A2(n_231), .B1(n_329), .B2(n_34), .C(n_35), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_532), .A2(n_329), .B1(n_155), .B2(n_159), .Y(n_643) );
NAND4xp25_ASAP7_75t_L g644 ( .A(n_523), .B(n_32), .C(n_33), .D(n_34), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_604), .B(n_32), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_548), .B(n_33), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_546), .B(n_155), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_597), .A2(n_155), .B1(n_159), .B2(n_288), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_567), .B(n_155), .C(n_159), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_535), .B(n_529), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_535), .B(n_35), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_529), .B(n_36), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_510), .B(n_37), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_529), .B(n_552), .Y(n_654) );
NAND3xp33_ASAP7_75t_L g655 ( .A(n_568), .B(n_155), .C(n_159), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_541), .B(n_155), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_514), .B(n_37), .Y(n_657) );
OAI221xp5_ASAP7_75t_L g658 ( .A1(n_547), .A2(n_159), .B1(n_228), .B2(n_226), .C(n_225), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_531), .A2(n_159), .B1(n_310), .B2(n_304), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g660 ( .A(n_601), .B(n_306), .C(n_304), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_529), .B(n_38), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_592), .B(n_306), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_602), .B(n_39), .Y(n_663) );
OAI221xp5_ASAP7_75t_SL g664 ( .A1(n_540), .A2(n_40), .B1(n_228), .B2(n_226), .C(n_225), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_552), .B(n_40), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_561), .B(n_42), .Y(n_666) );
OAI221xp5_ASAP7_75t_SL g667 ( .A1(n_540), .A2(n_221), .B1(n_310), .B2(n_246), .C(n_240), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_526), .B(n_43), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_542), .A2(n_310), .B1(n_306), .B2(n_304), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_591), .B(n_306), .C(n_304), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g671 ( .A(n_590), .B(n_563), .C(n_572), .Y(n_671) );
NAND3xp33_ASAP7_75t_L g672 ( .A(n_562), .B(n_306), .C(n_304), .Y(n_672) );
NAND3xp33_ASAP7_75t_L g673 ( .A(n_580), .B(n_306), .C(n_304), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_534), .B(n_556), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_603), .B(n_44), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_603), .B(n_45), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_594), .B(n_306), .Y(n_677) );
OA21x2_ASAP7_75t_L g678 ( .A1(n_551), .A2(n_265), .B(n_221), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_525), .A2(n_310), .B1(n_306), .B2(n_304), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_598), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_516), .B(n_565), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_564), .B(n_47), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_550), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_559), .B(n_48), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_539), .B(n_553), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_586), .B(n_50), .Y(n_686) );
OA21x2_ASAP7_75t_L g687 ( .A1(n_580), .A2(n_259), .B(n_246), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_571), .B(n_576), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_570), .B(n_53), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_557), .A2(n_310), .B1(n_306), .B2(n_304), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_573), .B(n_54), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_573), .B(n_55), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_569), .A2(n_304), .B1(n_283), .B2(n_259), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_558), .B(n_56), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_566), .B(n_57), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_537), .B(n_59), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_596), .B(n_63), .Y(n_697) );
NOR3xp33_ASAP7_75t_L g698 ( .A(n_545), .B(n_240), .C(n_275), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_574), .B(n_64), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_518), .B(n_65), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_555), .B(n_304), .Y(n_701) );
OAI21xp5_ASAP7_75t_SL g702 ( .A1(n_593), .A2(n_283), .B(n_68), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_578), .B(n_66), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_683), .B(n_599), .Y(n_704) );
NAND3xp33_ASAP7_75t_SL g705 ( .A(n_607), .B(n_549), .C(n_554), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g706 ( .A(n_626), .B(n_577), .C(n_595), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_685), .A2(n_575), .B1(n_584), .B2(n_589), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_650), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_605), .B(n_583), .Y(n_709) );
NOR3xp33_ASAP7_75t_L g710 ( .A(n_644), .B(n_581), .C(n_70), .Y(n_710) );
AND2x4_ASAP7_75t_L g711 ( .A(n_617), .B(n_71), .Y(n_711) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_673), .B(n_283), .C(n_72), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_688), .A2(n_283), .B1(n_74), .B2(n_75), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_674), .A2(n_283), .B1(n_79), .B2(n_80), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_652), .B(n_73), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_681), .A2(n_283), .B1(n_275), .B2(n_85), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_663), .B(n_82), .Y(n_717) );
AND2x4_ASAP7_75t_L g718 ( .A(n_650), .B(n_84), .Y(n_718) );
NOR3xp33_ASAP7_75t_L g719 ( .A(n_618), .B(n_86), .C(n_88), .Y(n_719) );
NAND3xp33_ASAP7_75t_L g720 ( .A(n_622), .B(n_283), .C(n_91), .Y(n_720) );
NAND3xp33_ASAP7_75t_L g721 ( .A(n_652), .B(n_283), .C(n_94), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g722 ( .A(n_649), .B(n_99), .C(n_100), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_627), .A2(n_102), .B1(n_186), .B2(n_671), .Y(n_723) );
NOR3xp33_ASAP7_75t_L g724 ( .A(n_655), .B(n_653), .C(n_657), .Y(n_724) );
INVxp67_ASAP7_75t_L g725 ( .A(n_661), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_680), .B(n_661), .Y(n_726) );
AO21x2_ASAP7_75t_L g727 ( .A1(n_619), .A2(n_633), .B(n_634), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_613), .B(n_616), .Y(n_728) );
NAND4xp25_ASAP7_75t_L g729 ( .A(n_664), .B(n_642), .C(n_615), .D(n_667), .Y(n_729) );
OR2x2_ASAP7_75t_L g730 ( .A(n_665), .B(n_651), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_625), .A2(n_698), .B1(n_648), .B2(n_656), .Y(n_731) );
INVxp67_ASAP7_75t_L g732 ( .A(n_630), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_665), .B(n_640), .Y(n_733) );
AND2x4_ASAP7_75t_L g734 ( .A(n_614), .B(n_630), .Y(n_734) );
NOR3xp33_ASAP7_75t_L g735 ( .A(n_610), .B(n_611), .C(n_608), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_651), .B(n_687), .Y(n_736) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_701), .Y(n_737) );
NOR3xp33_ASAP7_75t_L g738 ( .A(n_609), .B(n_646), .C(n_632), .Y(n_738) );
AO21x2_ASAP7_75t_L g739 ( .A1(n_623), .A2(n_628), .B(n_645), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_640), .B(n_641), .Y(n_740) );
NOR3xp33_ASAP7_75t_SL g741 ( .A(n_702), .B(n_612), .C(n_656), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_687), .B(n_641), .Y(n_742) );
OA211x2_ASAP7_75t_L g743 ( .A1(n_677), .A2(n_662), .B(n_647), .C(n_621), .Y(n_743) );
OR2x2_ASAP7_75t_L g744 ( .A(n_636), .B(n_639), .Y(n_744) );
AOI221xp5_ASAP7_75t_L g745 ( .A1(n_637), .A2(n_643), .B1(n_690), .B2(n_658), .C(n_606), .Y(n_745) );
OA211x2_ASAP7_75t_L g746 ( .A1(n_677), .A2(n_662), .B(n_647), .C(n_621), .Y(n_746) );
NOR2x1_ASAP7_75t_L g747 ( .A(n_660), .B(n_670), .Y(n_747) );
OAI211xp5_ASAP7_75t_L g748 ( .A1(n_629), .A2(n_620), .B(n_701), .C(n_624), .Y(n_748) );
NAND3xp33_ASAP7_75t_L g749 ( .A(n_678), .B(n_672), .C(n_636), .Y(n_749) );
NAND3xp33_ASAP7_75t_L g750 ( .A(n_678), .B(n_692), .C(n_691), .Y(n_750) );
NAND4xp75_ASAP7_75t_L g751 ( .A(n_678), .B(n_695), .C(n_699), .D(n_666), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_666), .B(n_699), .Y(n_752) );
NAND4xp75_ASAP7_75t_L g753 ( .A(n_682), .B(n_686), .C(n_676), .D(n_675), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_696), .B(n_700), .Y(n_754) );
NAND3xp33_ASAP7_75t_L g755 ( .A(n_668), .B(n_684), .C(n_694), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_679), .B(n_669), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_693), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_703), .B(n_689), .Y(n_758) );
AND2x4_ASAP7_75t_L g759 ( .A(n_703), .B(n_697), .Y(n_759) );
NOR3xp33_ASAP7_75t_SL g760 ( .A(n_659), .B(n_635), .C(n_638), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_631), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_605), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_685), .A2(n_644), .B1(n_681), .B2(n_307), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_607), .B(n_524), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_654), .B(n_683), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_663), .B(n_579), .Y(n_766) );
AO22x1_ASAP7_75t_L g767 ( .A1(n_617), .A2(n_451), .B1(n_478), .B2(n_442), .Y(n_767) );
NOR3xp33_ASAP7_75t_L g768 ( .A(n_764), .B(n_706), .C(n_705), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_725), .B(n_765), .Y(n_769) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_708), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_710), .A2(n_763), .B1(n_764), .B2(n_729), .Y(n_771) );
BUFx2_ASAP7_75t_L g772 ( .A(n_767), .Y(n_772) );
NAND4xp75_ASAP7_75t_L g773 ( .A(n_743), .B(n_746), .C(n_747), .D(n_741), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_726), .B(n_725), .Y(n_774) );
OR2x2_ASAP7_75t_L g775 ( .A(n_730), .B(n_762), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_757), .B(n_728), .Y(n_776) );
XNOR2xp5_ASAP7_75t_L g777 ( .A(n_763), .B(n_733), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_742), .B(n_736), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_737), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_732), .B(n_737), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_727), .B(n_739), .Y(n_781) );
XNOR2xp5_ASAP7_75t_L g782 ( .A(n_751), .B(n_740), .Y(n_782) );
INVx2_ASAP7_75t_SL g783 ( .A(n_734), .Y(n_783) );
AND2x2_ASAP7_75t_SL g784 ( .A(n_734), .B(n_752), .Y(n_784) );
NOR4xp25_ASAP7_75t_L g785 ( .A(n_766), .B(n_705), .C(n_732), .D(n_750), .Y(n_785) );
NAND4xp75_ASAP7_75t_SL g786 ( .A(n_756), .B(n_754), .C(n_758), .D(n_717), .Y(n_786) );
NAND4xp75_ASAP7_75t_L g787 ( .A(n_741), .B(n_723), .C(n_745), .D(n_760), .Y(n_787) );
NOR4xp25_ASAP7_75t_L g788 ( .A(n_749), .B(n_704), .C(n_748), .D(n_731), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_744), .B(n_739), .Y(n_789) );
NAND4xp75_ASAP7_75t_L g790 ( .A(n_745), .B(n_760), .C(n_761), .D(n_715), .Y(n_790) );
NAND4xp75_ASAP7_75t_L g791 ( .A(n_709), .B(n_714), .C(n_713), .D(n_710), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_727), .Y(n_792) );
XNOR2xp5_ASAP7_75t_L g793 ( .A(n_753), .B(n_724), .Y(n_793) );
INVx4_ASAP7_75t_L g794 ( .A(n_711), .Y(n_794) );
AND2x2_ASAP7_75t_L g795 ( .A(n_718), .B(n_759), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_759), .B(n_738), .Y(n_796) );
BUFx2_ASAP7_75t_L g797 ( .A(n_711), .Y(n_797) );
XOR2x2_ASAP7_75t_L g798 ( .A(n_738), .B(n_724), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_721), .Y(n_799) );
INVxp67_ASAP7_75t_SL g800 ( .A(n_712), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_755), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_735), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_720), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_735), .B(n_707), .Y(n_804) );
NAND4xp75_ASAP7_75t_L g805 ( .A(n_722), .B(n_719), .C(n_707), .D(n_716), .Y(n_805) );
XNOR2xp5_ASAP7_75t_L g806 ( .A(n_790), .B(n_716), .Y(n_806) );
BUFx3_ASAP7_75t_L g807 ( .A(n_797), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_775), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_770), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_790), .A2(n_719), .B1(n_722), .B2(n_768), .Y(n_810) );
XOR2x2_ASAP7_75t_L g811 ( .A(n_798), .B(n_786), .Y(n_811) );
OR2x2_ASAP7_75t_L g812 ( .A(n_801), .B(n_779), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_775), .Y(n_813) );
OR2x2_ASAP7_75t_L g814 ( .A(n_801), .B(n_779), .Y(n_814) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_783), .Y(n_815) );
INVxp67_ASAP7_75t_L g816 ( .A(n_796), .Y(n_816) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_783), .Y(n_817) );
NOR2xp33_ASAP7_75t_SL g818 ( .A(n_794), .B(n_773), .Y(n_818) );
XNOR2x1_ASAP7_75t_SL g819 ( .A(n_793), .B(n_782), .Y(n_819) );
AND2x2_ASAP7_75t_L g820 ( .A(n_778), .B(n_789), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_784), .A2(n_794), .B1(n_772), .B2(n_797), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_778), .B(n_789), .Y(n_822) );
XOR2x2_ASAP7_75t_L g823 ( .A(n_798), .B(n_793), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_802), .B(n_780), .Y(n_824) );
INVx1_ASAP7_75t_SL g825 ( .A(n_772), .Y(n_825) );
XNOR2x1_ASAP7_75t_L g826 ( .A(n_771), .B(n_787), .Y(n_826) );
XOR2x2_ASAP7_75t_L g827 ( .A(n_777), .B(n_771), .Y(n_827) );
XNOR2xp5_ASAP7_75t_L g828 ( .A(n_777), .B(n_773), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_774), .Y(n_829) );
XNOR2xp5_ASAP7_75t_L g830 ( .A(n_787), .B(n_782), .Y(n_830) );
CKINVDCx8_ASAP7_75t_R g831 ( .A(n_804), .Y(n_831) );
AOI22xp5_ASAP7_75t_SL g832 ( .A1(n_828), .A2(n_794), .B1(n_802), .B2(n_780), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_826), .A2(n_799), .B1(n_781), .B2(n_792), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_809), .Y(n_834) );
INVx3_ASAP7_75t_L g835 ( .A(n_807), .Y(n_835) );
INVx2_ASAP7_75t_SL g836 ( .A(n_815), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_809), .Y(n_837) );
INVxp67_ASAP7_75t_SL g838 ( .A(n_826), .Y(n_838) );
INVx1_ASAP7_75t_SL g839 ( .A(n_825), .Y(n_839) );
OAI22x1_ASAP7_75t_L g840 ( .A1(n_830), .A2(n_792), .B1(n_785), .B2(n_788), .Y(n_840) );
XNOR2x1_ASAP7_75t_L g841 ( .A(n_819), .B(n_805), .Y(n_841) );
AOI22xp5_ASAP7_75t_L g842 ( .A1(n_830), .A2(n_805), .B1(n_791), .B2(n_784), .Y(n_842) );
HB1xp67_ASAP7_75t_L g843 ( .A(n_812), .Y(n_843) );
OA22x2_ASAP7_75t_L g844 ( .A1(n_828), .A2(n_799), .B1(n_776), .B2(n_795), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_827), .A2(n_791), .B1(n_784), .B2(n_795), .Y(n_845) );
INVxp67_ASAP7_75t_L g846 ( .A(n_818), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_843), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_843), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_839), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_835), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_835), .Y(n_851) );
OAI322xp33_ASAP7_75t_L g852 ( .A1(n_838), .A2(n_816), .A3(n_810), .B1(n_824), .B2(n_819), .C1(n_821), .C2(n_806), .Y(n_852) );
OAI322xp33_ASAP7_75t_L g853 ( .A1(n_838), .A2(n_806), .A3(n_812), .B1(n_814), .B2(n_827), .C1(n_823), .C2(n_817), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_836), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_849), .Y(n_855) );
OAI322xp33_ASAP7_75t_L g856 ( .A1(n_854), .A2(n_841), .A3(n_832), .B1(n_842), .B2(n_844), .C1(n_845), .C2(n_846), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_848), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_848), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_852), .A2(n_823), .B1(n_844), .B2(n_840), .Y(n_859) );
OAI22xp33_ASAP7_75t_L g860 ( .A1(n_855), .A2(n_850), .B1(n_851), .B2(n_831), .Y(n_860) );
INVx1_ASAP7_75t_SL g861 ( .A(n_857), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_858), .Y(n_862) );
NAND4xp25_ASAP7_75t_SL g863 ( .A(n_861), .B(n_859), .C(n_856), .D(n_833), .Y(n_863) );
NOR2x1_ASAP7_75t_L g864 ( .A(n_860), .B(n_853), .Y(n_864) );
NOR2x1_ASAP7_75t_L g865 ( .A(n_862), .B(n_850), .Y(n_865) );
INVxp67_ASAP7_75t_L g866 ( .A(n_865), .Y(n_866) );
NOR2xp67_ASAP7_75t_L g867 ( .A(n_863), .B(n_847), .Y(n_867) );
AND4x1_ASAP7_75t_L g868 ( .A(n_867), .B(n_864), .C(n_859), .D(n_833), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_866), .A2(n_831), .B1(n_814), .B2(n_837), .Y(n_869) );
INVx4_ASAP7_75t_L g870 ( .A(n_868), .Y(n_870) );
INVxp67_ASAP7_75t_SL g871 ( .A(n_869), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_871), .A2(n_811), .B1(n_807), .B2(n_834), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_872), .Y(n_873) );
AOI221xp5_ASAP7_75t_L g874 ( .A1(n_873), .A2(n_870), .B1(n_837), .B2(n_834), .C(n_811), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_874), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_875), .A2(n_829), .B1(n_808), .B2(n_813), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_876), .Y(n_877) );
AOI221xp5_ASAP7_75t_L g878 ( .A1(n_877), .A2(n_820), .B1(n_822), .B2(n_800), .C(n_803), .Y(n_878) );
AOI211xp5_ASAP7_75t_L g879 ( .A1(n_878), .A2(n_822), .B(n_820), .C(n_769), .Y(n_879) );
endmodule