module real_aes_17502_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1583;
wire n_360;
wire n_1284;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1605;
wire n_1056;
wire n_1592;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1343;
wire n_465;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1596;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1595;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_1584;
wire n_1277;
wire n_559;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1352;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g775 ( .A(n_0), .Y(n_775) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1), .Y(n_1083) );
AOI221x1_ASAP7_75t_SL g786 ( .A1(n_2), .A2(n_264), .B1(n_787), .B2(n_788), .C(n_789), .Y(n_786) );
AOI21xp33_ASAP7_75t_L g854 ( .A1(n_2), .A2(n_480), .B(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g716 ( .A(n_3), .Y(n_716) );
OAI211xp5_ASAP7_75t_L g753 ( .A1(n_3), .A2(n_754), .B(n_755), .C(n_762), .Y(n_753) );
CKINVDCx5p33_ASAP7_75t_R g983 ( .A(n_4), .Y(n_983) );
INVx1_ASAP7_75t_L g581 ( .A(n_5), .Y(n_581) );
INVx1_ASAP7_75t_L g676 ( .A(n_6), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_6), .A2(n_120), .B1(n_706), .B2(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g343 ( .A(n_7), .Y(n_343) );
OAI22xp33_ASAP7_75t_L g470 ( .A1(n_7), .A2(n_132), .B1(n_471), .B2(n_477), .Y(n_470) );
AOI22xp33_ASAP7_75t_SL g1078 ( .A1(n_8), .A2(n_252), .B1(n_706), .B2(n_951), .Y(n_1078) );
AOI221xp5_ASAP7_75t_L g1095 ( .A1(n_8), .A2(n_135), .B1(n_321), .B2(n_330), .C(n_1096), .Y(n_1095) );
INVxp67_ASAP7_75t_SL g1147 ( .A(n_9), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_9), .A2(n_28), .B1(n_314), .B2(n_660), .Y(n_1155) );
INVx1_ASAP7_75t_L g1173 ( .A(n_10), .Y(n_1173) );
AOI221xp5_ASAP7_75t_L g1240 ( .A1(n_11), .A2(n_118), .B1(n_330), .B2(n_655), .C(n_657), .Y(n_1240) );
INVx1_ASAP7_75t_L g1262 ( .A(n_11), .Y(n_1262) );
INVx1_ASAP7_75t_L g292 ( .A(n_12), .Y(n_292) );
AND2x2_ASAP7_75t_L g317 ( .A(n_12), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g341 ( .A(n_12), .B(n_242), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_12), .B(n_302), .Y(n_558) );
AOI22xp5_ASAP7_75t_SL g1313 ( .A1(n_13), .A2(n_266), .B1(n_1296), .B2(n_1304), .Y(n_1313) );
OAI221xp5_ASAP7_75t_L g350 ( .A1(n_14), .A2(n_265), .B1(n_351), .B2(n_355), .C(n_361), .Y(n_350) );
INVx1_ASAP7_75t_L g460 ( .A(n_14), .Y(n_460) );
OAI211xp5_ASAP7_75t_L g505 ( .A1(n_15), .A2(n_506), .B(n_510), .C(n_517), .Y(n_505) );
INVx1_ASAP7_75t_L g538 ( .A(n_15), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_16), .A2(n_197), .B1(n_442), .B2(n_871), .Y(n_979) );
AOI221xp5_ASAP7_75t_L g1003 ( .A1(n_16), .A2(n_99), .B1(n_682), .B2(n_761), .C(n_1004), .Y(n_1003) );
INVx1_ASAP7_75t_L g1186 ( .A(n_17), .Y(n_1186) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_18), .A2(n_279), .B1(n_1085), .B2(n_1086), .Y(n_1084) );
OAI211xp5_ASAP7_75t_L g1088 ( .A1(n_18), .A2(n_1089), .B(n_1090), .C(n_1094), .Y(n_1088) );
INVx1_ASAP7_75t_L g973 ( .A(n_19), .Y(n_973) );
INVx2_ASAP7_75t_L g1291 ( .A(n_20), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_20), .B(n_1292), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_20), .B(n_111), .Y(n_1299) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_21), .A2(n_172), .B1(n_492), .B2(n_496), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_21), .A2(n_172), .B1(n_543), .B2(n_545), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_22), .A2(n_149), .B1(n_403), .B2(n_811), .Y(n_810) );
OAI221xp5_ASAP7_75t_L g818 ( .A1(n_22), .A2(n_244), .B1(n_819), .B2(n_821), .C(n_823), .Y(n_818) );
AOI22xp5_ASAP7_75t_SL g1327 ( .A1(n_23), .A2(n_148), .B1(n_1296), .B2(n_1304), .Y(n_1327) );
AOI22xp5_ASAP7_75t_SL g1322 ( .A1(n_24), .A2(n_259), .B1(n_1293), .B2(n_1298), .Y(n_1322) );
OAI22xp33_ASAP7_75t_L g502 ( .A1(n_25), .A2(n_41), .B1(n_294), .B2(n_503), .Y(n_502) );
OAI22xp33_ASAP7_75t_L g521 ( .A1(n_25), .A2(n_41), .B1(n_522), .B2(n_525), .Y(n_521) );
INVx1_ASAP7_75t_L g1080 ( .A(n_26), .Y(n_1080) );
OAI221xp5_ASAP7_75t_L g1100 ( .A1(n_26), .A2(n_170), .B1(n_1101), .B2(n_1102), .C(n_1103), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_27), .A2(n_213), .B1(n_438), .B2(n_442), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_27), .A2(n_134), .B1(n_1055), .B2(n_1067), .Y(n_1066) );
INVxp67_ASAP7_75t_SL g1136 ( .A(n_28), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_29), .A2(n_222), .B1(n_433), .B2(n_736), .Y(n_971) );
AOI221xp5_ASAP7_75t_L g988 ( .A1(n_29), .A2(n_64), .B1(n_935), .B2(n_989), .C(n_991), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_30), .A2(n_134), .B1(n_438), .B2(n_442), .Y(n_1044) );
AOI22xp33_ASAP7_75t_SL g1058 ( .A1(n_30), .A2(n_213), .B1(n_1059), .B2(n_1060), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_31), .A2(n_79), .B1(n_660), .B2(n_661), .Y(n_1241) );
INVx1_ASAP7_75t_L g1266 ( .A(n_31), .Y(n_1266) );
INVx1_ASAP7_75t_L g1122 ( .A(n_32), .Y(n_1122) );
INVx1_ASAP7_75t_L g624 ( .A(n_33), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g1576 ( .A1(n_34), .A2(n_127), .B1(n_503), .B2(n_1577), .Y(n_1576) );
OAI22xp5_ASAP7_75t_L g1579 ( .A1(n_34), .A2(n_280), .B1(n_1580), .B2(n_1581), .Y(n_1579) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_35), .A2(n_109), .B1(n_438), .B2(n_704), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_35), .A2(n_253), .B1(n_935), .B2(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g912 ( .A(n_36), .Y(n_912) );
INVx1_ASAP7_75t_L g1575 ( .A(n_37), .Y(n_1575) );
INVx1_ASAP7_75t_L g577 ( .A(n_38), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_39), .A2(n_245), .B1(n_744), .B2(n_746), .Y(n_743) );
INVx1_ASAP7_75t_L g756 ( .A(n_39), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g1287 ( .A1(n_40), .A2(n_195), .B1(n_1288), .B2(n_1293), .Y(n_1287) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_42), .A2(n_239), .B1(n_682), .B2(n_1153), .Y(n_1245) );
AOI22xp33_ASAP7_75t_L g1267 ( .A1(n_42), .A2(n_118), .B1(n_698), .B2(n_946), .Y(n_1267) );
CKINVDCx5p33_ASAP7_75t_R g879 ( .A(n_43), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_44), .A2(n_82), .B1(n_701), .B2(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g902 ( .A(n_44), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g1342 ( .A1(n_45), .A2(n_105), .B1(n_1296), .B2(n_1343), .Y(n_1342) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_46), .A2(n_145), .B1(n_321), .B2(n_324), .C(n_330), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_46), .A2(n_86), .B1(n_433), .B2(n_457), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g734 ( .A1(n_47), .A2(n_125), .B1(n_735), .B2(n_736), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_47), .A2(n_245), .B1(n_314), .B2(n_761), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g1295 ( .A1(n_48), .A2(n_199), .B1(n_1296), .B2(n_1298), .Y(n_1295) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_49), .A2(n_183), .B1(n_333), .B2(n_338), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_49), .A2(n_110), .B1(n_447), .B2(n_450), .Y(n_446) );
INVx1_ASAP7_75t_L g1139 ( .A(n_50), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_50), .A2(n_142), .B1(n_1099), .B2(n_1153), .Y(n_1152) );
AOI22xp5_ASAP7_75t_L g1305 ( .A1(n_51), .A2(n_92), .B1(n_1288), .B2(n_1296), .Y(n_1305) );
INVx1_ASAP7_75t_L g573 ( .A(n_52), .Y(n_573) );
INVx1_ASAP7_75t_L g389 ( .A(n_53), .Y(n_389) );
INVx1_ASAP7_75t_L g419 ( .A(n_53), .Y(n_419) );
INVx1_ASAP7_75t_L g742 ( .A(n_54), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_54), .A2(n_254), .B1(n_314), .B2(n_761), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_55), .A2(n_622), .B1(n_709), .B2(n_710), .Y(n_621) );
INVxp67_ASAP7_75t_L g710 ( .A(n_55), .Y(n_710) );
INVx1_ASAP7_75t_L g1216 ( .A(n_56), .Y(n_1216) );
AOI22xp5_ASAP7_75t_L g1307 ( .A1(n_57), .A2(n_273), .B1(n_1288), .B2(n_1293), .Y(n_1307) );
CKINVDCx5p33_ASAP7_75t_R g793 ( .A(n_58), .Y(n_793) );
CKINVDCx5p33_ASAP7_75t_R g648 ( .A(n_59), .Y(n_648) );
INVx1_ASAP7_75t_L g1574 ( .A(n_60), .Y(n_1574) );
INVx1_ASAP7_75t_L g1250 ( .A(n_61), .Y(n_1250) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_62), .A2(n_712), .B1(n_713), .B2(n_769), .Y(n_711) );
INVxp67_ASAP7_75t_L g769 ( .A(n_62), .Y(n_769) );
INVx1_ASAP7_75t_L g286 ( .A(n_63), .Y(n_286) );
AOI22xp33_ASAP7_75t_SL g980 ( .A1(n_64), .A2(n_204), .B1(n_434), .B2(n_868), .Y(n_980) );
INVx2_ASAP7_75t_L g395 ( .A(n_65), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g1590 ( .A1(n_66), .A2(n_228), .B1(n_1055), .B2(n_1063), .Y(n_1590) );
AOI22xp33_ASAP7_75t_L g1602 ( .A1(n_66), .A2(n_101), .B1(n_1603), .B2(n_1605), .Y(n_1602) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_67), .A2(n_164), .B1(n_503), .B2(n_1125), .Y(n_1124) );
OAI22xp5_ASAP7_75t_L g1160 ( .A1(n_67), .A2(n_164), .B1(n_1161), .B2(n_1163), .Y(n_1160) );
INVx1_ASAP7_75t_L g1121 ( .A(n_68), .Y(n_1121) );
AOI22xp5_ASAP7_75t_L g1323 ( .A1(n_69), .A2(n_73), .B1(n_1288), .B2(n_1296), .Y(n_1323) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_70), .A2(n_235), .B1(n_402), .B2(n_413), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_71), .A2(n_276), .B1(n_681), .B2(n_682), .Y(n_680) );
INVx1_ASAP7_75t_L g696 ( .A(n_71), .Y(n_696) );
INVx1_ASAP7_75t_L g589 ( .A(n_72), .Y(n_589) );
OAI22xp33_ASAP7_75t_SL g1531 ( .A1(n_74), .A2(n_277), .B1(n_524), .B2(n_1532), .Y(n_1531) );
OAI22xp33_ASAP7_75t_L g1542 ( .A1(n_74), .A2(n_277), .B1(n_1543), .B2(n_1544), .Y(n_1542) );
INVx1_ASAP7_75t_L g400 ( .A(n_75), .Y(n_400) );
OAI22xp33_ASAP7_75t_L g1540 ( .A1(n_76), .A2(n_268), .B1(n_544), .B2(n_546), .Y(n_1540) );
OAI22xp5_ASAP7_75t_L g1553 ( .A1(n_76), .A2(n_268), .B1(n_1554), .B2(n_1555), .Y(n_1553) );
INVx1_ASAP7_75t_L g1171 ( .A(n_77), .Y(n_1171) );
AOI221xp5_ASAP7_75t_L g1244 ( .A1(n_78), .A2(n_113), .B1(n_657), .B2(n_930), .C(n_1097), .Y(n_1244) );
INVxp67_ASAP7_75t_SL g1254 ( .A(n_78), .Y(n_1254) );
INVxp67_ASAP7_75t_SL g1256 ( .A(n_79), .Y(n_1256) );
INVx1_ASAP7_75t_L g1509 ( .A(n_80), .Y(n_1509) );
INVxp67_ASAP7_75t_SL g717 ( .A(n_81), .Y(n_717) );
OAI221xp5_ASAP7_75t_L g766 ( .A1(n_81), .A2(n_231), .B1(n_356), .B2(n_399), .C(n_767), .Y(n_766) );
AOI221xp5_ASAP7_75t_L g881 ( .A1(n_82), .A2(n_133), .B1(n_682), .B2(n_882), .C(n_884), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_83), .A2(n_120), .B1(n_660), .B2(n_661), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_83), .A2(n_212), .B1(n_698), .B2(n_701), .Y(n_697) );
INVx1_ASAP7_75t_L g516 ( .A(n_84), .Y(n_516) );
OAI211xp5_ASAP7_75t_L g528 ( .A1(n_84), .A2(n_529), .B(n_531), .C(n_533), .Y(n_528) );
INVx1_ASAP7_75t_L g1175 ( .A(n_85), .Y(n_1175) );
INVxp67_ASAP7_75t_SL g369 ( .A(n_86), .Y(n_369) );
INVx1_ASAP7_75t_L g977 ( .A(n_87), .Y(n_977) );
XOR2x2_ASAP7_75t_L g485 ( .A(n_88), .B(n_486), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g921 ( .A1(n_89), .A2(n_188), .B1(n_563), .B2(n_791), .Y(n_921) );
NOR2xp33_ASAP7_75t_L g964 ( .A(n_89), .B(n_543), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g1210 ( .A1(n_90), .A2(n_96), .B1(n_522), .B2(n_1211), .Y(n_1210) );
OAI22xp33_ASAP7_75t_L g1221 ( .A1(n_90), .A2(n_123), .B1(n_294), .B2(n_1222), .Y(n_1221) );
AOI22xp5_ASAP7_75t_L g1303 ( .A1(n_91), .A2(n_209), .B1(n_1293), .B2(n_1304), .Y(n_1303) );
INVx1_ASAP7_75t_L g1506 ( .A(n_93), .Y(n_1506) );
CKINVDCx5p33_ASAP7_75t_R g878 ( .A(n_94), .Y(n_878) );
OAI221xp5_ASAP7_75t_SL g642 ( .A1(n_95), .A2(n_97), .B1(n_643), .B2(n_645), .C(n_647), .Y(n_642) );
INVx1_ASAP7_75t_L g669 ( .A(n_95), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g1223 ( .A1(n_96), .A2(n_193), .B1(n_492), .B2(n_1224), .Y(n_1223) );
INVx1_ASAP7_75t_L g685 ( .A(n_97), .Y(n_685) );
CKINVDCx5p33_ASAP7_75t_R g723 ( .A(n_98), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_99), .A2(n_136), .B1(n_447), .B2(n_450), .Y(n_970) );
INVx1_ASAP7_75t_L g1024 ( .A(n_100), .Y(n_1024) );
AOI22xp33_ASAP7_75t_SL g1596 ( .A1(n_101), .A2(n_221), .B1(n_1055), .B2(n_1067), .Y(n_1596) );
OA222x2_ASAP7_75t_L g777 ( .A1(n_102), .A2(n_223), .B1(n_244), .B2(n_778), .C1(n_780), .C2(n_784), .Y(n_777) );
INVx1_ASAP7_75t_L g835 ( .A(n_102), .Y(n_835) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_103), .Y(n_288) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_103), .B(n_286), .Y(n_1289) );
INVx1_ASAP7_75t_L g1027 ( .A(n_104), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g1033 ( .A1(n_104), .A2(n_262), .B1(n_1034), .B2(n_1035), .Y(n_1033) );
INVx1_ASAP7_75t_L g1276 ( .A(n_105), .Y(n_1276) );
INVx1_ASAP7_75t_L g1187 ( .A(n_106), .Y(n_1187) );
CKINVDCx5p33_ASAP7_75t_R g875 ( .A(n_107), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g1345 ( .A1(n_108), .A2(n_171), .B1(n_1288), .B2(n_1293), .Y(n_1345) );
INVxp67_ASAP7_75t_SL g1104 ( .A(n_109), .Y(n_1104) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_110), .A2(n_168), .B1(n_326), .B2(n_371), .C(n_373), .Y(n_370) );
INVx1_ASAP7_75t_L g1292 ( .A(n_111), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_111), .B(n_1291), .Y(n_1297) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_112), .A2(n_210), .B1(n_314), .B2(n_761), .Y(n_926) );
INVxp67_ASAP7_75t_SL g944 ( .A(n_112), .Y(n_944) );
INVx1_ASAP7_75t_L g1264 ( .A(n_113), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_114), .A2(n_122), .B1(n_438), .B2(n_836), .Y(n_869) );
INVx1_ASAP7_75t_L g905 ( .A(n_114), .Y(n_905) );
AOI22xp5_ASAP7_75t_L g1314 ( .A1(n_115), .A2(n_208), .B1(n_1288), .B2(n_1293), .Y(n_1314) );
AOI22xp33_ASAP7_75t_SL g1587 ( .A1(n_116), .A2(n_143), .B1(n_1588), .B2(n_1589), .Y(n_1587) );
AOI22xp33_ASAP7_75t_L g1598 ( .A1(n_116), .A2(n_180), .B1(n_1049), .B2(n_1599), .Y(n_1598) );
INVx1_ASAP7_75t_L g1028 ( .A(n_117), .Y(n_1028) );
INVx1_ASAP7_75t_L g864 ( .A(n_119), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_119), .A2(n_249), .B1(n_364), .B2(n_367), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_121), .A2(n_253), .B1(n_438), .B2(n_1076), .Y(n_1075) );
AOI21xp33_ASAP7_75t_L g1106 ( .A1(n_121), .A2(n_373), .B(n_759), .Y(n_1106) );
INVx1_ASAP7_75t_L g887 ( .A(n_122), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g1218 ( .A1(n_123), .A2(n_193), .B1(n_545), .B2(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g633 ( .A(n_124), .Y(n_633) );
AOI21xp33_ASAP7_75t_L g758 ( .A1(n_125), .A2(n_679), .B(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_126), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g423 ( .A(n_126), .Y(n_423) );
INVx1_ASAP7_75t_L g455 ( .A(n_126), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g1584 ( .A1(n_127), .A2(n_275), .B1(n_522), .B2(n_1038), .Y(n_1584) );
INVx1_ASAP7_75t_L g1517 ( .A(n_128), .Y(n_1517) );
INVx1_ASAP7_75t_L g1021 ( .A(n_129), .Y(n_1021) );
AOI22xp33_ASAP7_75t_SL g1042 ( .A1(n_130), .A2(n_158), .B1(n_434), .B2(n_1043), .Y(n_1042) );
AOI22xp33_ASAP7_75t_SL g1062 ( .A1(n_130), .A2(n_233), .B1(n_1059), .B2(n_1063), .Y(n_1062) );
OAI22xp33_ASAP7_75t_L g1071 ( .A1(n_131), .A2(n_220), .B1(n_477), .B2(n_632), .Y(n_1071) );
INVx1_ASAP7_75t_L g1092 ( .A(n_131), .Y(n_1092) );
INVx1_ASAP7_75t_L g346 ( .A(n_132), .Y(n_346) );
AOI22xp33_ASAP7_75t_SL g873 ( .A1(n_133), .A2(n_173), .B1(n_457), .B2(n_868), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_135), .A2(n_205), .B1(n_434), .B2(n_744), .Y(n_1074) );
INVx1_ASAP7_75t_L g993 ( .A(n_136), .Y(n_993) );
INVx1_ASAP7_75t_L g1123 ( .A(n_137), .Y(n_1123) );
INVxp67_ASAP7_75t_SL g976 ( .A(n_138), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_138), .A2(n_250), .B1(n_364), .B2(n_997), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_139), .A2(n_263), .B1(n_333), .B2(n_338), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_139), .A2(n_247), .B1(n_444), .B2(n_706), .Y(n_856) );
NOR2xp33_ASAP7_75t_L g1247 ( .A(n_140), .B(n_356), .Y(n_1247) );
INVxp67_ASAP7_75t_SL g1272 ( .A(n_140), .Y(n_1272) );
XNOR2xp5_ASAP7_75t_L g1068 ( .A(n_141), .B(n_1069), .Y(n_1068) );
INVxp67_ASAP7_75t_SL g1130 ( .A(n_142), .Y(n_1130) );
AOI22xp33_ASAP7_75t_SL g1606 ( .A1(n_143), .A2(n_241), .B1(n_735), .B2(n_946), .Y(n_1606) );
INVx1_ASAP7_75t_L g727 ( .A(n_144), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_144), .A2(n_184), .B1(n_751), .B2(n_752), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_145), .A2(n_190), .B1(n_431), .B2(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g1514 ( .A(n_146), .Y(n_1514) );
INVx1_ASAP7_75t_L g934 ( .A(n_147), .Y(n_934) );
INVx1_ASAP7_75t_L g837 ( .A(n_149), .Y(n_837) );
INVx1_ASAP7_75t_L g1341 ( .A(n_150), .Y(n_1341) );
CKINVDCx5p33_ASAP7_75t_R g741 ( .A(n_151), .Y(n_741) );
CKINVDCx5p33_ASAP7_75t_R g802 ( .A(n_152), .Y(n_802) );
INVx1_ASAP7_75t_L g588 ( .A(n_153), .Y(n_588) );
INVx1_ASAP7_75t_L g984 ( .A(n_154), .Y(n_984) );
INVx1_ASAP7_75t_L g731 ( .A(n_155), .Y(n_731) );
AOI21xp33_ASAP7_75t_L g763 ( .A1(n_155), .A2(n_326), .B(n_373), .Y(n_763) );
INVx1_ASAP7_75t_L g1180 ( .A(n_156), .Y(n_1180) );
INVx1_ASAP7_75t_L g1246 ( .A(n_157), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_158), .A2(n_272), .B1(n_1055), .B2(n_1056), .Y(n_1054) );
INVx1_ASAP7_75t_L g1249 ( .A(n_159), .Y(n_1249) );
OAI322xp33_ASAP7_75t_L g1252 ( .A1(n_159), .A2(n_615), .A3(n_635), .B1(n_737), .B2(n_1253), .C1(n_1257), .C2(n_1263), .Y(n_1252) );
INVx1_ASAP7_75t_L g1539 ( .A(n_160), .Y(n_1539) );
OAI211xp5_ASAP7_75t_L g1545 ( .A1(n_160), .A2(n_939), .B(n_1546), .C(n_1548), .Y(n_1545) );
AOI22xp5_ASAP7_75t_L g1346 ( .A1(n_161), .A2(n_206), .B1(n_1296), .B2(n_1343), .Y(n_1346) );
BUFx3_ASAP7_75t_L g388 ( .A(n_162), .Y(n_388) );
AOI22xp33_ASAP7_75t_SL g931 ( .A1(n_163), .A2(n_278), .B1(n_761), .B2(n_932), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_163), .A2(n_211), .B1(n_825), .B2(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g1237 ( .A(n_165), .Y(n_1237) );
INVx1_ASAP7_75t_L g1507 ( .A(n_166), .Y(n_1507) );
INVx1_ASAP7_75t_L g1510 ( .A(n_167), .Y(n_1510) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_168), .A2(n_183), .B1(n_438), .B2(n_442), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g1537 ( .A(n_169), .Y(n_1537) );
INVx1_ASAP7_75t_L g1081 ( .A(n_170), .Y(n_1081) );
XNOR2x1_ASAP7_75t_L g1501 ( .A(n_171), .B(n_1502), .Y(n_1501) );
AOI22xp33_ASAP7_75t_L g1561 ( .A1(n_171), .A2(n_1562), .B1(n_1607), .B2(n_1609), .Y(n_1561) );
AOI211xp5_ASAP7_75t_SL g899 ( .A1(n_173), .A2(n_900), .B(n_901), .C(n_904), .Y(n_899) );
CKINVDCx5p33_ASAP7_75t_R g975 ( .A(n_174), .Y(n_975) );
INVx1_ASAP7_75t_L g1007 ( .A(n_175), .Y(n_1007) );
AOI22xp5_ASAP7_75t_L g1308 ( .A1(n_175), .A2(n_236), .B1(n_1296), .B2(n_1304), .Y(n_1308) );
INVx1_ASAP7_75t_L g1131 ( .A(n_176), .Y(n_1131) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_177), .Y(n_299) );
INVx1_ASAP7_75t_L g627 ( .A(n_178), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_179), .A2(n_214), .B1(n_450), .B2(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g886 ( .A(n_179), .Y(n_886) );
AOI22xp33_ASAP7_75t_SL g1594 ( .A1(n_180), .A2(n_241), .B1(n_1060), .B2(n_1595), .Y(n_1594) );
OAI221xp5_ASAP7_75t_L g936 ( .A1(n_181), .A2(n_215), .B1(n_937), .B2(n_938), .C(n_939), .Y(n_936) );
INVx1_ASAP7_75t_L g956 ( .A(n_181), .Y(n_956) );
OAI22xp33_ASAP7_75t_SL g922 ( .A1(n_182), .A2(n_229), .B1(n_801), .B2(n_903), .Y(n_922) );
INVx1_ASAP7_75t_L g959 ( .A(n_182), .Y(n_959) );
INVx1_ASAP7_75t_L g726 ( .A(n_184), .Y(n_726) );
INVx1_ASAP7_75t_L g924 ( .A(n_185), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_185), .A2(n_278), .B1(n_825), .B2(n_951), .Y(n_950) );
AOI21xp5_ASAP7_75t_SL g929 ( .A1(n_186), .A2(n_678), .B(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g943 ( .A(n_186), .Y(n_943) );
CKINVDCx5p33_ASAP7_75t_R g928 ( .A(n_187), .Y(n_928) );
INVx1_ASAP7_75t_L g958 ( .A(n_188), .Y(n_958) );
INVx1_ASAP7_75t_L g1573 ( .A(n_189), .Y(n_1573) );
OAI211xp5_ASAP7_75t_L g1582 ( .A1(n_189), .A2(n_531), .B(n_1213), .C(n_1583), .Y(n_1582) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_190), .Y(n_365) );
OAI211xp5_ASAP7_75t_L g1212 ( .A1(n_191), .A2(n_1213), .B(n_1214), .C(n_1215), .Y(n_1212) );
INVx1_ASAP7_75t_L g1228 ( .A(n_191), .Y(n_1228) );
INVx1_ASAP7_75t_L g1145 ( .A(n_192), .Y(n_1145) );
INVx1_ASAP7_75t_L g560 ( .A(n_194), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g1269 ( .A(n_196), .Y(n_1269) );
INVx1_ASAP7_75t_L g992 ( .A(n_197), .Y(n_992) );
INVx1_ASAP7_75t_L g1116 ( .A(n_198), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_200), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g861 ( .A(n_201), .Y(n_861) );
XOR2x2_ASAP7_75t_L g308 ( .A(n_202), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g513 ( .A(n_203), .Y(n_513) );
INVx1_ASAP7_75t_L g1005 ( .A(n_204), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_205), .A2(n_252), .B1(n_682), .B2(n_935), .Y(n_1107) );
INVx1_ASAP7_75t_L g1242 ( .A(n_207), .Y(n_1242) );
INVxp67_ASAP7_75t_L g949 ( .A(n_210), .Y(n_949) );
AOI21xp33_ASAP7_75t_L g925 ( .A1(n_211), .A2(n_678), .B(n_679), .Y(n_925) );
AOI21xp33_ASAP7_75t_L g677 ( .A1(n_212), .A2(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_L g908 ( .A(n_214), .Y(n_908) );
INVxp67_ASAP7_75t_SL g961 ( .A(n_215), .Y(n_961) );
INVx1_ASAP7_75t_L g1140 ( .A(n_216), .Y(n_1140) );
INVx1_ASAP7_75t_L g564 ( .A(n_217), .Y(n_564) );
INVx1_ASAP7_75t_L g1177 ( .A(n_218), .Y(n_1177) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_219), .Y(n_298) );
INVx1_ASAP7_75t_L g1091 ( .A(n_220), .Y(n_1091) );
AOI22xp33_ASAP7_75t_SL g1600 ( .A1(n_221), .A2(n_228), .B1(n_442), .B2(n_735), .Y(n_1600) );
INVx1_ASAP7_75t_L g1006 ( .A(n_222), .Y(n_1006) );
INVx1_ASAP7_75t_L g824 ( .A(n_223), .Y(n_824) );
INVx1_ASAP7_75t_L g722 ( .A(n_224), .Y(n_722) );
INVx1_ASAP7_75t_L g1134 ( .A(n_225), .Y(n_1134) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_226), .Y(n_815) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_227), .A2(n_237), .B1(n_655), .B2(n_657), .C(n_658), .Y(n_654) );
INVx1_ASAP7_75t_L g692 ( .A(n_227), .Y(n_692) );
INVx1_ASAP7_75t_L g963 ( .A(n_229), .Y(n_963) );
XNOR2xp5_ASAP7_75t_L g1014 ( .A(n_230), .B(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g720 ( .A(n_231), .Y(n_720) );
INVx1_ASAP7_75t_L g1183 ( .A(n_232), .Y(n_1183) );
AOI22xp33_ASAP7_75t_SL g1048 ( .A1(n_233), .A2(n_272), .B1(n_868), .B2(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g1513 ( .A(n_234), .Y(n_1513) );
OAI211xp5_ASAP7_75t_L g311 ( .A1(n_235), .A2(n_312), .B(n_319), .C(n_342), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_237), .A2(n_276), .B1(n_603), .B2(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g1019 ( .A(n_238), .Y(n_1019) );
INVxp67_ASAP7_75t_SL g1258 ( .A(n_239), .Y(n_1258) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_240), .Y(n_650) );
BUFx3_ASAP7_75t_L g302 ( .A(n_242), .Y(n_302) );
INVx1_ASAP7_75t_L g318 ( .A(n_242), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g1165 ( .A(n_243), .Y(n_1165) );
INVx1_ASAP7_75t_L g575 ( .A(n_246), .Y(n_575) );
INVx1_ASAP7_75t_L g790 ( .A(n_247), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_248), .Y(n_798) );
INVx1_ASAP7_75t_L g910 ( .A(n_249), .Y(n_910) );
INVxp67_ASAP7_75t_SL g986 ( .A(n_250), .Y(n_986) );
INVx1_ASAP7_75t_L g1217 ( .A(n_251), .Y(n_1217) );
OAI211xp5_ASAP7_75t_L g1225 ( .A1(n_251), .A2(n_1226), .B(n_1227), .C(n_1229), .Y(n_1225) );
INVx1_ASAP7_75t_L g733 ( .A(n_254), .Y(n_733) );
INVx1_ASAP7_75t_L g1518 ( .A(n_255), .Y(n_1518) );
INVx2_ASAP7_75t_L g380 ( .A(n_256), .Y(n_380) );
INVx1_ASAP7_75t_L g393 ( .A(n_256), .Y(n_393) );
INVx1_ASAP7_75t_L g398 ( .A(n_256), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g1326 ( .A1(n_257), .A2(n_271), .B1(n_1288), .B2(n_1293), .Y(n_1326) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_258), .Y(n_816) );
INVx1_ASAP7_75t_L g915 ( .A(n_260), .Y(n_915) );
INVx1_ASAP7_75t_L g1339 ( .A(n_261), .Y(n_1339) );
INVx1_ASAP7_75t_L g1026 ( .A(n_262), .Y(n_1026) );
INVx1_ASAP7_75t_L g850 ( .A(n_263), .Y(n_850) );
INVx1_ASAP7_75t_L g849 ( .A(n_264), .Y(n_849) );
INVx1_ASAP7_75t_L g465 ( .A(n_265), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g1563 ( .A1(n_267), .A2(n_1564), .B1(n_1565), .B2(n_1566), .Y(n_1563) );
CKINVDCx5p33_ASAP7_75t_R g1564 ( .A(n_267), .Y(n_1564) );
CKINVDCx5p33_ASAP7_75t_R g865 ( .A(n_269), .Y(n_865) );
INVx1_ASAP7_75t_L g1023 ( .A(n_270), .Y(n_1023) );
XOR2x2_ASAP7_75t_L g1166 ( .A(n_274), .B(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g1571 ( .A(n_275), .Y(n_1571) );
INVx1_ASAP7_75t_L g1570 ( .A(n_280), .Y(n_1570) );
OAI211xp5_ASAP7_75t_L g1534 ( .A1(n_281), .A2(n_614), .B(n_1214), .C(n_1535), .Y(n_1534) );
INVx1_ASAP7_75t_L g1552 ( .A(n_281), .Y(n_1552) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_303), .B(n_1278), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_289), .Y(n_283) );
INVx1_ASAP7_75t_L g1560 ( .A(n_284), .Y(n_1560) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g1608 ( .A(n_285), .B(n_288), .Y(n_1608) );
INVx1_ASAP7_75t_L g1610 ( .A(n_285), .Y(n_1610) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g1613 ( .A(n_288), .B(n_1610), .Y(n_1613) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x4_ASAP7_75t_L g488 ( .A(n_291), .B(n_489), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g1559 ( .A(n_291), .B(n_1560), .Y(n_1559) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g331 ( .A(n_292), .B(n_302), .Y(n_331) );
AND2x4_ASAP7_75t_L g374 ( .A(n_292), .B(n_301), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_293), .A2(n_504), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
INVx1_ASAP7_75t_L g1125 ( .A(n_293), .Y(n_1125) );
AND2x4_ASAP7_75t_SL g1558 ( .A(n_293), .B(n_1559), .Y(n_1558) );
INVxp67_ASAP7_75t_SL g1577 ( .A(n_293), .Y(n_1577) );
INVx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x6_ASAP7_75t_L g294 ( .A(n_295), .B(n_300), .Y(n_294) );
OR2x6_ASAP7_75t_L g494 ( .A(n_295), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g1207 ( .A(n_295), .Y(n_1207) );
OR2x2_ASAP7_75t_L g1554 ( .A(n_295), .B(n_495), .Y(n_1554) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx3_ASAP7_75t_L g364 ( .A(n_296), .Y(n_364) );
BUFx4f_ASAP7_75t_L g907 ( .A(n_296), .Y(n_907) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx2_ASAP7_75t_L g316 ( .A(n_298), .Y(n_316) );
AND2x2_ASAP7_75t_L g323 ( .A(n_298), .B(n_299), .Y(n_323) );
AND2x2_ASAP7_75t_L g328 ( .A(n_298), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g336 ( .A(n_298), .Y(n_336) );
INVx1_ASAP7_75t_L g406 ( .A(n_298), .Y(n_406) );
NAND2x1_ASAP7_75t_L g509 ( .A(n_298), .B(n_299), .Y(n_509) );
AND2x2_ASAP7_75t_L g315 ( .A(n_299), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g329 ( .A(n_299), .Y(n_329) );
INVx1_ASAP7_75t_L g337 ( .A(n_299), .Y(n_337) );
BUFx2_ASAP7_75t_L g359 ( .A(n_299), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_299), .B(n_316), .Y(n_368) );
OR2x2_ASAP7_75t_L g572 ( .A(n_299), .B(n_336), .Y(n_572) );
OR2x6_ASAP7_75t_L g1543 ( .A(n_300), .B(n_364), .Y(n_1543) );
INVxp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g519 ( .A(n_301), .Y(n_519) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx2_ASAP7_75t_L g501 ( .A(n_302), .Y(n_501) );
AND2x4_ASAP7_75t_L g515 ( .A(n_302), .B(n_405), .Y(n_515) );
OAI21xp33_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_1011), .B(n_1277), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_770), .B1(n_1009), .B2(n_1010), .Y(n_304) );
INVx2_ASAP7_75t_SL g1009 ( .A(n_305), .Y(n_1009) );
OAI221xp5_ASAP7_75t_L g1277 ( .A1(n_305), .A2(n_770), .B1(n_1009), .B2(n_1010), .C(n_1011), .Y(n_1277) );
AO22x1_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B1(n_619), .B2(n_620), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
XNOR2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_485), .Y(n_307) );
NAND3xp33_ASAP7_75t_L g309 ( .A(n_310), .B(n_381), .C(n_425), .Y(n_309) );
OAI21xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_350), .B(n_375), .Y(n_310) );
INVx2_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
INVx3_ASAP7_75t_L g1089 ( .A(n_313), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_313), .A2(n_348), .B1(n_1249), .B2(n_1250), .Y(n_1248) );
AND2x4_ASAP7_75t_L g313 ( .A(n_314), .B(n_317), .Y(n_313) );
INVx1_ASAP7_75t_L g990 ( .A(n_314), .Y(n_990) );
BUFx2_ASAP7_75t_L g1067 ( .A(n_314), .Y(n_1067) );
HB1xp67_ASAP7_75t_L g1099 ( .A(n_314), .Y(n_1099) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g339 ( .A(n_315), .Y(n_339) );
BUFx3_ASAP7_75t_L g661 ( .A(n_315), .Y(n_661) );
BUFx3_ASAP7_75t_L g682 ( .A(n_315), .Y(n_682) );
AND2x2_ASAP7_75t_L g345 ( .A(n_317), .B(n_335), .Y(n_345) );
AND2x4_ASAP7_75t_L g348 ( .A(n_317), .B(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_SL g354 ( .A(n_317), .B(n_322), .Y(n_354) );
AND2x2_ASAP7_75t_L g640 ( .A(n_317), .B(n_349), .Y(n_640) );
AND2x2_ASAP7_75t_L g684 ( .A(n_317), .B(n_338), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_317), .B(n_398), .Y(n_783) );
BUFx2_ASAP7_75t_L g891 ( .A(n_317), .Y(n_891) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_318), .Y(n_495) );
AOI21xp5_ASAP7_75t_SL g319 ( .A1(n_320), .A2(n_332), .B(n_340), .Y(n_319) );
AOI222xp33_ASAP7_75t_L g1120 ( .A1(n_321), .A2(n_511), .B1(n_1029), .B2(n_1121), .C1(n_1122), .C2(n_1123), .Y(n_1120) );
AOI222xp33_ASAP7_75t_L g1572 ( .A1(n_321), .A2(n_1029), .B1(n_1549), .B2(n_1573), .C1(n_1574), .C2(n_1575), .Y(n_1572) );
BUFx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x6_ASAP7_75t_L g340 ( .A(n_322), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g372 ( .A(n_322), .Y(n_372) );
AND2x2_ASAP7_75t_L g518 ( .A(n_322), .B(n_519), .Y(n_518) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_322), .Y(n_657) );
BUFx3_ASAP7_75t_L g900 ( .A(n_322), .Y(n_900) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g672 ( .A(n_323), .Y(n_672) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g787 ( .A(n_325), .Y(n_787) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
HB1xp67_ASAP7_75t_L g1595 ( .A(n_326), .Y(n_1595) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g759 ( .A(n_327), .Y(n_759) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_328), .Y(n_349) );
AND2x4_ASAP7_75t_L g504 ( .A(n_328), .B(n_495), .Y(n_504) );
BUFx3_ASAP7_75t_L g1097 ( .A(n_328), .Y(n_1097) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_331), .B(n_585), .Y(n_584) );
INVx4_ASAP7_75t_L g679 ( .A(n_331), .Y(n_679) );
AND2x4_ASAP7_75t_L g805 ( .A(n_331), .B(n_585), .Y(n_805) );
OAI21xp33_ASAP7_75t_L g901 ( .A1(n_331), .A2(n_902), .B(n_903), .Y(n_901) );
OAI221xp5_ASAP7_75t_L g1004 ( .A1(n_331), .A2(n_508), .B1(n_903), .B2(n_1005), .C(n_1006), .Y(n_1004) );
AND2x2_ASAP7_75t_SL g1528 ( .A(n_331), .B(n_391), .Y(n_1528) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g660 ( .A(n_334), .Y(n_660) );
INVx2_ASAP7_75t_SL g664 ( .A(n_334), .Y(n_664) );
INVx1_ASAP7_75t_L g681 ( .A(n_334), .Y(n_681) );
INVx1_ASAP7_75t_L g1055 ( .A(n_334), .Y(n_1055) );
INVx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_335), .B(n_341), .Y(n_399) );
BUFx6f_ASAP7_75t_L g761 ( .A(n_335), .Y(n_761) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_336), .Y(n_667) );
AND2x4_ASAP7_75t_L g781 ( .A(n_338), .B(n_782), .Y(n_781) );
INVx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g932 ( .A(n_339), .Y(n_932) );
AOI211xp5_ASAP7_75t_SL g765 ( .A1(n_340), .A2(n_686), .B(n_722), .C(n_766), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g1094 ( .A1(n_340), .A2(n_1095), .B(n_1098), .Y(n_1094) );
AOI221xp5_ASAP7_75t_L g1239 ( .A1(n_340), .A2(n_686), .B1(n_1240), .B2(n_1241), .C(n_1242), .Y(n_1239) );
INVx1_ASAP7_75t_L g360 ( .A(n_341), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_341), .B(n_405), .Y(n_404) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_341), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_341), .B(n_380), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_344), .B1(n_346), .B2(n_347), .Y(n_342) );
INVx1_ASAP7_75t_L g751 ( .A(n_344), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_344), .A2(n_1091), .B1(n_1092), .B2(n_1093), .Y(n_1090) );
AOI221xp5_ASAP7_75t_SL g1243 ( .A1(n_344), .A2(n_1244), .B1(n_1245), .B2(n_1246), .C(n_1247), .Y(n_1243) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g630 ( .A(n_345), .B(n_631), .Y(n_630) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g754 ( .A(n_348), .Y(n_754) );
BUFx6f_ASAP7_75t_L g1093 ( .A(n_348), .Y(n_1093) );
INVx1_ASAP7_75t_L g656 ( .A(n_349), .Y(n_656) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_349), .Y(n_678) );
INVx2_ASAP7_75t_L g894 ( .A(n_349), .Y(n_894) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g1101 ( .A(n_352), .Y(n_1101) );
INVx4_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx3_ASAP7_75t_L g686 ( .A(n_354), .Y(n_686) );
BUFx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g1102 ( .A(n_357), .Y(n_1102) );
NOR2x1_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
INVx1_ASAP7_75t_L g668 ( .A(n_358), .Y(n_668) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g512 ( .A(n_359), .B(n_501), .Y(n_512) );
INVx1_ASAP7_75t_L g813 ( .A(n_359), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_359), .A2(n_666), .B1(n_861), .B2(n_878), .Y(n_898) );
BUFx2_ASAP7_75t_L g1001 ( .A(n_359), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_359), .B(n_501), .Y(n_1549) );
INVx1_ASAP7_75t_L g1002 ( .A(n_360), .Y(n_1002) );
OAI221xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B1(n_366), .B2(n_369), .C(n_370), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
BUFx3_ASAP7_75t_L g563 ( .A(n_364), .Y(n_563) );
BUFx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g500 ( .A(n_367), .B(n_501), .Y(n_500) );
INVx8_ASAP7_75t_L g568 ( .A(n_367), .Y(n_568) );
OR2x2_ASAP7_75t_L g1555 ( .A(n_367), .B(n_519), .Y(n_1555) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g658 ( .A(n_374), .Y(n_658) );
OAI221xp5_ASAP7_75t_L g884 ( .A1(n_374), .A2(n_885), .B1(n_886), .B2(n_887), .C(n_888), .Y(n_884) );
INVx1_ASAP7_75t_L g930 ( .A(n_374), .Y(n_930) );
OAI221xp5_ASAP7_75t_L g991 ( .A1(n_374), .A2(n_570), .B1(n_885), .B2(n_992), .C(n_993), .Y(n_991) );
OAI21xp5_ASAP7_75t_SL g1087 ( .A1(n_375), .A2(n_1088), .B(n_1100), .Y(n_1087) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI21xp33_ASAP7_75t_L g748 ( .A1(n_376), .A2(n_749), .B(n_765), .Y(n_748) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI31xp33_ASAP7_75t_L g880 ( .A1(n_378), .A2(n_881), .A3(n_889), .B(n_899), .Y(n_880) );
HB1xp67_ASAP7_75t_L g918 ( .A(n_378), .Y(n_918) );
OAI31xp33_ASAP7_75t_L g987 ( .A1(n_378), .A2(n_988), .A3(n_994), .B(n_1003), .Y(n_987) );
BUFx2_ASAP7_75t_L g1251 ( .A(n_378), .Y(n_1251) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND3x4_ASAP7_75t_L g428 ( .A(n_379), .B(n_423), .C(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx2_ASAP7_75t_L g453 ( .A(n_380), .Y(n_453) );
AOI21xp33_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_400), .B(n_401), .Y(n_381) );
AOI21xp33_ASAP7_75t_L g1082 ( .A1(n_382), .A2(n_1083), .B(n_1084), .Y(n_1082) );
AOI21xp5_ASAP7_75t_L g1268 ( .A1(n_382), .A2(n_1269), .B(n_1270), .Y(n_1268) );
INVx8_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_396), .Y(n_383) );
INVx1_ASAP7_75t_L g649 ( .A(n_384), .Y(n_649) );
OR2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_390), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_386), .Y(n_606) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx2_ASAP7_75t_L g547 ( .A(n_387), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_388), .Y(n_412) );
INVx2_ASAP7_75t_L g416 ( .A(n_388), .Y(n_416) );
AND2x4_ASAP7_75t_L g435 ( .A(n_388), .B(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g474 ( .A(n_388), .B(n_418), .Y(n_474) );
INVx1_ASAP7_75t_L g411 ( .A(n_389), .Y(n_411) );
INVx2_ASAP7_75t_L g436 ( .A(n_389), .Y(n_436) );
OR2x2_ASAP7_75t_L g408 ( .A(n_390), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g476 ( .A(n_390), .Y(n_476) );
INVx1_ASAP7_75t_L g479 ( .A(n_390), .Y(n_479) );
OR2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_394), .Y(n_390) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_391), .Y(n_553) );
INVx1_ASAP7_75t_L g586 ( .A(n_391), .Y(n_586) );
OR2x2_ASAP7_75t_L g592 ( .A(n_391), .B(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx2_ASAP7_75t_L g407 ( .A(n_392), .Y(n_407) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g840 ( .A(n_394), .Y(n_840) );
INVx3_ASAP7_75t_L g421 ( .A(n_395), .Y(n_421) );
BUFx3_ASAP7_75t_L g429 ( .A(n_395), .Y(n_429) );
NAND2xp33_ASAP7_75t_SL g593 ( .A(n_395), .B(n_423), .Y(n_593) );
INVx1_ASAP7_75t_L g779 ( .A(n_396), .Y(n_779) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_399), .Y(n_396) );
AND2x4_ASAP7_75t_L g464 ( .A(n_397), .B(n_420), .Y(n_464) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g618 ( .A(n_398), .Y(n_618) );
INVx2_ASAP7_75t_L g1236 ( .A(n_402), .Y(n_1236) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_408), .Y(n_402) );
AND2x4_ASAP7_75t_L g1085 ( .A(n_403), .B(n_408), .Y(n_1085) );
OR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_407), .Y(n_403) );
INVx1_ASAP7_75t_L g768 ( .A(n_404), .Y(n_768) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVxp67_ASAP7_75t_L g424 ( .A(n_407), .Y(n_424) );
INVx1_ASAP7_75t_L g489 ( .A(n_407), .Y(n_489) );
INVx1_ASAP7_75t_L g631 ( .A(n_407), .Y(n_631) );
INVx2_ASAP7_75t_L g651 ( .A(n_408), .Y(n_651) );
INVx4_ASAP7_75t_L g530 ( .A(n_409), .Y(n_530) );
INVx3_ASAP7_75t_L g853 ( .A(n_409), .Y(n_853) );
BUFx6f_ASAP7_75t_L g1142 ( .A(n_409), .Y(n_1142) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx3_ASAP7_75t_L g600 ( .A(n_410), .Y(n_600) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
BUFx2_ASAP7_75t_L g541 ( .A(n_411), .Y(n_541) );
AND2x4_ASAP7_75t_L g444 ( .A(n_412), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g463 ( .A(n_412), .Y(n_463) );
BUFx2_ASAP7_75t_L g537 ( .A(n_412), .Y(n_537) );
INVx3_ASAP7_75t_L g625 ( .A(n_413), .Y(n_625) );
INVx5_ASAP7_75t_L g911 ( .A(n_413), .Y(n_911) );
OR2x6_ASAP7_75t_L g413 ( .A(n_414), .B(n_424), .Y(n_413) );
OR2x2_ASAP7_75t_L g1086 ( .A(n_414), .B(n_424), .Y(n_1086) );
NAND2x1p5_ASAP7_75t_L g414 ( .A(n_415), .B(n_420), .Y(n_414) );
BUFx3_ASAP7_75t_L g433 ( .A(n_415), .Y(n_433) );
BUFx3_ASAP7_75t_L g700 ( .A(n_415), .Y(n_700) );
INVx8_ASAP7_75t_L g707 ( .A(n_415), .Y(n_707) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_415), .Y(n_831) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
AND2x4_ASAP7_75t_L g440 ( .A(n_416), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVxp67_ASAP7_75t_L g441 ( .A(n_419), .Y(n_441) );
AND2x6_ASAP7_75t_L g820 ( .A(n_420), .B(n_462), .Y(n_820) );
AND2x2_ASAP7_75t_L g822 ( .A(n_420), .B(n_469), .Y(n_822) );
INVx1_ASAP7_75t_L g828 ( .A(n_420), .Y(n_828) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
NAND2x1p5_ASAP7_75t_L g454 ( .A(n_421), .B(n_455), .Y(n_454) );
OR2x4_ASAP7_75t_L g524 ( .A(n_421), .B(n_474), .Y(n_524) );
INVx1_ASAP7_75t_L g527 ( .A(n_421), .Y(n_527) );
AND2x4_ASAP7_75t_L g532 ( .A(n_421), .B(n_435), .Y(n_532) );
OR2x6_ASAP7_75t_L g546 ( .A(n_421), .B(n_547), .Y(n_546) );
NAND3x1_ASAP7_75t_L g617 ( .A(n_421), .B(n_455), .C(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_423), .Y(n_551) );
NOR3xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_470), .C(n_481), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_427), .B(n_459), .Y(n_426) );
AOI33xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .A3(n_437), .B1(n_446), .B2(n_451), .B3(n_456), .Y(n_427) );
AOI33xp33_ASAP7_75t_L g866 ( .A1(n_428), .A2(n_451), .A3(n_867), .B1(n_869), .B2(n_870), .B3(n_873), .Y(n_866) );
NAND3xp33_ASAP7_75t_L g969 ( .A(n_428), .B(n_970), .C(n_971), .Y(n_969) );
BUFx3_ASAP7_75t_L g1041 ( .A(n_428), .Y(n_1041) );
AOI33xp33_ASAP7_75t_L g1073 ( .A1(n_428), .A2(n_451), .A3(n_1074), .B1(n_1075), .B2(n_1077), .B3(n_1078), .Y(n_1073) );
INVx3_ASAP7_75t_L g536 ( .A(n_429), .Y(n_536) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
BUFx3_ASAP7_75t_L g735 ( .A(n_433), .Y(n_735) );
INVx1_ASAP7_75t_L g745 ( .A(n_433), .Y(n_745) );
BUFx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g458 ( .A(n_435), .Y(n_458) );
BUFx2_ASAP7_75t_L g484 ( .A(n_435), .Y(n_484) );
BUFx2_ASAP7_75t_L g701 ( .A(n_435), .Y(n_701) );
BUFx2_ASAP7_75t_L g724 ( .A(n_435), .Y(n_724) );
BUFx3_ASAP7_75t_L g826 ( .A(n_435), .Y(n_826) );
BUFx2_ASAP7_75t_L g951 ( .A(n_435), .Y(n_951) );
INVx1_ASAP7_75t_L g445 ( .A(n_436), .Y(n_445) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g526 ( .A(n_439), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g691 ( .A(n_439), .Y(n_691) );
BUFx6f_ASAP7_75t_L g848 ( .A(n_439), .Y(n_848) );
INVx2_ASAP7_75t_L g1135 ( .A(n_439), .Y(n_1135) );
INVx1_ASAP7_75t_L g1146 ( .A(n_439), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_439), .B(n_527), .Y(n_1533) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_440), .Y(n_449) );
BUFx8_ASAP7_75t_L g480 ( .A(n_440), .Y(n_480) );
INVx2_ASAP7_75t_L g604 ( .A(n_440), .Y(n_604) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_R g1076 ( .A(n_443), .Y(n_1076) );
INVx1_ASAP7_75t_L g1605 ( .A(n_443), .Y(n_1605) );
INVx5_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx3_ASAP7_75t_L g450 ( .A(n_444), .Y(n_450) );
BUFx12f_ASAP7_75t_L g704 ( .A(n_444), .Y(n_704) );
BUFx3_ASAP7_75t_L g836 ( .A(n_444), .Y(n_836) );
INVx1_ASAP7_75t_L g469 ( .A(n_445), .Y(n_469) );
INVx8_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx3_ASAP7_75t_L g1255 ( .A(n_448), .Y(n_1255) );
INVx5_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_449), .Y(n_609) );
INVx3_ASAP7_75t_L g833 ( .A(n_449), .Y(n_833) );
INVx2_ASAP7_75t_SL g872 ( .A(n_449), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_449), .A2(n_868), .B1(n_958), .B2(n_959), .Y(n_957) );
NAND3xp33_ASAP7_75t_L g978 ( .A(n_451), .B(n_979), .C(n_980), .Y(n_978) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR2x6_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
AND2x4_ASAP7_75t_L g557 ( .A(n_453), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g688 ( .A(n_453), .Y(n_688) );
OR2x2_ASAP7_75t_L g1515 ( .A(n_453), .B(n_454), .Y(n_1515) );
INVx3_ASAP7_75t_L g845 ( .A(n_454), .Y(n_845) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g708 ( .A(n_458), .Y(n_708) );
INVx1_ASAP7_75t_L g736 ( .A(n_458), .Y(n_736) );
INVx2_ASAP7_75t_L g946 ( .A(n_458), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B1(n_465), .B2(n_466), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_461), .A2(n_466), .B1(n_1080), .B2(n_1081), .Y(n_1079) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
AND2x4_ASAP7_75t_SL g644 ( .A(n_462), .B(n_464), .Y(n_644) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x4_ASAP7_75t_L g466 ( .A(n_464), .B(n_467), .Y(n_466) );
AND2x4_ASAP7_75t_L g483 ( .A(n_464), .B(n_484), .Y(n_483) );
AND2x4_ASAP7_75t_SL g646 ( .A(n_464), .B(n_467), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g1271 ( .A1(n_466), .A2(n_483), .B1(n_644), .B2(n_1242), .C(n_1272), .Y(n_1271) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_475), .Y(n_471) );
INVx2_ASAP7_75t_SL g613 ( .A(n_472), .Y(n_613) );
OR2x6_ASAP7_75t_L g632 ( .A(n_472), .B(n_475), .Y(n_632) );
INVx2_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OR2x4_ASAP7_75t_L g544 ( .A(n_474), .B(n_527), .Y(n_544) );
BUFx4f_ASAP7_75t_L g597 ( .A(n_474), .Y(n_597) );
BUFx3_ASAP7_75t_L g844 ( .A(n_474), .Y(n_844) );
BUFx3_ASAP7_75t_L g1261 ( .A(n_474), .Y(n_1261) );
INVxp67_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g636 ( .A(n_476), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_478), .B(n_875), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_478), .B(n_973), .Y(n_972) );
AND2x4_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
AND2x4_ASAP7_75t_L g862 ( .A(n_479), .B(n_863), .Y(n_862) );
AND2x4_ASAP7_75t_L g1275 ( .A(n_479), .B(n_863), .Y(n_1275) );
INVx3_ASAP7_75t_L g1604 ( .A(n_480), .Y(n_1604) );
NOR3xp33_ASAP7_75t_L g1070 ( .A(n_481), .B(n_1071), .C(n_1072), .Y(n_1070) );
INVx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
OAI211xp5_ASAP7_75t_SL g689 ( .A1(n_482), .A2(n_591), .B(n_690), .C(n_702), .Y(n_689) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g877 ( .A1(n_483), .A2(n_644), .B1(n_646), .B2(n_878), .C(n_879), .Y(n_877) );
AOI221xp5_ASAP7_75t_L g982 ( .A1(n_483), .A2(n_644), .B1(n_646), .B2(n_983), .C(n_984), .Y(n_982) );
OAI221xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_490), .B1(n_520), .B2(n_548), .C(n_554), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g1016 ( .A1(n_488), .A2(n_549), .B1(n_1017), .B2(n_1031), .Y(n_1016) );
BUFx2_ASAP7_75t_L g1126 ( .A(n_488), .Y(n_1126) );
BUFx2_ASAP7_75t_SL g1230 ( .A(n_488), .Y(n_1230) );
NOR3xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_502), .C(n_505), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g1569 ( .A1(n_497), .A2(n_1020), .B1(n_1570), .B2(n_1571), .Y(n_1569) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_499), .A2(n_1019), .B1(n_1020), .B2(n_1021), .Y(n_1018) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g1119 ( .A(n_500), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_501), .B(n_761), .Y(n_1020) );
INVx3_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g1222 ( .A(n_504), .Y(n_1222) );
INVx4_ASAP7_75t_L g1544 ( .A(n_504), .Y(n_1544) );
OAI22xp33_ASAP7_75t_L g1203 ( .A1(n_506), .A2(n_1177), .B1(n_1183), .B2(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g885 ( .A(n_507), .Y(n_885) );
INVx2_ASAP7_75t_L g1105 ( .A(n_507), .Y(n_1105) );
INVx2_ASAP7_75t_L g1526 ( .A(n_507), .Y(n_1526) );
INVx4_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx4f_ASAP7_75t_L g574 ( .A(n_508), .Y(n_574) );
BUFx4f_ASAP7_75t_L g801 ( .A(n_508), .Y(n_801) );
OR2x6_ASAP7_75t_L g806 ( .A(n_508), .B(n_807), .Y(n_806) );
BUFx6f_ASAP7_75t_L g939 ( .A(n_508), .Y(n_939) );
BUFx4f_ASAP7_75t_L g1151 ( .A(n_508), .Y(n_1151) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx3_ASAP7_75t_L g580 ( .A(n_509), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_513), .B1(n_514), .B2(n_516), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g1227 ( .A1(n_511), .A2(n_514), .B1(n_1216), .B2(n_1228), .Y(n_1227) );
BUFx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AOI222xp33_ASAP7_75t_L g1025 ( .A1(n_512), .A2(n_900), .B1(n_1026), .B2(n_1027), .C1(n_1028), .C2(n_1029), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_513), .A2(n_534), .B1(n_538), .B2(n_539), .Y(n_533) );
BUFx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g1030 ( .A(n_515), .Y(n_1030) );
INVx2_ASAP7_75t_L g1551 ( .A(n_515), .Y(n_1551) );
NAND4xp25_ASAP7_75t_L g1017 ( .A(n_517), .B(n_1018), .C(n_1022), .D(n_1025), .Y(n_1017) );
NAND3xp33_ASAP7_75t_L g1114 ( .A(n_517), .B(n_1115), .C(n_1120), .Y(n_1114) );
NAND3xp33_ASAP7_75t_L g1568 ( .A(n_517), .B(n_1569), .C(n_1572), .Y(n_1568) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g1229 ( .A(n_518), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1547 ( .A(n_519), .B(n_1065), .Y(n_1547) );
NOR3xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_528), .C(n_542), .Y(n_520) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_523), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_523), .A2(n_526), .B1(n_1023), .B2(n_1024), .Y(n_1039) );
INVx2_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g1162 ( .A(n_524), .Y(n_1162) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_526), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_715) );
INVx2_ASAP7_75t_L g1163 ( .A(n_526), .Y(n_1163) );
INVx1_ASAP7_75t_L g1219 ( .A(n_526), .Y(n_1219) );
INVxp67_ASAP7_75t_L g1580 ( .A(n_526), .Y(n_1580) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g843 ( .A(n_530), .Y(n_843) );
NAND4xp25_ASAP7_75t_L g714 ( .A(n_531), .B(n_715), .C(n_719), .D(n_725), .Y(n_714) );
NAND3xp33_ASAP7_75t_L g1157 ( .A(n_531), .B(n_1158), .C(n_1159), .Y(n_1157) );
CKINVDCx8_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
OAI31xp33_ASAP7_75t_L g953 ( .A1(n_532), .A2(n_954), .A3(n_964), .B(n_965), .Y(n_953) );
AOI211xp5_ASAP7_75t_L g1032 ( .A1(n_532), .A2(n_736), .B(n_1028), .C(n_1033), .Y(n_1032) );
CKINVDCx8_ASAP7_75t_R g1214 ( .A(n_532), .Y(n_1214) );
AOI22xp33_ASAP7_75t_L g1583 ( .A1(n_534), .A2(n_539), .B1(n_1574), .B2(n_1575), .Y(n_1583) );
BUFx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx3_ASAP7_75t_L g721 ( .A(n_535), .Y(n_721) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
AND2x4_ASAP7_75t_L g540 ( .A(n_536), .B(n_541), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g954 ( .A1(n_536), .A2(n_955), .B(n_957), .C(n_960), .Y(n_954) );
AND2x4_ASAP7_75t_L g962 ( .A(n_536), .B(n_537), .Y(n_962) );
AND2x4_ASAP7_75t_L g1536 ( .A(n_536), .B(n_537), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1538 ( .A(n_536), .B(n_541), .Y(n_1538) );
AOI222xp33_ASAP7_75t_L g719 ( .A1(n_539), .A2(n_720), .B1(n_721), .B2(n_722), .C1(n_723), .C2(n_724), .Y(n_719) );
AOI222xp33_ASAP7_75t_L g1158 ( .A1(n_539), .A2(n_721), .B1(n_746), .B2(n_1121), .C1(n_1122), .C2(n_1123), .Y(n_1158) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g960 ( .A1(n_540), .A2(n_961), .B1(n_962), .B2(n_963), .Y(n_960) );
INVx1_ASAP7_75t_L g1035 ( .A(n_540), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g1215 ( .A1(n_540), .A2(n_962), .B1(n_1216), .B2(n_1217), .Y(n_1215) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_SL g728 ( .A(n_544), .Y(n_728) );
BUFx3_ASAP7_75t_L g1038 ( .A(n_544), .Y(n_1038) );
BUFx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g718 ( .A(n_546), .Y(n_718) );
INVx1_ASAP7_75t_L g695 ( .A(n_547), .Y(n_695) );
BUFx3_ASAP7_75t_L g1137 ( .A(n_547), .Y(n_1137) );
CKINVDCx14_ASAP7_75t_R g548 ( .A(n_549), .Y(n_548) );
AOI211xp5_ASAP7_75t_L g713 ( .A1(n_549), .A2(n_714), .B(n_729), .C(n_748), .Y(n_713) );
OAI31xp33_ASAP7_75t_L g1578 ( .A1(n_549), .A2(n_1579), .A3(n_1582), .B(n_1584), .Y(n_1578) );
AND2x4_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
AND2x2_ASAP7_75t_L g965 ( .A(n_550), .B(n_552), .Y(n_965) );
AND2x2_ASAP7_75t_SL g1164 ( .A(n_550), .B(n_552), .Y(n_1164) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_590), .Y(n_554) );
OAI33xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_559), .A3(n_569), .B1(n_576), .B2(n_582), .B3(n_587), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g795 ( .A(n_557), .Y(n_795) );
INVx2_ASAP7_75t_L g1053 ( .A(n_557), .Y(n_1053) );
INVx2_ASAP7_75t_L g1189 ( .A(n_557), .Y(n_1189) );
INVx4_ASAP7_75t_L g1592 ( .A(n_557), .Y(n_1592) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B1(n_564), .B2(n_565), .Y(n_559) );
OAI22xp33_ASAP7_75t_L g594 ( .A1(n_560), .A2(n_577), .B1(n_595), .B2(n_598), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_561), .A2(n_565), .B1(n_588), .B2(n_589), .Y(n_587) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_563), .A2(n_790), .B1(n_791), .B2(n_793), .Y(n_789) );
OAI22xp33_ASAP7_75t_L g611 ( .A1(n_564), .A2(n_581), .B1(n_612), .B2(n_614), .Y(n_611) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_567), .A2(n_905), .B1(n_906), .B2(n_908), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g1529 ( .A1(n_567), .A2(n_906), .B1(n_1507), .B2(n_1518), .Y(n_1529) );
INVx4_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g792 ( .A(n_568), .Y(n_792) );
INVx2_ASAP7_75t_L g997 ( .A(n_568), .Y(n_997) );
INVx2_ASAP7_75t_SL g1195 ( .A(n_568), .Y(n_1195) );
INVx1_ASAP7_75t_L g1521 ( .A(n_568), .Y(n_1521) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_573), .B1(n_574), .B2(n_575), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_570), .A2(n_577), .B1(n_578), .B2(n_581), .Y(n_576) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g888 ( .A(n_571), .Y(n_888) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g800 ( .A(n_572), .Y(n_800) );
BUFx3_ASAP7_75t_L g903 ( .A(n_572), .Y(n_903) );
BUFx2_ASAP7_75t_L g1199 ( .A(n_572), .Y(n_1199) );
BUFx2_ASAP7_75t_L g1523 ( .A(n_572), .Y(n_1523) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_573), .A2(n_588), .B1(n_602), .B2(n_605), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_575), .A2(n_589), .B1(n_608), .B2(n_610), .Y(n_607) );
OAI211xp5_ASAP7_75t_L g675 ( .A1(n_578), .A2(n_676), .B(n_677), .C(n_680), .Y(n_675) );
INVx5_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
BUFx3_ASAP7_75t_L g757 ( .A(n_580), .Y(n_757) );
OR2x2_ASAP7_75t_L g784 ( .A(n_580), .B(n_783), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_580), .B(n_898), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_580), .B(n_1000), .Y(n_999) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OAI33xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_594), .A3(n_601), .B1(n_607), .B2(n_611), .B3(n_615), .Y(n_590) );
BUFx4f_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
BUFx4f_ASAP7_75t_L g738 ( .A(n_592), .Y(n_738) );
BUFx2_ASAP7_75t_L g855 ( .A(n_593), .Y(n_855) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
HB1xp67_ASAP7_75t_L g1172 ( .A(n_597), .Y(n_1172) );
HB1xp67_ASAP7_75t_L g1185 ( .A(n_597), .Y(n_1185) );
OAI22xp5_ASAP7_75t_SL g1508 ( .A1(n_597), .A2(n_1509), .B1(n_1510), .B2(n_1511), .Y(n_1508) );
OAI22xp33_ASAP7_75t_L g1512 ( .A1(n_597), .A2(n_600), .B1(n_1513), .B2(n_1514), .Y(n_1512) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g1132 ( .A(n_599), .Y(n_1132) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_600), .Y(n_614) );
OAI221xp5_ASAP7_75t_L g730 ( .A1(n_602), .A2(n_731), .B1(n_732), .B2(n_733), .C(n_734), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g1179 ( .A1(n_602), .A2(n_1180), .B1(n_1181), .B2(n_1183), .Y(n_1179) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx3_ASAP7_75t_L g637 ( .A(n_604), .Y(n_637) );
BUFx2_ASAP7_75t_L g740 ( .A(n_604), .Y(n_740) );
INVx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx3_ASAP7_75t_L g610 ( .A(n_606), .Y(n_610) );
CKINVDCx8_ASAP7_75t_R g732 ( .A(n_606), .Y(n_732) );
INVx3_ASAP7_75t_L g1148 ( .A(n_606), .Y(n_1148) );
INVx1_ASAP7_75t_L g1265 ( .A(n_606), .Y(n_1265) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI221xp5_ASAP7_75t_L g739 ( .A1(n_610), .A2(n_740), .B1(n_741), .B2(n_742), .C(n_743), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g1505 ( .A1(n_610), .A2(n_833), .B1(n_1506), .B2(n_1507), .Y(n_1505) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI22xp33_ASAP7_75t_L g1170 ( .A1(n_614), .A2(n_1171), .B1(n_1172), .B2(n_1173), .Y(n_1170) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_614), .A2(n_1258), .B1(n_1259), .B2(n_1262), .Y(n_1257) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_615), .A2(n_730), .B1(n_737), .B2(n_739), .Y(n_729) );
OAI33xp33_ASAP7_75t_L g1169 ( .A1(n_615), .A2(n_737), .A3(n_1170), .B1(n_1174), .B2(n_1179), .B3(n_1184), .Y(n_1169) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_616), .B(n_703), .C(n_705), .Y(n_702) );
INVx2_ASAP7_75t_L g952 ( .A(n_616), .Y(n_952) );
CKINVDCx5p33_ASAP7_75t_R g1143 ( .A(n_616), .Y(n_1143) );
NAND3xp33_ASAP7_75t_L g1601 ( .A(n_616), .B(n_1602), .C(n_1606), .Y(n_1601) );
INVx3_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx3_ASAP7_75t_L g1047 ( .A(n_617), .Y(n_1047) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
XOR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_711), .Y(n_620) );
INVx1_ASAP7_75t_L g709 ( .A(n_622), .Y(n_709) );
NAND3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_626), .C(n_641), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_624), .A2(n_684), .B1(n_685), .B2(n_686), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B1(n_633), .B2(n_634), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_632), .Y(n_628) );
INVx3_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_630), .A2(n_639), .B1(n_815), .B2(n_816), .Y(n_814) );
AND2x4_ASAP7_75t_L g639 ( .A(n_631), .B(n_640), .Y(n_639) );
NAND2x1_ASAP7_75t_L g634 ( .A(n_635), .B(n_638), .Y(n_634) );
INVx2_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g948 ( .A(n_637), .Y(n_948) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR3xp33_ASAP7_75t_SL g641 ( .A(n_642), .B(n_652), .C(n_689), .Y(n_641) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B1(n_650), .B2(n_651), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_648), .B(n_664), .Y(n_663) );
AOI222xp33_ASAP7_75t_L g860 ( .A1(n_649), .A2(n_651), .B1(n_861), .B2(n_862), .C1(n_864), .C2(n_865), .Y(n_860) );
AOI222xp33_ASAP7_75t_L g974 ( .A1(n_649), .A2(n_651), .B1(n_862), .B2(n_975), .C1(n_976), .C2(n_977), .Y(n_974) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_650), .A2(n_666), .B1(n_668), .B2(n_669), .C(n_670), .Y(n_665) );
AOI31xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_675), .A3(n_683), .B(n_687), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_659), .B(n_662), .Y(n_653) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
BUFx2_ASAP7_75t_L g788 ( .A(n_657), .Y(n_788) );
AOI221xp5_ASAP7_75t_L g892 ( .A1(n_657), .A2(n_875), .B1(n_879), .B2(n_893), .C(n_895), .Y(n_892) );
AOI221xp5_ASAP7_75t_L g995 ( .A1(n_657), .A2(n_893), .B1(n_973), .B2(n_984), .C(n_996), .Y(n_995) );
INVx1_ASAP7_75t_SL g1057 ( .A(n_661), .Y(n_1057) );
BUFx3_ASAP7_75t_L g1589 ( .A(n_661), .Y(n_1589) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_665), .B(n_673), .Y(n_662) );
INVx1_ASAP7_75t_L g938 ( .A(n_666), .Y(n_938) );
AOI22xp5_ASAP7_75t_L g1000 ( .A1(n_666), .A2(n_975), .B1(n_983), .B2(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g937 ( .A(n_668), .Y(n_937) );
INVx1_ASAP7_75t_L g1061 ( .A(n_670), .Y(n_1061) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
BUFx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g1065 ( .A(n_672), .Y(n_1065) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g896 ( .A1(n_674), .A2(n_761), .B(n_865), .C(n_897), .Y(n_896) );
A2O1A1Ixp33_ASAP7_75t_SL g933 ( .A1(n_674), .A2(n_934), .B(n_935), .C(n_936), .Y(n_933) );
BUFx3_ASAP7_75t_L g1059 ( .A(n_678), .Y(n_1059) );
INVx2_ASAP7_75t_L g752 ( .A(n_684), .Y(n_752) );
OAI31xp67_ASAP7_75t_L g817 ( .A1(n_687), .A2(n_818), .A3(n_829), .B(n_841), .Y(n_817) );
BUFx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .B1(n_693), .B2(n_696), .C(n_697), .Y(n_690) );
INVx3_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
BUFx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g1178 ( .A(n_695), .Y(n_1178) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
BUFx2_ASAP7_75t_L g1043 ( .A(n_700), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_701), .A2(n_835), .B1(n_836), .B2(n_837), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_704), .A2(n_826), .B1(n_934), .B2(n_956), .Y(n_955) );
INVx3_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_707), .Y(n_825) );
INVx2_ASAP7_75t_L g863 ( .A(n_707), .Y(n_863) );
INVx8_ASAP7_75t_L g868 ( .A(n_707), .Y(n_868) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_718), .A2(n_1019), .B1(n_1021), .B2(n_1037), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_718), .A2(n_728), .B1(n_1116), .B2(n_1117), .Y(n_1159) );
INVx2_ASAP7_75t_L g1581 ( .A(n_718), .Y(n_1581) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_723), .B(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g747 ( .A(n_724), .Y(n_747) );
INVx2_ASAP7_75t_L g1211 ( .A(n_728), .Y(n_1211) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_732), .A2(n_847), .B1(n_849), .B2(n_850), .Y(n_846) );
OAI221xp5_ASAP7_75t_L g941 ( .A1(n_732), .A2(n_942), .B1(n_943), .B2(n_944), .C(n_945), .Y(n_941) );
OAI221xp5_ASAP7_75t_L g947 ( .A1(n_732), .A2(n_928), .B1(n_948), .B2(n_949), .C(n_950), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g1253 ( .A1(n_732), .A2(n_1254), .B1(n_1255), .B2(n_1256), .Y(n_1253) );
OAI22xp33_ASAP7_75t_L g940 ( .A1(n_737), .A2(n_941), .B1(n_947), .B2(n_952), .Y(n_940) );
OAI33xp33_ASAP7_75t_L g1128 ( .A1(n_737), .A2(n_1129), .A3(n_1133), .B1(n_1138), .B2(n_1143), .B3(n_1144), .Y(n_1128) );
BUFx3_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OAI33xp33_ASAP7_75t_L g1504 ( .A1(n_738), .A2(n_1505), .A3(n_1508), .B1(n_1512), .B2(n_1515), .B3(n_1516), .Y(n_1504) );
INVx2_ASAP7_75t_L g1599 ( .A(n_740), .Y(n_1599) );
OAI211xp5_ASAP7_75t_SL g762 ( .A1(n_741), .A2(n_757), .B(n_763), .C(n_764), .Y(n_762) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_753), .Y(n_749) );
OAI211xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B(n_758), .C(n_760), .Y(n_755) );
BUFx2_ASAP7_75t_L g1226 ( .A(n_757), .Y(n_1226) );
INVx3_ASAP7_75t_L g883 ( .A(n_761), .Y(n_883) );
BUFx6f_ASAP7_75t_L g935 ( .A(n_761), .Y(n_935) );
A2O1A1Ixp33_ASAP7_75t_L g998 ( .A1(n_761), .A2(n_977), .B(n_999), .C(n_1002), .Y(n_998) );
INVx3_ASAP7_75t_SL g1010 ( .A(n_770), .Y(n_1010) );
BUFx3_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
OA22x2_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .B1(n_913), .B2(n_1008), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
XOR2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_857), .Y(n_773) );
XNOR2x1_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
NAND4xp75_ASAP7_75t_L g776 ( .A(n_777), .B(n_785), .C(n_814), .D(n_817), .Y(n_776) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AOI211x1_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_794), .B(n_796), .C(n_810), .Y(n_785) );
BUFx6f_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
OAI221xp5_ASAP7_75t_L g842 ( .A1(n_793), .A2(n_802), .B1(n_843), .B2(n_844), .C(n_845), .Y(n_842) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_804), .B(n_806), .Y(n_796) );
OAI221xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .B1(n_801), .B2(n_802), .C(n_803), .Y(n_797) );
OAI211xp5_ASAP7_75t_L g851 ( .A1(n_798), .A2(n_852), .B(n_854), .C(n_856), .Y(n_851) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g1525 ( .A(n_800), .Y(n_1525) );
OAI211xp5_ASAP7_75t_SL g923 ( .A1(n_801), .A2(n_924), .B(n_925), .C(n_926), .Y(n_923) );
OAI211xp5_ASAP7_75t_SL g927 ( .A1(n_801), .A2(n_928), .B(n_929), .C(n_931), .Y(n_927) );
OAI22xp5_ASAP7_75t_L g1149 ( .A1(n_804), .A2(n_1052), .B1(n_1150), .B2(n_1154), .Y(n_1149) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
AOI33xp33_ASAP7_75t_L g1050 ( .A1(n_805), .A2(n_1051), .A3(n_1054), .B1(n_1058), .B2(n_1062), .B3(n_1066), .Y(n_1050) );
INVx2_ASAP7_75t_L g1208 ( .A(n_805), .Y(n_1208) );
NAND3xp33_ASAP7_75t_L g1593 ( .A(n_805), .B(n_1594), .C(n_1596), .Y(n_1593) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
NAND2x2_ASAP7_75t_L g811 ( .A(n_808), .B(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx2_ASAP7_75t_SL g812 ( .A(n_813), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_815), .A2(n_816), .B1(n_831), .B2(n_832), .Y(n_830) );
INVx4_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
A2O1A1Ixp33_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_825), .B(n_826), .C(n_827), .Y(n_823) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AOI21xp33_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_834), .B(n_838), .Y(n_829) );
INVx2_ASAP7_75t_L g1176 ( .A(n_832), .Y(n_1176) );
INVx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OAI21xp5_ASAP7_75t_SL g841 ( .A1(n_842), .A2(n_846), .B(n_851), .Y(n_841) );
OAI22xp33_ASAP7_75t_L g1129 ( .A1(n_844), .A2(n_1130), .B1(n_1131), .B2(n_1132), .Y(n_1129) );
OAI22xp33_ASAP7_75t_L g1138 ( .A1(n_844), .A2(n_1139), .B1(n_1140), .B2(n_1141), .Y(n_1138) );
OAI221xp5_ASAP7_75t_L g1263 ( .A1(n_847), .A2(n_1264), .B1(n_1265), .B2(n_1266), .C(n_1267), .Y(n_1263) );
INVx2_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx2_ASAP7_75t_SL g942 ( .A(n_848), .Y(n_942) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx2_ASAP7_75t_L g1213 ( .A(n_853), .Y(n_1213) );
INVx3_ASAP7_75t_L g1511 ( .A(n_853), .Y(n_1511) );
XNOR2x1_ASAP7_75t_L g857 ( .A(n_858), .B(n_912), .Y(n_857) );
OR2x2_ASAP7_75t_L g858 ( .A(n_859), .B(n_876), .Y(n_858) );
NAND3xp33_ASAP7_75t_L g859 ( .A(n_860), .B(n_866), .C(n_874), .Y(n_859) );
INVx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
OAI22xp5_ASAP7_75t_L g1516 ( .A1(n_872), .A2(n_1178), .B1(n_1517), .B2(n_1518), .Y(n_1516) );
NAND3xp33_ASAP7_75t_SL g876 ( .A(n_877), .B(n_880), .C(n_909), .Y(n_876) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx2_ASAP7_75t_SL g1153 ( .A(n_883), .Y(n_1153) );
OAI221xp5_ASAP7_75t_SL g1150 ( .A1(n_888), .A2(n_1134), .B1(n_1145), .B2(n_1151), .C(n_1152), .Y(n_1150) );
OAI221xp5_ASAP7_75t_SL g1154 ( .A1(n_888), .A2(n_1131), .B1(n_1140), .B2(n_1151), .C(n_1155), .Y(n_1154) );
OAI21xp33_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_892), .B(n_896), .Y(n_889) );
OAI21xp5_ASAP7_75t_SL g994 ( .A1(n_890), .A2(n_995), .B(n_998), .Y(n_994) );
INVxp67_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
OAI21xp5_ASAP7_75t_L g920 ( .A1(n_891), .A2(n_921), .B(n_922), .Y(n_920) );
INVx2_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx2_ASAP7_75t_L g1202 ( .A(n_903), .Y(n_1202) );
OAI22xp33_ASAP7_75t_L g1520 ( .A1(n_906), .A2(n_1509), .B1(n_1513), .B2(n_1521), .Y(n_1520) );
INVx4_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
BUFx6f_ASAP7_75t_L g1192 ( .A(n_907), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_910), .B(n_911), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_911), .B(n_986), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_911), .B(n_1250), .Y(n_1273) );
XNOR2xp5_ASAP7_75t_L g913 ( .A(n_914), .B(n_966), .Y(n_913) );
XOR2xp5_ASAP7_75t_L g1008 ( .A(n_914), .B(n_966), .Y(n_1008) );
XNOR2x1_ASAP7_75t_L g914 ( .A(n_915), .B(n_916), .Y(n_914) );
AND2x2_ASAP7_75t_L g916 ( .A(n_917), .B(n_953), .Y(n_916) );
AOI21xp5_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_919), .B(n_940), .Y(n_917) );
NAND4xp25_ASAP7_75t_L g919 ( .A(n_920), .B(n_923), .C(n_927), .D(n_933), .Y(n_919) );
HB1xp67_ASAP7_75t_L g1049 ( .A(n_951), .Y(n_1049) );
INVx1_ASAP7_75t_L g1034 ( .A(n_962), .Y(n_1034) );
OAI31xp33_ASAP7_75t_L g1530 ( .A1(n_965), .A2(n_1531), .A3(n_1534), .B(n_1540), .Y(n_1530) );
XNOR2x1_ASAP7_75t_L g966 ( .A(n_967), .B(n_1007), .Y(n_966) );
OR2x2_ASAP7_75t_L g967 ( .A(n_968), .B(n_981), .Y(n_967) );
NAND4xp25_ASAP7_75t_SL g968 ( .A(n_969), .B(n_972), .C(n_974), .D(n_978), .Y(n_968) );
NAND3xp33_ASAP7_75t_SL g981 ( .A(n_982), .B(n_985), .C(n_987), .Y(n_981) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
XNOR2xp5_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1108), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
XNOR2x1_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1068), .Y(n_1013) );
NAND3x1_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1040), .C(n_1050), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_1020), .A2(n_1116), .B1(n_1117), .B2(n_1118), .Y(n_1115) );
INVx2_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
NAND3xp33_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1036), .C(n_1039), .Y(n_1031) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
AOI33xp33_ASAP7_75t_L g1040 ( .A1(n_1041), .A2(n_1042), .A3(n_1044), .B1(n_1045), .B2(n_1046), .B3(n_1048), .Y(n_1040) );
NAND3xp33_ASAP7_75t_L g1597 ( .A(n_1041), .B(n_1598), .C(n_1600), .Y(n_1597) );
BUFx2_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
BUFx6f_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx1_ASAP7_75t_SL g1056 ( .A(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
INVx2_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
AND3x1_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1082), .C(n_1087), .Y(n_1069) );
NAND2xp5_ASAP7_75t_SL g1072 ( .A(n_1073), .B(n_1079), .Y(n_1072) );
HB1xp67_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
BUFx2_ASAP7_75t_L g1588 ( .A(n_1097), .Y(n_1588) );
OAI211xp5_ASAP7_75t_SL g1103 ( .A1(n_1104), .A2(n_1105), .B(n_1106), .C(n_1107), .Y(n_1103) );
XOR2xp5_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1232), .Y(n_1108) );
AOI22xp5_ASAP7_75t_L g1109 ( .A1(n_1110), .A2(n_1111), .B1(n_1166), .B2(n_1231), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
XOR2x2_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1165), .Y(n_1111) );
NAND3x1_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1127), .C(n_1156), .Y(n_1112) );
OAI21xp5_ASAP7_75t_L g1113 ( .A1(n_1114), .A2(n_1124), .B(n_1126), .Y(n_1113) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1118), .Y(n_1224) );
INVx2_ASAP7_75t_SL g1118 ( .A(n_1119), .Y(n_1118) );
OAI31xp33_ASAP7_75t_SL g1541 ( .A1(n_1126), .A2(n_1542), .A3(n_1545), .B(n_1553), .Y(n_1541) );
OAI21xp5_ASAP7_75t_L g1567 ( .A1(n_1126), .A2(n_1568), .B(n_1576), .Y(n_1567) );
NOR2x1_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1149), .Y(n_1127) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_1134), .A2(n_1135), .B1(n_1136), .B2(n_1137), .Y(n_1133) );
HB1xp67_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1142), .Y(n_1182) );
OAI22xp5_ASAP7_75t_L g1144 ( .A1(n_1145), .A2(n_1146), .B1(n_1147), .B2(n_1148), .Y(n_1144) );
OAI22xp5_ASAP7_75t_L g1184 ( .A1(n_1148), .A2(n_1185), .B1(n_1186), .B2(n_1187), .Y(n_1184) );
OAI22xp5_ASAP7_75t_L g1196 ( .A1(n_1151), .A2(n_1175), .B1(n_1180), .B2(n_1197), .Y(n_1196) );
OAI22xp5_ASAP7_75t_L g1522 ( .A1(n_1151), .A2(n_1506), .B1(n_1517), .B2(n_1523), .Y(n_1522) );
OAI21xp33_ASAP7_75t_L g1156 ( .A1(n_1157), .A2(n_1160), .B(n_1164), .Y(n_1156) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
OAI31xp33_ASAP7_75t_SL g1209 ( .A1(n_1164), .A2(n_1210), .A3(n_1212), .B(n_1218), .Y(n_1209) );
INVx2_ASAP7_75t_SL g1231 ( .A(n_1166), .Y(n_1231) );
NAND3xp33_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1209), .C(n_1220), .Y(n_1167) );
NOR2xp33_ASAP7_75t_SL g1168 ( .A(n_1169), .B(n_1188), .Y(n_1168) );
OAI22xp5_ASAP7_75t_L g1190 ( .A1(n_1171), .A2(n_1186), .B1(n_1191), .B2(n_1193), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g1200 ( .A1(n_1173), .A2(n_1187), .B1(n_1193), .B2(n_1201), .Y(n_1200) );
OAI22xp33_ASAP7_75t_SL g1174 ( .A1(n_1175), .A2(n_1176), .B1(n_1177), .B2(n_1178), .Y(n_1174) );
INVx2_ASAP7_75t_SL g1181 ( .A(n_1182), .Y(n_1181) );
OAI33xp33_ASAP7_75t_L g1188 ( .A1(n_1189), .A2(n_1190), .A3(n_1196), .B1(n_1200), .B2(n_1203), .B3(n_1208), .Y(n_1188) );
OAI33xp33_ASAP7_75t_L g1519 ( .A1(n_1189), .A2(n_1520), .A3(n_1522), .B1(n_1524), .B2(n_1527), .B3(n_1529), .Y(n_1519) );
INVx2_ASAP7_75t_SL g1191 ( .A(n_1192), .Y(n_1191) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
INVx2_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
INVx4_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
INVx3_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
OAI31xp33_ASAP7_75t_L g1220 ( .A1(n_1221), .A2(n_1223), .A3(n_1225), .B(n_1230), .Y(n_1220) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
XNOR2xp5_ASAP7_75t_L g1233 ( .A(n_1234), .B(n_1276), .Y(n_1233) );
NAND2xp5_ASAP7_75t_SL g1234 ( .A(n_1235), .B(n_1268), .Y(n_1234) );
AOI221xp5_ASAP7_75t_L g1235 ( .A1(n_1236), .A2(n_1237), .B1(n_1238), .B2(n_1251), .C(n_1252), .Y(n_1235) );
NAND3xp33_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1243), .C(n_1248), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1246), .B(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
INVxp67_ASAP7_75t_SL g1260 ( .A(n_1261), .Y(n_1260) );
NAND3xp33_ASAP7_75t_L g1270 ( .A(n_1271), .B(n_1273), .C(n_1274), .Y(n_1270) );
OAI221xp5_ASAP7_75t_L g1278 ( .A1(n_1279), .A2(n_1497), .B1(n_1499), .B2(n_1556), .C(n_1561), .Y(n_1278) );
AND3x1_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1426), .C(n_1462), .Y(n_1279) );
NOR3xp33_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1357), .C(n_1415), .Y(n_1280) );
OAI221xp5_ASAP7_75t_L g1281 ( .A1(n_1282), .A2(n_1284), .B1(n_1334), .B2(n_1347), .C(n_1350), .Y(n_1281) );
AOI221xp5_ASAP7_75t_L g1282 ( .A1(n_1283), .A2(n_1309), .B1(n_1315), .B2(n_1324), .C(n_1328), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1300), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1374 ( .A(n_1285), .B(n_1375), .Y(n_1374) );
CKINVDCx5p33_ASAP7_75t_R g1410 ( .A(n_1285), .Y(n_1410) );
NAND2xp5_ASAP7_75t_L g1428 ( .A(n_1285), .B(n_1429), .Y(n_1428) );
OAI211xp5_ASAP7_75t_SL g1463 ( .A1(n_1285), .A2(n_1464), .B(n_1467), .C(n_1479), .Y(n_1463) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1285), .B(n_1361), .Y(n_1476) );
NOR2xp33_ASAP7_75t_L g1494 ( .A(n_1285), .B(n_1495), .Y(n_1494) );
INVx4_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
INVx4_ASAP7_75t_L g1317 ( .A(n_1286), .Y(n_1317) );
NAND2xp5_ASAP7_75t_SL g1332 ( .A(n_1286), .B(n_1333), .Y(n_1332) );
OR2x2_ASAP7_75t_L g1365 ( .A(n_1286), .B(n_1333), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1286), .B(n_1418), .Y(n_1417) );
NOR2xp33_ASAP7_75t_L g1425 ( .A(n_1286), .B(n_1349), .Y(n_1425) );
NAND2xp5_ASAP7_75t_L g1472 ( .A(n_1286), .B(n_1385), .Y(n_1472) );
AND2x4_ASAP7_75t_SL g1286 ( .A(n_1287), .B(n_1295), .Y(n_1286) );
AND2x4_ASAP7_75t_L g1288 ( .A(n_1289), .B(n_1290), .Y(n_1288) );
AND2x6_ASAP7_75t_L g1293 ( .A(n_1289), .B(n_1294), .Y(n_1293) );
AND2x6_ASAP7_75t_L g1296 ( .A(n_1289), .B(n_1297), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1289), .B(n_1299), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1289), .B(n_1299), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1338 ( .A(n_1289), .B(n_1290), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1289), .B(n_1299), .Y(n_1343) );
HB1xp67_ASAP7_75t_L g1611 ( .A(n_1290), .Y(n_1611) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1291), .B(n_1292), .Y(n_1290) );
INVx2_ASAP7_75t_L g1340 ( .A(n_1293), .Y(n_1340) );
INVxp67_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
NOR2xp33_ASAP7_75t_L g1460 ( .A(n_1301), .B(n_1317), .Y(n_1460) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1302), .B(n_1306), .Y(n_1301) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1302), .Y(n_1331) );
OR2x2_ASAP7_75t_L g1366 ( .A(n_1302), .B(n_1325), .Y(n_1366) );
NAND2xp5_ASAP7_75t_L g1372 ( .A(n_1302), .B(n_1333), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1383 ( .A(n_1302), .B(n_1324), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1389 ( .A(n_1302), .B(n_1325), .Y(n_1389) );
NOR2xp33_ASAP7_75t_L g1471 ( .A(n_1302), .B(n_1472), .Y(n_1471) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1302), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1303), .B(n_1305), .Y(n_1302) );
OR2x2_ASAP7_75t_L g1356 ( .A(n_1306), .B(n_1330), .Y(n_1356) );
OR2x2_ASAP7_75t_L g1387 ( .A(n_1306), .B(n_1388), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_1306), .B(n_1383), .Y(n_1407) );
AOI222xp33_ASAP7_75t_L g1493 ( .A1(n_1306), .A2(n_1429), .B1(n_1435), .B2(n_1443), .C1(n_1494), .C2(n_1496), .Y(n_1493) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1308), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1333 ( .A(n_1307), .B(n_1308), .Y(n_1333) );
OAI321xp33_ASAP7_75t_L g1415 ( .A1(n_1309), .A2(n_1416), .A3(n_1419), .B1(n_1420), .B2(n_1421), .C(n_1422), .Y(n_1415) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1310), .B(n_1344), .Y(n_1379) );
NOR2xp33_ASAP7_75t_L g1449 ( .A(n_1310), .B(n_1317), .Y(n_1449) );
NOR2xp33_ASAP7_75t_L g1452 ( .A(n_1310), .B(n_1453), .Y(n_1452) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1311), .B(n_1320), .Y(n_1319) );
OR2x2_ASAP7_75t_L g1349 ( .A(n_1311), .B(n_1321), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1311), .B(n_1352), .Y(n_1367) );
OR2x2_ASAP7_75t_L g1369 ( .A(n_1311), .B(n_1362), .Y(n_1369) );
INVx2_ASAP7_75t_L g1398 ( .A(n_1311), .Y(n_1398) );
OR2x2_ASAP7_75t_L g1406 ( .A(n_1311), .B(n_1344), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1474 ( .A(n_1311), .B(n_1344), .Y(n_1474) );
INVx2_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
OR2x2_ASAP7_75t_L g1414 ( .A(n_1312), .B(n_1362), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1314), .Y(n_1312) );
NOR2xp33_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1318), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1316), .B(n_1348), .Y(n_1371) );
NAND3xp33_ASAP7_75t_L g1378 ( .A(n_1316), .B(n_1376), .C(n_1379), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1316), .B(n_1320), .Y(n_1455) );
AND2x2_ASAP7_75t_L g1496 ( .A(n_1316), .B(n_1319), .Y(n_1496) );
CKINVDCx5p33_ASAP7_75t_R g1316 ( .A(n_1317), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1317), .B(n_1320), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1409 ( .A(n_1317), .B(n_1337), .Y(n_1409) );
NAND2x1_ASAP7_75t_L g1486 ( .A(n_1317), .B(n_1487), .Y(n_1486) );
NOR2xp33_ASAP7_75t_L g1328 ( .A(n_1318), .B(n_1329), .Y(n_1328) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_1319), .B(n_1418), .Y(n_1421) );
INVx2_ASAP7_75t_L g1385 ( .A(n_1320), .Y(n_1385) );
NAND2xp5_ASAP7_75t_L g1431 ( .A(n_1320), .B(n_1352), .Y(n_1431) );
OAI31xp33_ASAP7_75t_L g1477 ( .A1(n_1320), .A2(n_1325), .A3(n_1370), .B(n_1478), .Y(n_1477) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1321), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1323), .Y(n_1321) );
NOR2xp33_ASAP7_75t_L g1375 ( .A(n_1324), .B(n_1376), .Y(n_1375) );
OR2x2_ASAP7_75t_L g1424 ( .A(n_1324), .B(n_1333), .Y(n_1424) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1324), .B(n_1333), .Y(n_1458) );
INVx2_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1330 ( .A(n_1325), .B(n_1331), .Y(n_1330) );
NAND2x1p5_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1327), .Y(n_1325) );
OR2x2_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1332), .Y(n_1329) );
NAND2xp5_ASAP7_75t_L g1381 ( .A(n_1330), .B(n_1382), .Y(n_1381) );
OR2x2_ASAP7_75t_L g1430 ( .A(n_1330), .B(n_1376), .Y(n_1430) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1330), .Y(n_1465) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1332), .Y(n_1394) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1333), .Y(n_1376) );
AND2x2_ASAP7_75t_L g1481 ( .A(n_1333), .B(n_1482), .Y(n_1481) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1333), .B(n_1389), .Y(n_1487) );
OR2x2_ASAP7_75t_L g1495 ( .A(n_1333), .B(n_1482), .Y(n_1495) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
NOR2xp33_ASAP7_75t_SL g1335 ( .A(n_1336), .B(n_1344), .Y(n_1335) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1336), .Y(n_1397) );
A2O1A1Ixp33_ASAP7_75t_L g1403 ( .A1(n_1336), .A2(n_1385), .B(n_1404), .C(n_1406), .Y(n_1403) );
NAND2xp5_ASAP7_75t_L g1484 ( .A(n_1336), .B(n_1351), .Y(n_1484) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
OAI221xp5_ASAP7_75t_L g1337 ( .A1(n_1338), .A2(n_1339), .B1(n_1340), .B2(n_1341), .C(n_1342), .Y(n_1337) );
CKINVDCx5p33_ASAP7_75t_R g1498 ( .A(n_1338), .Y(n_1498) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1344), .Y(n_1348) );
INVx3_ASAP7_75t_L g1352 ( .A(n_1344), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1345), .B(n_1346), .Y(n_1344) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1347), .Y(n_1466) );
OR2x2_ASAP7_75t_L g1347 ( .A(n_1348), .B(n_1349), .Y(n_1347) );
NAND3xp33_ASAP7_75t_L g1478 ( .A(n_1348), .B(n_1355), .C(n_1383), .Y(n_1478) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1351), .B(n_1353), .Y(n_1350) );
NAND3xp33_ASAP7_75t_L g1475 ( .A(n_1351), .B(n_1383), .C(n_1476), .Y(n_1475) );
CKINVDCx14_ASAP7_75t_R g1351 ( .A(n_1352), .Y(n_1351) );
OR2x2_ASAP7_75t_L g1405 ( .A(n_1352), .B(n_1361), .Y(n_1405) );
OR2x2_ASAP7_75t_L g1413 ( .A(n_1352), .B(n_1414), .Y(n_1413) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_1352), .B(n_1435), .Y(n_1434) );
NOR2xp33_ASAP7_75t_L g1353 ( .A(n_1354), .B(n_1356), .Y(n_1353) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
NAND3xp33_ASAP7_75t_L g1357 ( .A(n_1358), .B(n_1384), .C(n_1399), .Y(n_1357) );
AOI21xp5_ASAP7_75t_L g1358 ( .A1(n_1359), .A2(n_1367), .B(n_1368), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1360), .B(n_1363), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1360), .B(n_1392), .Y(n_1391) );
O2A1O1Ixp33_ASAP7_75t_L g1456 ( .A1(n_1360), .A2(n_1457), .B(n_1459), .C(n_1461), .Y(n_1456) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1377 ( .A(n_1361), .B(n_1367), .Y(n_1377) );
OAI22xp5_ASAP7_75t_SL g1408 ( .A1(n_1361), .A2(n_1396), .B1(n_1409), .B2(n_1410), .Y(n_1408) );
OAI221xp5_ASAP7_75t_L g1485 ( .A1(n_1361), .A2(n_1486), .B1(n_1488), .B2(n_1489), .C(n_1493), .Y(n_1485) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
AOI222xp33_ASAP7_75t_L g1479 ( .A1(n_1363), .A2(n_1379), .B1(n_1407), .B2(n_1434), .C1(n_1480), .C2(n_1481), .Y(n_1479) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
OR2x2_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1366), .Y(n_1364) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1365), .Y(n_1402) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1366), .Y(n_1393) );
OAI211xp5_ASAP7_75t_SL g1432 ( .A1(n_1366), .A2(n_1433), .B(n_1436), .C(n_1438), .Y(n_1432) );
OR2x2_ASAP7_75t_L g1440 ( .A(n_1366), .B(n_1376), .Y(n_1440) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1367), .Y(n_1461) );
OAI322xp33_ASAP7_75t_L g1368 ( .A1(n_1369), .A2(n_1370), .A3(n_1372), .B1(n_1373), .B2(n_1377), .C1(n_1378), .C2(n_1380), .Y(n_1368) );
CKINVDCx5p33_ASAP7_75t_R g1435 ( .A(n_1369), .Y(n_1435) );
CKINVDCx14_ASAP7_75t_R g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1372), .Y(n_1454) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1376), .B(n_1393), .Y(n_1411) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1376), .B(n_1383), .Y(n_1418) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
NAND2xp5_ASAP7_75t_L g1442 ( .A(n_1383), .B(n_1402), .Y(n_1442) );
A2O1A1Ixp33_ASAP7_75t_R g1384 ( .A1(n_1385), .A2(n_1386), .B(n_1390), .C(n_1395), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1436 ( .A(n_1385), .B(n_1437), .Y(n_1436) );
OR2x2_ASAP7_75t_L g1450 ( .A(n_1385), .B(n_1406), .Y(n_1450) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1385), .Y(n_1488) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
AOI21xp33_ASAP7_75t_SL g1427 ( .A1(n_1387), .A2(n_1428), .B(n_1431), .Y(n_1427) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
NAND2xp5_ASAP7_75t_L g1401 ( .A(n_1389), .B(n_1402), .Y(n_1401) );
AOI211xp5_ASAP7_75t_L g1467 ( .A1(n_1389), .A2(n_1468), .B(n_1469), .C(n_1477), .Y(n_1467) );
AND2x2_ASAP7_75t_L g1492 ( .A(n_1389), .B(n_1394), .Y(n_1492) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
AND2x2_ASAP7_75t_L g1392 ( .A(n_1393), .B(n_1394), .Y(n_1392) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
NAND2xp5_ASAP7_75t_L g1396 ( .A(n_1397), .B(n_1398), .Y(n_1396) );
INVx2_ASAP7_75t_L g1420 ( .A(n_1397), .Y(n_1420) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1398), .Y(n_1480) );
AOI222xp33_ASAP7_75t_L g1399 ( .A1(n_1400), .A2(n_1403), .B1(n_1407), .B2(n_1408), .C1(n_1411), .C2(n_1412), .Y(n_1399) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
OAI21xp5_ASAP7_75t_L g1422 ( .A1(n_1407), .A2(n_1423), .B(n_1425), .Y(n_1422) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1407), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1437 ( .A(n_1410), .B(n_1411), .Y(n_1437) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1411), .Y(n_1446) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
CKINVDCx5p33_ASAP7_75t_R g1443 ( .A(n_1414), .Y(n_1443) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
AOI22xp5_ASAP7_75t_L g1462 ( .A1(n_1419), .A2(n_1463), .B1(n_1483), .B2(n_1485), .Y(n_1462) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
OAI31xp33_ASAP7_75t_L g1426 ( .A1(n_1420), .A2(n_1427), .A3(n_1432), .B(n_1444), .Y(n_1426) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
OAI221xp5_ASAP7_75t_L g1444 ( .A1(n_1430), .A2(n_1445), .B1(n_1448), .B2(n_1450), .C(n_1451), .Y(n_1444) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
OAI21xp33_ASAP7_75t_L g1438 ( .A1(n_1439), .A2(n_1441), .B(n_1443), .Y(n_1438) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
NAND2xp5_ASAP7_75t_L g1490 ( .A(n_1440), .B(n_1491), .Y(n_1490) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1446), .B(n_1447), .Y(n_1445) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1450), .Y(n_1468) );
NOR2xp33_ASAP7_75t_L g1451 ( .A(n_1452), .B(n_1456), .Y(n_1451) );
NAND2xp5_ASAP7_75t_L g1453 ( .A(n_1454), .B(n_1455), .Y(n_1453) );
CKINVDCx14_ASAP7_75t_R g1457 ( .A(n_1458), .Y(n_1457) );
INVxp67_ASAP7_75t_SL g1459 ( .A(n_1460), .Y(n_1459) );
NAND2xp5_ASAP7_75t_L g1464 ( .A(n_1465), .B(n_1466), .Y(n_1464) );
OAI21xp33_ASAP7_75t_L g1469 ( .A1(n_1470), .A2(n_1473), .B(n_1475), .Y(n_1469) );
INVxp33_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
INVxp67_ASAP7_75t_SL g1489 ( .A(n_1490), .Y(n_1489) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
CKINVDCx20_ASAP7_75t_R g1497 ( .A(n_1498), .Y(n_1497) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
AND3x1_ASAP7_75t_L g1502 ( .A(n_1503), .B(n_1530), .C(n_1541), .Y(n_1502) );
NOR2xp33_ASAP7_75t_L g1503 ( .A(n_1504), .B(n_1519), .Y(n_1503) );
OAI22xp5_ASAP7_75t_L g1524 ( .A1(n_1510), .A2(n_1514), .B1(n_1525), .B2(n_1526), .Y(n_1524) );
INVx2_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
INVx2_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
AOI22xp33_ASAP7_75t_SL g1535 ( .A1(n_1536), .A2(n_1537), .B1(n_1538), .B2(n_1539), .Y(n_1535) );
AOI22xp33_ASAP7_75t_L g1548 ( .A1(n_1537), .A2(n_1549), .B1(n_1550), .B2(n_1552), .Y(n_1548) );
INVx2_ASAP7_75t_L g1546 ( .A(n_1547), .Y(n_1546) );
INVx2_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
INVx1_ASAP7_75t_L g1556 ( .A(n_1557), .Y(n_1556) );
BUFx3_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
INVxp33_ASAP7_75t_SL g1562 ( .A(n_1563), .Y(n_1562) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1566), .Y(n_1565) );
NAND3xp33_ASAP7_75t_L g1566 ( .A(n_1567), .B(n_1578), .C(n_1585), .Y(n_1566) );
AND4x1_ASAP7_75t_L g1585 ( .A(n_1586), .B(n_1593), .C(n_1597), .D(n_1601), .Y(n_1585) );
NAND3xp33_ASAP7_75t_L g1586 ( .A(n_1587), .B(n_1590), .C(n_1591), .Y(n_1586) );
INVx2_ASAP7_75t_SL g1591 ( .A(n_1592), .Y(n_1591) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
BUFx3_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
OAI21xp5_ASAP7_75t_L g1609 ( .A1(n_1610), .A2(n_1611), .B(n_1612), .Y(n_1609) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
endmodule