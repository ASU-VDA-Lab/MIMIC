module fake_ibex_643_n_961 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_188, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_961);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_188;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_961;

wire n_599;
wire n_822;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_510;
wire n_193;
wire n_845;
wire n_947;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_708;
wire n_280;
wire n_375;
wire n_340;
wire n_317;
wire n_698;
wire n_901;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_276;
wire n_470;
wire n_339;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_857;
wire n_849;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_560;
wire n_429;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_648;
wire n_571;
wire n_472;
wire n_209;
wire n_229;
wire n_589;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_433;
wire n_299;
wire n_439;
wire n_262;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_567;
wire n_516;
wire n_548;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_200;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_397;
wire n_366;
wire n_283;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_379;
wire n_288;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_385;
wire n_233;
wire n_414;
wire n_342;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_450;
wire n_302;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_890;
wire n_912;
wire n_921;
wire n_816;
wire n_874;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

NOR2xp67_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_86),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_39),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_61),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_52),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_29),
.Y(n_197)
);

INVxp33_ASAP7_75t_SL g198 ( 
.A(n_184),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_22),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_51),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_38),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_63),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_91),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_102),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_100),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_11),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_29),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_82),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_0),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_16),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_154),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_158),
.Y(n_216)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_147),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_92),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_104),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_108),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_143),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_70),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_95),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_39),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_121),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_38),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_157),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

NOR2xp67_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_72),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_176),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_25),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_46),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_77),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_133),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_11),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_27),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_54),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_96),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_113),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_181),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_32),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_27),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_187),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_156),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_162),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_4),
.B(n_137),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_106),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_75),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_139),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_166),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_87),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_128),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_99),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_85),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_98),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_57),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_81),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_141),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_14),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_76),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_21),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_111),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_191),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_136),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_71),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_49),
.B(n_90),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_118),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_84),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_172),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_18),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_182),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_140),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_129),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_5),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_23),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_30),
.Y(n_277)
);

INVxp33_ASAP7_75t_SL g278 ( 
.A(n_168),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_97),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_171),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_135),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_12),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_125),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_10),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_74),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_174),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_149),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_53),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_130),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_89),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_83),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_66),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_186),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_192),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_25),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_124),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_80),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_188),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_101),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_179),
.B(n_109),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g301 ( 
.A(n_132),
.B(n_22),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_47),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_60),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_117),
.B(n_19),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_68),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_48),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_43),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_94),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_20),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_64),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_146),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_33),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_126),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_148),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_119),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_3),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_73),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_16),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_4),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_112),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_161),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_203),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_281),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_282),
.B(n_1),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_282),
.B(n_2),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_226),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_209),
.B(n_3),
.Y(n_327)
);

OA21x2_ASAP7_75t_L g328 ( 
.A1(n_201),
.A2(n_78),
.B(n_189),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_226),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_217),
.B(n_6),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_269),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_217),
.B(n_6),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_269),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_269),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_269),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_204),
.B(n_7),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_221),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_208),
.B(n_8),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_195),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_212),
.B(n_8),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_221),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_196),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_257),
.B(n_9),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_202),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_303),
.B(n_9),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_205),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_223),
.B(n_10),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_221),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_206),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_199),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_245),
.B(n_13),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_221),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_199),
.A2(n_319),
.B1(n_266),
.B2(n_280),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_207),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_210),
.Y(n_356)
);

OAI22x1_ASAP7_75t_R g357 ( 
.A1(n_247),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_215),
.Y(n_358)
);

AND2x6_ASAP7_75t_L g359 ( 
.A(n_256),
.B(n_45),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_235),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_239),
.B(n_15),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_285),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_218),
.B(n_50),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_281),
.B(n_17),
.Y(n_364)
);

NOR2x1_ASAP7_75t_L g365 ( 
.A(n_301),
.B(n_19),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_247),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_259),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_219),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_216),
.B(n_24),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_297),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_251),
.B(n_24),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_225),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_285),
.B(n_26),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_305),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_297),
.B(n_26),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_218),
.B(n_55),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_227),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_305),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_201),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_228),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_214),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_284),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_222),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_230),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_266),
.Y(n_385)
);

OA21x2_ASAP7_75t_L g386 ( 
.A1(n_222),
.A2(n_103),
.B(n_183),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_280),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_240),
.B(n_28),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_289),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_289),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_233),
.Y(n_391)
);

OA21x2_ASAP7_75t_L g392 ( 
.A1(n_253),
.A2(n_107),
.B(n_178),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_194),
.B(n_34),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_388),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_323),
.B(n_264),
.Y(n_395)
);

BUFx4f_ASAP7_75t_L g396 ( 
.A(n_346),
.Y(n_396)
);

INVx6_ASAP7_75t_L g397 ( 
.A(n_371),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_L g398 ( 
.A1(n_388),
.A2(n_213),
.B1(n_318),
.B2(n_316),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_388),
.A2(n_211),
.B1(n_197),
.B2(n_224),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_323),
.B(n_315),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_323),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_340),
.B(n_272),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_323),
.B(n_198),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_388),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_362),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_324),
.Y(n_406)
);

BUFx10_ASAP7_75t_L g407 ( 
.A(n_346),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_324),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_374),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_340),
.B(n_272),
.Y(n_410)
);

NAND3xp33_ASAP7_75t_L g411 ( 
.A(n_343),
.B(n_237),
.C(n_234),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_324),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g413 ( 
.A(n_373),
.B(n_293),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_SL g414 ( 
.A1(n_351),
.A2(n_290),
.B1(n_320),
.B2(n_231),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_333),
.B(n_198),
.Y(n_415)
);

NAND3xp33_ASAP7_75t_L g416 ( 
.A(n_343),
.B(n_243),
.C(n_238),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_345),
.B(n_293),
.Y(n_417)
);

OR2x6_ASAP7_75t_L g418 ( 
.A(n_322),
.B(n_236),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_324),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_333),
.B(n_278),
.Y(n_420)
);

NOR2x1p5_ASAP7_75t_L g421 ( 
.A(n_333),
.B(n_241),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_331),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_330),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_354),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_325),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_331),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_325),
.Y(n_427)
);

OR2x6_ASAP7_75t_L g428 ( 
.A(n_322),
.B(n_242),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_345),
.A2(n_276),
.B1(n_261),
.B2(n_309),
.Y(n_429)
);

OR2x6_ASAP7_75t_L g430 ( 
.A(n_389),
.B(n_271),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_333),
.B(n_370),
.Y(n_431)
);

AO22x2_ASAP7_75t_L g432 ( 
.A1(n_325),
.A2(n_304),
.B1(n_277),
.B2(n_275),
.Y(n_432)
);

INVx5_ASAP7_75t_L g433 ( 
.A(n_359),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_347),
.A2(n_312),
.B1(n_278),
.B2(n_214),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_347),
.B(n_321),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_359),
.B(n_290),
.Y(n_436)
);

INVx6_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_338),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_334),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_371),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_330),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_332),
.A2(n_320),
.B1(n_220),
.B2(n_260),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_367),
.B(n_260),
.Y(n_443)
);

AND3x1_ASAP7_75t_L g444 ( 
.A(n_366),
.B(n_246),
.C(n_254),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_373),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_370),
.B(n_200),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_382),
.B(n_307),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_335),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_332),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_350),
.B(n_321),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_373),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g453 ( 
.A(n_373),
.B(n_255),
.Y(n_453)
);

NAND3xp33_ASAP7_75t_L g454 ( 
.A(n_350),
.B(n_298),
.C(n_314),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_378),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_359),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_355),
.B(n_263),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_355),
.B(n_265),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_360),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_337),
.B(n_214),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_346),
.A2(n_246),
.B1(n_214),
.B2(n_295),
.Y(n_462)
);

OR2x6_ASAP7_75t_L g463 ( 
.A(n_389),
.B(n_295),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_356),
.B(n_268),
.Y(n_464)
);

INVxp33_ASAP7_75t_L g465 ( 
.A(n_354),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_336),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_336),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_385),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_356),
.A2(n_295),
.B1(n_313),
.B2(n_311),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_337),
.B(n_341),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_378),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_393),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_359),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_379),
.Y(n_474)
);

BUFx6f_ASAP7_75t_SL g475 ( 
.A(n_359),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_358),
.B(n_273),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_359),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_358),
.B(n_274),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_368),
.B(n_279),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_364),
.B(n_286),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_383),
.Y(n_482)
);

AND2x6_ASAP7_75t_L g483 ( 
.A(n_364),
.B(n_288),
.Y(n_483)
);

OR2x6_ASAP7_75t_L g484 ( 
.A(n_375),
.B(n_348),
.Y(n_484)
);

OR2x6_ASAP7_75t_L g485 ( 
.A(n_375),
.B(n_295),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_348),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_372),
.B(n_292),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_372),
.B(n_294),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_328),
.Y(n_489)
);

AO21x2_ASAP7_75t_L g490 ( 
.A1(n_369),
.A2(n_300),
.B(n_310),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_423),
.B(n_341),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_423),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_450),
.B(n_361),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_461),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_456),
.B(n_377),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_422),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_485),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_403),
.B(n_380),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_460),
.B(n_387),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_443),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_426),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_432),
.A2(n_380),
.B1(n_384),
.B2(n_391),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_474),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_432),
.A2(n_384),
.B1(n_391),
.B2(n_361),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_485),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_481),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_473),
.B(n_363),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_415),
.B(n_420),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_470),
.B(n_339),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_441),
.B(n_344),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_486),
.B(n_327),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_485),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_468),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_449),
.B(n_352),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_439),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_482),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_395),
.B(n_326),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_394),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_484),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_448),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_404),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_473),
.B(n_376),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_477),
.B(n_433),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_421),
.B(n_365),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_480),
.A2(n_366),
.B1(n_390),
.B2(n_365),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_445),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_400),
.B(n_326),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_431),
.B(n_329),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_480),
.B(n_329),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_440),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_480),
.B(n_232),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_477),
.B(n_296),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_466),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_467),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_483),
.B(n_244),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_445),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_483),
.B(n_249),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_458),
.B(n_302),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_486),
.B(n_351),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_413),
.B(n_250),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_413),
.B(n_252),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_472),
.B(n_306),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_447),
.B(n_390),
.Y(n_543)
);

A2O1A1Ixp33_ASAP7_75t_L g544 ( 
.A1(n_396),
.A2(n_193),
.B(n_229),
.C(n_267),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_413),
.B(n_258),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g546 ( 
.A(n_436),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_397),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_401),
.B(n_270),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_433),
.B(n_248),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_437),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_433),
.B(n_248),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_433),
.B(n_248),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_484),
.A2(n_317),
.B1(n_308),
.B2(n_283),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_455),
.B(n_287),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_446),
.B(n_299),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_471),
.B(n_291),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_442),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_396),
.B(n_453),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_453),
.B(n_328),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_490),
.B(n_328),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_436),
.B(n_248),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_490),
.B(n_386),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_405),
.Y(n_563)
);

OAI22xp33_ASAP7_75t_L g564 ( 
.A1(n_465),
.A2(n_357),
.B1(n_386),
.B2(n_392),
.Y(n_564)
);

A2O1A1Ixp33_ASAP7_75t_L g565 ( 
.A1(n_406),
.A2(n_267),
.B(n_381),
.C(n_262),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_398),
.B(n_386),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_414),
.B(n_386),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_489),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_407),
.B(n_392),
.Y(n_569)
);

AND2x6_ASAP7_75t_SL g570 ( 
.A(n_430),
.B(n_357),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_398),
.A2(n_381),
.B1(n_392),
.B2(n_262),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_399),
.B(n_392),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_452),
.B(n_262),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_408),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_424),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_444),
.A2(n_381),
.B1(n_262),
.B2(n_349),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_452),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_511),
.B(n_434),
.Y(n_578)
);

BUFx12f_ASAP7_75t_L g579 ( 
.A(n_570),
.Y(n_579)
);

A2O1A1Ixp33_ASAP7_75t_L g580 ( 
.A1(n_498),
.A2(n_427),
.B(n_425),
.C(n_419),
.Y(n_580)
);

O2A1O1Ixp33_ASAP7_75t_L g581 ( 
.A1(n_509),
.A2(n_514),
.B(n_492),
.C(n_491),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_560),
.A2(n_412),
.B(n_479),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_498),
.B(n_434),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_557),
.A2(n_444),
.B1(n_463),
.B2(n_418),
.Y(n_584)
);

AOI221xp5_ASAP7_75t_L g585 ( 
.A1(n_543),
.A2(n_414),
.B1(n_429),
.B2(n_488),
.C(n_464),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_504),
.A2(n_462),
.B1(n_463),
.B2(n_429),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_502),
.A2(n_463),
.B1(n_469),
.B2(n_428),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_510),
.B(n_459),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_568),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_569),
.A2(n_478),
.B(n_459),
.Y(n_590)
);

A2O1A1Ixp33_ASAP7_75t_L g591 ( 
.A1(n_508),
.A2(n_487),
.B(n_476),
.C(n_457),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_494),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_500),
.B(n_418),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_519),
.B(n_430),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_499),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_493),
.B(n_402),
.Y(n_596)
);

AOI33xp33_ASAP7_75t_L g597 ( 
.A1(n_539),
.A2(n_409),
.A3(n_402),
.B1(n_451),
.B2(n_410),
.B3(n_435),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_510),
.B(n_410),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_536),
.B(n_411),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_546),
.A2(n_475),
.B1(n_454),
.B2(n_416),
.Y(n_600)
);

BUFx12f_ASAP7_75t_L g601 ( 
.A(n_513),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_512),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_497),
.Y(n_603)
);

O2A1O1Ixp33_ASAP7_75t_SL g604 ( 
.A1(n_565),
.A2(n_451),
.B(n_435),
.C(n_417),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_525),
.B(n_417),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_569),
.A2(n_416),
.B(n_438),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_497),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_553),
.B(n_34),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_524),
.B(n_35),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_558),
.A2(n_338),
.B1(n_342),
.B2(n_349),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_575),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_505),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_566),
.A2(n_572),
.B1(n_574),
.B2(n_576),
.Y(n_613)
);

AOI21x1_ASAP7_75t_L g614 ( 
.A1(n_571),
.A2(n_353),
.B(n_349),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_538),
.B(n_542),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_567),
.A2(n_353),
.B1(n_349),
.B2(n_342),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_563),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_495),
.A2(n_353),
.B(n_349),
.Y(n_618)
);

INVx8_ASAP7_75t_L g619 ( 
.A(n_526),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_530),
.B(n_36),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_550),
.B(n_36),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_518),
.B(n_37),
.Y(n_622)
);

A2O1A1Ixp33_ASAP7_75t_L g623 ( 
.A1(n_521),
.A2(n_37),
.B(n_40),
.C(n_41),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_503),
.B(n_40),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_577),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_550),
.B(n_41),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_532),
.A2(n_114),
.B(n_175),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_506),
.B(n_42),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_529),
.Y(n_629)
);

AOI21xp33_ASAP7_75t_L g630 ( 
.A1(n_531),
.A2(n_42),
.B(n_43),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_517),
.B(n_44),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_555),
.B(n_44),
.Y(n_632)
);

O2A1O1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_544),
.A2(n_56),
.B(n_58),
.C(n_59),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_527),
.B(n_190),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_523),
.A2(n_62),
.B(n_65),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_523),
.A2(n_67),
.B(n_69),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_496),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_528),
.A2(n_79),
.B1(n_88),
.B2(n_93),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_507),
.A2(n_522),
.B(n_573),
.Y(n_639)
);

CKINVDCx8_ASAP7_75t_R g640 ( 
.A(n_535),
.Y(n_640)
);

BUFx4f_ASAP7_75t_L g641 ( 
.A(n_516),
.Y(n_641)
);

O2A1O1Ixp33_ASAP7_75t_L g642 ( 
.A1(n_547),
.A2(n_105),
.B(n_110),
.C(n_115),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_522),
.A2(n_573),
.B(n_561),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_537),
.B(n_116),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_501),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_645)
);

AO21x1_ASAP7_75t_L g646 ( 
.A1(n_549),
.A2(n_127),
.B(n_131),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_515),
.A2(n_134),
.B1(n_138),
.B2(n_142),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_SL g648 ( 
.A1(n_540),
.A2(n_144),
.B1(n_145),
.B2(n_150),
.Y(n_648)
);

A2O1A1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_520),
.A2(n_151),
.B(n_152),
.C(n_155),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_612),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_601),
.Y(n_651)
);

OAI21x1_ASAP7_75t_L g652 ( 
.A1(n_639),
.A2(n_551),
.B(n_552),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_590),
.A2(n_548),
.B(n_541),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_612),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_592),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_596),
.B(n_533),
.Y(n_656)
);

AND2x2_ASAP7_75t_SL g657 ( 
.A(n_641),
.B(n_545),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_595),
.B(n_556),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_584),
.B(n_534),
.Y(n_659)
);

AO21x2_ASAP7_75t_L g660 ( 
.A1(n_616),
.A2(n_533),
.B(n_554),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_582),
.A2(n_159),
.B(n_163),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_620),
.Y(n_662)
);

OAI22x1_ASAP7_75t_L g663 ( 
.A1(n_608),
.A2(n_173),
.B1(n_169),
.B2(n_170),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_643),
.A2(n_606),
.B(n_581),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_612),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_587),
.A2(n_586),
.B1(n_585),
.B2(n_605),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_619),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_593),
.B(n_594),
.Y(n_668)
);

INVx3_ASAP7_75t_SL g669 ( 
.A(n_617),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_607),
.B(n_602),
.Y(n_670)
);

A2O1A1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_615),
.A2(n_597),
.B(n_632),
.C(n_591),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_583),
.A2(n_578),
.B1(n_631),
.B2(n_580),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_622),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_604),
.A2(n_599),
.B(n_600),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_634),
.A2(n_618),
.B(n_625),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_602),
.Y(n_676)
);

BUFx12f_ASAP7_75t_L g677 ( 
.A(n_579),
.Y(n_677)
);

NAND2x1p5_ASAP7_75t_L g678 ( 
.A(n_603),
.B(n_641),
.Y(n_678)
);

O2A1O1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_623),
.A2(n_630),
.B(n_609),
.C(n_624),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_628),
.A2(n_633),
.B(n_644),
.C(n_642),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_SL g681 ( 
.A1(n_603),
.A2(n_621),
.B(n_626),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_611),
.Y(n_682)
);

AOI221x1_ASAP7_75t_L g683 ( 
.A1(n_638),
.A2(n_648),
.B1(n_649),
.B2(n_647),
.C(n_610),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_629),
.A2(n_637),
.B1(n_640),
.B2(n_589),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_589),
.Y(n_685)
);

AOI211x1_ASAP7_75t_L g686 ( 
.A1(n_646),
.A2(n_627),
.B(n_635),
.C(n_636),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_645),
.B(n_598),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_617),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_595),
.B(n_499),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_592),
.Y(n_690)
);

AO21x1_ASAP7_75t_L g691 ( 
.A1(n_633),
.A2(n_564),
.B(n_613),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_617),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_588),
.A2(n_598),
.B1(n_586),
.B2(n_504),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_639),
.A2(n_559),
.B(n_560),
.Y(n_694)
);

AO31x2_ASAP7_75t_L g695 ( 
.A1(n_613),
.A2(n_571),
.A3(n_560),
.B(n_562),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_589),
.Y(n_696)
);

NOR2xp67_ASAP7_75t_L g697 ( 
.A(n_612),
.B(n_598),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_639),
.A2(n_559),
.B(n_560),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_639),
.A2(n_559),
.B(n_560),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_595),
.B(n_497),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_595),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_612),
.Y(n_702)
);

BUFx12f_ASAP7_75t_L g703 ( 
.A(n_601),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_598),
.B(n_588),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_595),
.B(n_557),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_SL g706 ( 
.A(n_587),
.B(n_247),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_595),
.B(n_497),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_598),
.B(n_588),
.Y(n_708)
);

A2O1A1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_581),
.A2(n_590),
.B(n_508),
.C(n_498),
.Y(n_709)
);

O2A1O1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_581),
.A2(n_615),
.B(n_591),
.C(n_508),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_617),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_SL g712 ( 
.A(n_587),
.B(n_456),
.Y(n_712)
);

AO31x2_ASAP7_75t_L g713 ( 
.A1(n_613),
.A2(n_571),
.A3(n_560),
.B(n_562),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_639),
.A2(n_559),
.B(n_560),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_598),
.B(n_588),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_639),
.A2(n_559),
.B(n_560),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_617),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_598),
.B(n_588),
.Y(n_718)
);

AOI31xp67_ASAP7_75t_L g719 ( 
.A1(n_616),
.A2(n_562),
.A3(n_560),
.B(n_561),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_612),
.B(n_592),
.Y(n_720)
);

AO31x2_ASAP7_75t_L g721 ( 
.A1(n_613),
.A2(n_571),
.A3(n_560),
.B(n_562),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_592),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_598),
.B(n_588),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_595),
.B(n_557),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_639),
.A2(n_559),
.B(n_560),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_592),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_595),
.B(n_557),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_639),
.A2(n_559),
.B(n_560),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_595),
.Y(n_729)
);

AO31x2_ASAP7_75t_L g730 ( 
.A1(n_613),
.A2(n_571),
.A3(n_560),
.B(n_562),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_596),
.B(n_484),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_639),
.A2(n_559),
.B(n_560),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_588),
.A2(n_598),
.B1(n_586),
.B2(n_504),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_587),
.A2(n_586),
.B1(n_585),
.B2(n_584),
.Y(n_734)
);

OAI22x1_ASAP7_75t_L g735 ( 
.A1(n_595),
.A2(n_387),
.B1(n_385),
.B2(n_366),
.Y(n_735)
);

A2O1A1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_581),
.A2(n_590),
.B(n_508),
.C(n_498),
.Y(n_736)
);

AO21x2_ASAP7_75t_L g737 ( 
.A1(n_614),
.A2(n_616),
.B(n_604),
.Y(n_737)
);

O2A1O1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_581),
.A2(n_615),
.B(n_591),
.C(n_508),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_588),
.A2(n_598),
.B1(n_586),
.B2(n_504),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_598),
.B(n_588),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_598),
.B(n_588),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_592),
.Y(n_742)
);

INVx4_ASAP7_75t_SL g743 ( 
.A(n_579),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_595),
.B(n_557),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_639),
.A2(n_559),
.B(n_560),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_639),
.A2(n_559),
.B(n_560),
.Y(n_746)
);

CKINVDCx11_ASAP7_75t_R g747 ( 
.A(n_703),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_690),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_722),
.Y(n_749)
);

A2O1A1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_710),
.A2(n_738),
.B(n_666),
.C(n_734),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_704),
.B(n_708),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_726),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_669),
.Y(n_753)
);

OAI21x1_ASAP7_75t_SL g754 ( 
.A1(n_734),
.A2(n_661),
.B(n_702),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_715),
.B(n_718),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_723),
.B(n_740),
.Y(n_756)
);

AO21x2_ASAP7_75t_L g757 ( 
.A1(n_674),
.A2(n_691),
.B(n_737),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_741),
.Y(n_758)
);

OAI22xp33_ASAP7_75t_SL g759 ( 
.A1(n_676),
.A2(n_689),
.B1(n_678),
.B2(n_701),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_742),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_731),
.B(n_656),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_668),
.B(n_659),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_697),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_666),
.B(n_709),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_697),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_692),
.Y(n_766)
);

OAI21xp5_ASAP7_75t_L g767 ( 
.A1(n_736),
.A2(n_671),
.B(n_687),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_729),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_693),
.B(n_733),
.Y(n_769)
);

OR2x6_ASAP7_75t_L g770 ( 
.A(n_667),
.B(n_688),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_706),
.A2(n_724),
.B1(n_744),
.B2(n_705),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_727),
.B(n_670),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_739),
.B(n_658),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_720),
.B(n_735),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_662),
.B(n_673),
.Y(n_775)
);

OAI21xp5_ASAP7_75t_L g776 ( 
.A1(n_679),
.A2(n_653),
.B(n_680),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_681),
.A2(n_684),
.B1(n_665),
.B2(n_650),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_657),
.B(n_700),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_707),
.B(n_665),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_654),
.B(n_696),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_694),
.A2(n_746),
.B(n_745),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_698),
.A2(n_725),
.B(n_716),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_685),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_663),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_682),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_711),
.Y(n_786)
);

AO21x2_ASAP7_75t_L g787 ( 
.A1(n_660),
.A2(n_732),
.B(n_714),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_717),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_652),
.Y(n_789)
);

AO31x2_ASAP7_75t_L g790 ( 
.A1(n_683),
.A2(n_699),
.A3(n_728),
.B(n_675),
.Y(n_790)
);

OA21x2_ASAP7_75t_L g791 ( 
.A1(n_719),
.A2(n_713),
.B(n_730),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_651),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_695),
.Y(n_793)
);

OAI21x1_ASAP7_75t_L g794 ( 
.A1(n_686),
.A2(n_695),
.B(n_713),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_721),
.B(n_743),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_743),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_677),
.B(n_704),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_655),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_704),
.B(n_708),
.Y(n_799)
);

AND2x2_ASAP7_75t_SL g800 ( 
.A(n_666),
.B(n_712),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_669),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_655),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_704),
.B(n_708),
.Y(n_803)
);

AO31x2_ASAP7_75t_L g804 ( 
.A1(n_691),
.A2(n_664),
.A3(n_672),
.B(n_674),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_655),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_655),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_704),
.B(n_708),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_702),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_704),
.B(n_708),
.Y(n_809)
);

NAND2x1p5_ASAP7_75t_L g810 ( 
.A(n_667),
.B(n_612),
.Y(n_810)
);

AO21x2_ASAP7_75t_L g811 ( 
.A1(n_674),
.A2(n_691),
.B(n_737),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_704),
.B(n_708),
.Y(n_812)
);

AO21x1_ASAP7_75t_L g813 ( 
.A1(n_706),
.A2(n_564),
.B(n_734),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_667),
.Y(n_814)
);

OR2x6_ASAP7_75t_L g815 ( 
.A(n_754),
.B(n_795),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_758),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_803),
.B(n_809),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_758),
.Y(n_818)
);

AO21x2_ASAP7_75t_L g819 ( 
.A1(n_776),
.A2(n_782),
.B(n_781),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_751),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_755),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_756),
.B(n_799),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_807),
.B(n_756),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_812),
.B(n_762),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_793),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_771),
.B(n_775),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_813),
.A2(n_800),
.B1(n_764),
.B2(n_773),
.Y(n_827)
);

INVx1_ASAP7_75t_SL g828 ( 
.A(n_753),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_768),
.Y(n_829)
);

OR2x6_ASAP7_75t_L g830 ( 
.A(n_795),
.B(n_784),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_748),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_749),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_752),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_769),
.B(n_750),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_814),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_760),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_798),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_802),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_766),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_805),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_769),
.B(n_806),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_777),
.B(n_814),
.Y(n_842)
);

OR2x6_ASAP7_75t_L g843 ( 
.A(n_814),
.B(n_808),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_800),
.B(n_761),
.Y(n_844)
);

BUFx12f_ASAP7_75t_L g845 ( 
.A(n_747),
.Y(n_845)
);

AO21x2_ASAP7_75t_L g846 ( 
.A1(n_794),
.A2(n_767),
.B(n_757),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_810),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_810),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_772),
.B(n_797),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_789),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_804),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_770),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_770),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_804),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_834),
.B(n_804),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_834),
.B(n_791),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_850),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_842),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_823),
.B(n_811),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_819),
.B(n_811),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_842),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_843),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_842),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_825),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_820),
.B(n_757),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_843),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_819),
.B(n_787),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_841),
.B(n_790),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_815),
.B(n_787),
.Y(n_869)
);

NAND2x1_ASAP7_75t_L g870 ( 
.A(n_842),
.B(n_783),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_842),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_815),
.B(n_780),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_SL g873 ( 
.A1(n_844),
.A2(n_759),
.B1(n_774),
.B2(n_801),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_827),
.B(n_763),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_868),
.B(n_821),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_864),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_862),
.Y(n_877)
);

INVx4_ASAP7_75t_L g878 ( 
.A(n_862),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_859),
.B(n_854),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_859),
.B(n_851),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_856),
.B(n_854),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_856),
.B(n_846),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_865),
.B(n_830),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_857),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_867),
.B(n_846),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_869),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_884),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_882),
.B(n_855),
.Y(n_888)
);

OAI31xp33_ASAP7_75t_L g889 ( 
.A1(n_877),
.A2(n_835),
.A3(n_817),
.B(n_852),
.Y(n_889)
);

OR2x2_ASAP7_75t_L g890 ( 
.A(n_875),
.B(n_865),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_876),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_882),
.B(n_867),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_875),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_884),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_885),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_882),
.B(n_867),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_881),
.B(n_860),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_877),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_881),
.B(n_860),
.Y(n_899)
);

AND2x4_ASAP7_75t_SL g900 ( 
.A(n_878),
.B(n_872),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_880),
.A2(n_871),
.B1(n_861),
.B2(n_863),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_877),
.A2(n_835),
.B(n_873),
.C(n_870),
.Y(n_902)
);

OAI21xp33_ASAP7_75t_L g903 ( 
.A1(n_895),
.A2(n_873),
.B(n_885),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_891),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_887),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_893),
.B(n_880),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_890),
.B(n_879),
.Y(n_907)
);

OAI32xp33_ASAP7_75t_L g908 ( 
.A1(n_895),
.A2(n_878),
.A3(n_828),
.B1(n_886),
.B2(n_883),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_887),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_894),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_892),
.B(n_885),
.Y(n_911)
);

AO22x1_ASAP7_75t_L g912 ( 
.A1(n_898),
.A2(n_878),
.B1(n_862),
.B2(n_866),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_890),
.B(n_879),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_888),
.B(n_839),
.Y(n_914)
);

NAND4xp25_ASAP7_75t_SL g915 ( 
.A(n_906),
.B(n_902),
.C(n_889),
.D(n_901),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_903),
.A2(n_888),
.B1(n_896),
.B2(n_892),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_904),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_904),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_905),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_914),
.B(n_845),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_909),
.Y(n_921)
);

AOI21xp33_ASAP7_75t_L g922 ( 
.A1(n_914),
.A2(n_849),
.B(n_818),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_907),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_913),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_910),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_911),
.A2(n_896),
.B1(n_897),
.B2(n_899),
.Y(n_926)
);

OAI221xp5_ASAP7_75t_L g927 ( 
.A1(n_916),
.A2(n_889),
.B1(n_898),
.B2(n_858),
.C(n_863),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_925),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_917),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_915),
.A2(n_912),
.B(n_908),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_919),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_921),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_930),
.A2(n_927),
.B1(n_920),
.B2(n_929),
.Y(n_933)
);

NOR3x1_ASAP7_75t_L g934 ( 
.A(n_931),
.B(n_786),
.C(n_796),
.Y(n_934)
);

AOI221x1_ASAP7_75t_L g935 ( 
.A1(n_932),
.A2(n_918),
.B1(n_922),
.B2(n_924),
.C(n_923),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_933),
.B(n_926),
.Y(n_936)
);

NOR3xp33_ASAP7_75t_L g937 ( 
.A(n_935),
.B(n_747),
.C(n_785),
.Y(n_937)
);

NOR4xp25_ASAP7_75t_SL g938 ( 
.A(n_937),
.B(n_845),
.C(n_922),
.D(n_934),
.Y(n_938)
);

NOR3xp33_ASAP7_75t_L g939 ( 
.A(n_936),
.B(n_788),
.C(n_765),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_939),
.B(n_928),
.Y(n_940)
);

NOR3xp33_ASAP7_75t_SL g941 ( 
.A(n_938),
.B(n_792),
.C(n_826),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_940),
.Y(n_942)
);

AOI22x1_ASAP7_75t_L g943 ( 
.A1(n_941),
.A2(n_792),
.B1(n_853),
.B2(n_816),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_942),
.B(n_943),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_942),
.B(n_928),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_943),
.A2(n_770),
.B1(n_874),
.B2(n_900),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_944),
.A2(n_942),
.B(n_945),
.Y(n_947)
);

OAI22x1_ASAP7_75t_L g948 ( 
.A1(n_946),
.A2(n_829),
.B1(n_847),
.B2(n_848),
.Y(n_948)
);

OAI22xp33_ASAP7_75t_L g949 ( 
.A1(n_944),
.A2(n_843),
.B1(n_874),
.B2(n_822),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_944),
.A2(n_778),
.B(n_824),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_947),
.B(n_910),
.Y(n_951)
);

NAND2x1p5_ASAP7_75t_L g952 ( 
.A(n_950),
.B(n_948),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_949),
.A2(n_817),
.B1(n_843),
.B2(n_900),
.Y(n_953)
);

AOI21xp33_ASAP7_75t_L g954 ( 
.A1(n_947),
.A2(n_779),
.B(n_840),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_947),
.A2(n_843),
.B(n_831),
.Y(n_955)
);

OAI31xp33_ASAP7_75t_SL g956 ( 
.A1(n_953),
.A2(n_836),
.A3(n_833),
.B(n_832),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_951),
.A2(n_866),
.B1(n_838),
.B2(n_837),
.Y(n_957)
);

NAND3xp33_ASAP7_75t_L g958 ( 
.A(n_955),
.B(n_838),
.C(n_837),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_957),
.B(n_952),
.Y(n_959)
);

OA21x2_ASAP7_75t_L g960 ( 
.A1(n_958),
.A2(n_954),
.B(n_832),
.Y(n_960)
);

AOI21xp33_ASAP7_75t_L g961 ( 
.A1(n_959),
.A2(n_960),
.B(n_956),
.Y(n_961)
);


endmodule