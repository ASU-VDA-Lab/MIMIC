module fake_jpeg_3597_n_197 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_197);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_1),
.B(n_23),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_20),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_11),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_12),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_80),
.Y(n_84)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_80),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_49),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_56),
.B1(n_66),
.B2(n_54),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_94),
.B1(n_62),
.B2(n_50),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_66),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_90),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_49),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_91),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_58),
.B1(n_57),
.B2(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_95),
.B(n_63),
.Y(n_102)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_97),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_91),
.A2(n_76),
.B(n_71),
.C(n_67),
.Y(n_98)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_98),
.A2(n_9),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_103),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_58),
.B1(n_55),
.B2(n_50),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_107),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_84),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_106),
.B1(n_108),
.B2(n_5),
.Y(n_128)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_51),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_61),
.B1(n_69),
.B2(n_5),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_4),
.Y(n_124)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_112),
.Y(n_117)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_96),
.B(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_18),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_2),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_119),
.B(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_122),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_89),
.Y(n_122)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_4),
.Y(n_127)
);

NAND2xp33_ASAP7_75t_R g150 ( 
.A(n_128),
.B(n_135),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_100),
.B(n_6),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_133),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_134),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_7),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_98),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_15),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_142),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_113),
.C(n_97),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_132),
.C(n_112),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_16),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_16),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_143),
.B(n_146),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_154),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_21),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_22),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_152),
.Y(n_158)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_25),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_26),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_157),
.Y(n_159)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_156),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_28),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_162),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_137),
.A2(n_30),
.B(n_32),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_161),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_47),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_145),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_163)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_145),
.A3(n_152),
.B1(n_155),
.B2(n_151),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_167),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_148),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_37),
.B(n_39),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_41),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_179),
.B(n_181),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_164),
.Y(n_177)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_166),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_167),
.C(n_160),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_163),
.C(n_173),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_138),
.B1(n_170),
.B2(n_171),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_138),
.B1(n_159),
.B2(n_172),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_182),
.B(n_158),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_189),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_178),
.B(n_162),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_190),
.B(n_174),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_192),
.B(n_184),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_185),
.C(n_191),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_140),
.B(n_43),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_136),
.Y(n_197)
);


endmodule