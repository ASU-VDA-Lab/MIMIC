module fake_jpeg_322_n_467 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_467);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_467;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_48),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_50),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_23),
.B(n_16),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_62),
.Y(n_103)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_55),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_15),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_43),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_65),
.B(n_66),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_34),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_72),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_77),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_92),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_91),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_94),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_47),
.A2(n_40),
.B1(n_26),
.B2(n_45),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_98),
.A2(n_108),
.B1(n_150),
.B2(n_34),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_49),
.A2(n_26),
.B1(n_41),
.B2(n_38),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_101),
.A2(n_94),
.B1(n_93),
.B2(n_88),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_55),
.A2(n_28),
.B1(n_41),
.B2(n_38),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_104),
.A2(n_114),
.B1(n_122),
.B2(n_146),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_26),
.B1(n_41),
.B2(n_38),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_66),
.C(n_20),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_109),
.B(n_34),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_50),
.A2(n_28),
.B1(n_41),
.B2(n_18),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_56),
.B(n_27),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_130),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_69),
.A2(n_28),
.B1(n_18),
.B2(n_46),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_64),
.B(n_27),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_77),
.B(n_43),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_132),
.B(n_151),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_87),
.A2(n_46),
.B1(n_24),
.B2(n_39),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_L g150 ( 
.A1(n_78),
.A2(n_42),
.B1(n_39),
.B2(n_20),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_92),
.B(n_29),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_152),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_153),
.Y(n_225)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_154),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_155),
.Y(n_239)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_159),
.Y(n_217)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_160),
.Y(n_229)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_161),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_162),
.A2(n_188),
.B1(n_192),
.B2(n_193),
.Y(n_228)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_163),
.Y(n_234)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_165),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_166),
.B(n_178),
.Y(n_226)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_171),
.Y(n_210)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_169),
.Y(n_238)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_172),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_173),
.B(n_176),
.Y(n_218)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_174),
.Y(n_241)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_177),
.Y(n_219)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_95),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_117),
.A2(n_73),
.B1(n_76),
.B2(n_91),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_179),
.A2(n_142),
.B1(n_140),
.B2(n_105),
.Y(n_221)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_107),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_180),
.B(n_181),
.Y(n_223)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_182),
.B(n_183),
.Y(n_240)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_95),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_184),
.A2(n_86),
.B1(n_144),
.B2(n_120),
.Y(n_220)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_185),
.B(n_186),
.Y(n_247)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_124),
.Y(n_186)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_137),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_99),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_201),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_120),
.Y(n_190)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_103),
.B(n_112),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_191),
.B(n_195),
.Y(n_237)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_135),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_134),
.B(n_24),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_194),
.B(n_196),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_34),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_123),
.B(n_29),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_110),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_135),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_148),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_102),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_203),
.B(n_205),
.Y(n_249)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_102),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_144),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_105),
.B(n_22),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_99),
.B(n_34),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_206),
.A2(n_113),
.B1(n_35),
.B2(n_42),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_197),
.A2(n_104),
.B1(n_114),
.B2(n_146),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_208),
.A2(n_220),
.B1(n_221),
.B2(n_227),
.Y(n_268)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_209),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_164),
.B(n_122),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_216),
.B(n_222),
.C(n_236),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_142),
.C(n_140),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_174),
.B(n_22),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_248),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_184),
.A2(n_35),
.B1(n_42),
.B2(n_113),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_242),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_176),
.B(n_136),
.C(n_42),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_177),
.B1(n_181),
.B2(n_200),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_167),
.B(n_0),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_185),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_250),
.A2(n_251),
.B1(n_1),
.B2(n_3),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_198),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_211),
.B(n_172),
.Y(n_254)
);

NAND3xp33_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_259),
.C(n_274),
.Y(n_293)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_215),
.Y(n_255)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_255),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_155),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_257),
.B(n_258),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_157),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_210),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_169),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_263),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_183),
.C(n_178),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_261),
.B(n_235),
.C(n_244),
.Y(n_302)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_215),
.Y(n_262)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_262),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_170),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_264),
.Y(n_325)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_217),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_265),
.Y(n_303)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_266),
.B(n_270),
.Y(n_307)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_272),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_208),
.A2(n_179),
.B1(n_197),
.B2(n_190),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_269),
.A2(n_279),
.B1(n_1),
.B2(n_7),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_225),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_229),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_273),
.B(n_275),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_211),
.B(n_189),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_223),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_276),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_192),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_277),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_218),
.B(n_165),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_280),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_218),
.A2(n_207),
.B1(n_221),
.B2(n_209),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_152),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_241),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_281),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_207),
.A2(n_193),
.B(n_136),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_282),
.A2(n_285),
.B(n_289),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_283),
.A2(n_284),
.B1(n_287),
.B2(n_291),
.Y(n_311)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_245),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_241),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_224),
.B(n_219),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_288),
.Y(n_300)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_225),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_240),
.B(n_1),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_239),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_228),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_213),
.B1(n_245),
.B2(n_214),
.Y(n_295)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_230),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g294 ( 
.A(n_256),
.B(n_236),
.CI(n_233),
.CON(n_294),
.SN(n_294)
);

OA21x2_ASAP7_75t_SL g354 ( 
.A1(n_294),
.A2(n_267),
.B(n_291),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_295),
.B(n_310),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_269),
.A2(n_232),
.B1(n_213),
.B2(n_214),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_298),
.A2(n_305),
.B1(n_309),
.B2(n_316),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_302),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_268),
.A2(n_230),
.B1(n_234),
.B2(n_244),
.Y(n_305)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_256),
.B(n_234),
.C(n_239),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_306),
.B(n_284),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_268),
.A2(n_238),
.B1(n_235),
.B2(n_212),
.Y(n_309)
);

OAI32xp33_ASAP7_75t_L g310 ( 
.A1(n_260),
.A2(n_238),
.A3(n_212),
.B1(n_231),
.B2(n_243),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_278),
.A2(n_231),
.B(n_243),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_312),
.A2(n_313),
.B(n_315),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_279),
.A2(n_13),
.B(n_5),
.Y(n_313)
);

OAI32xp33_ASAP7_75t_L g314 ( 
.A1(n_253),
.A2(n_13),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_290),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_263),
.A2(n_1),
.B(n_6),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_282),
.A2(n_7),
.B(n_8),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_318),
.A2(n_321),
.B(n_264),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_253),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_319),
.A2(n_322),
.B1(n_255),
.B2(n_262),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_271),
.A2(n_9),
.B(n_10),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_271),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_261),
.B(n_12),
.C(n_275),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_324),
.B(n_315),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_300),
.B(n_252),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_327),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_299),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_328),
.B(n_331),
.Y(n_358)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_299),
.Y(n_330)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_330),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_299),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_297),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_335),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_308),
.A2(n_276),
.B(n_286),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_333),
.A2(n_349),
.B(n_350),
.Y(n_360)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_297),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_317),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_336),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_337),
.B(n_354),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_316),
.A2(n_252),
.B1(n_280),
.B2(n_285),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_338),
.A2(n_305),
.B1(n_309),
.B2(n_296),
.Y(n_361)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_317),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_342),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_301),
.B(n_288),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_340),
.B(n_341),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_326),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_344),
.A2(n_353),
.B1(n_355),
.B2(n_283),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_301),
.B(n_287),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_346),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_307),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_347),
.Y(n_368)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_304),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_348),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_308),
.A2(n_265),
.B(n_272),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_293),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_351),
.A2(n_352),
.B(n_313),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_312),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_325),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_325),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_356),
.B(n_292),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_361),
.B(n_329),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_354),
.B(n_306),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_362),
.B(n_365),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_292),
.C(n_296),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_364),
.B(n_367),
.C(n_369),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_334),
.A2(n_298),
.B1(n_320),
.B2(n_294),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_366),
.A2(n_378),
.B1(n_362),
.B2(n_363),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_356),
.B(n_302),
.C(n_294),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_300),
.C(n_324),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_330),
.B(n_303),
.C(n_323),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_372),
.B(n_373),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_303),
.C(n_323),
.Y(n_373)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_374),
.Y(n_386)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_377),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_310),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_378),
.B(n_380),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_314),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_334),
.B(n_295),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_329),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_383),
.A2(n_384),
.B1(n_391),
.B2(n_395),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_358),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_385),
.B(n_397),
.Y(n_419)
);

BUFx24_ASAP7_75t_SL g388 ( 
.A(n_368),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_388),
.B(n_399),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_382),
.A2(n_352),
.B1(n_331),
.B2(n_328),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_372),
.Y(n_392)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_392),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_361),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_376),
.B(n_340),
.Y(n_394)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_394),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_375),
.A2(n_338),
.B1(n_344),
.B2(n_341),
.Y(n_395)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_375),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_370),
.Y(n_398)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_398),
.Y(n_417)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_359),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_379),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_401),
.B(n_347),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_360),
.A2(n_343),
.B(n_349),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_402),
.A2(n_360),
.B(n_380),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_343),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_403),
.B(n_375),
.Y(n_414)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_404),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_384),
.B(n_363),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_405),
.B(n_410),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_406),
.A2(n_402),
.B(n_391),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_367),
.C(n_373),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_408),
.B(n_409),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_396),
.B(n_369),
.C(n_366),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_389),
.B(n_365),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_414),
.C(n_400),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_395),
.A2(n_374),
.B1(n_371),
.B2(n_381),
.Y(n_415)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_415),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_386),
.A2(n_357),
.B1(n_344),
.B2(n_346),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_418),
.A2(n_393),
.B1(n_311),
.B2(n_387),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_389),
.B(n_332),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_387),
.C(n_353),
.Y(n_432)
);

BUFx24_ASAP7_75t_SL g422 ( 
.A(n_412),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_422),
.B(n_432),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_428),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_407),
.B(n_351),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_424),
.B(n_426),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_396),
.C(n_400),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_416),
.A2(n_383),
.B1(n_390),
.B2(n_397),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_429),
.A2(n_414),
.B(n_420),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_411),
.B(n_403),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_430),
.Y(n_440)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_431),
.Y(n_435)
);

OAI321xp33_ASAP7_75t_L g434 ( 
.A1(n_427),
.A2(n_419),
.A3(n_417),
.B1(n_418),
.B2(n_406),
.C(n_339),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_434),
.B(n_335),
.Y(n_445)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_421),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_436),
.B(n_437),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_428),
.A2(n_410),
.B1(n_405),
.B2(n_311),
.Y(n_437)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_432),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_441),
.B(n_444),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_443),
.B(n_437),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_336),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_445),
.B(n_448),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_446),
.B(n_435),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_426),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_442),
.B(n_433),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_449),
.B(n_450),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_439),
.B(n_423),
.C(n_409),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_440),
.B(n_444),
.Y(n_452)
);

NOR3xp33_ASAP7_75t_SL g457 ( 
.A(n_452),
.B(n_355),
.C(n_443),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_453),
.B(n_455),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_451),
.B(n_439),
.Y(n_455)
);

AO21x1_ASAP7_75t_L g460 ( 
.A1(n_457),
.A2(n_447),
.B(n_321),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_456),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_459),
.A2(n_460),
.B(n_446),
.Y(n_462)
);

MAJx2_ASAP7_75t_L g461 ( 
.A(n_458),
.B(n_454),
.C(n_450),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_461),
.A2(n_462),
.B(n_413),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_463),
.A2(n_318),
.B(n_342),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_464),
.A2(n_322),
.B(n_319),
.Y(n_465)
);

NOR3xp33_ASAP7_75t_SL g466 ( 
.A(n_465),
.B(n_266),
.C(n_273),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_466),
.B(n_281),
.Y(n_467)
);


endmodule