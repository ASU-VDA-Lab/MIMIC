module fake_jpeg_3180_n_89 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_89);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_89;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_22),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_23),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_35),
.Y(n_48)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_25),
.C(n_31),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_2),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_32),
.B1(n_35),
.B2(n_29),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_46),
.B1(n_3),
.B2(n_4),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_13),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_56),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_36),
.B1(n_27),
.B2(n_38),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_53),
.B1(n_47),
.B2(n_6),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_55),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_3),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_47),
.B(n_7),
.Y(n_62)
);

BUFx24_ASAP7_75t_SL g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_18),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_65),
.B1(n_17),
.B2(n_19),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_15),
.Y(n_75)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_64),
.B(n_67),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_11),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_14),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVxp33_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_75),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_77),
.C(n_65),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_74),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_82),
.A2(n_81),
.B1(n_73),
.B2(n_75),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_83),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_80),
.B(n_78),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_69),
.B1(n_71),
.B2(n_62),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_20),
.C(n_21),
.Y(n_89)
);


endmodule