module real_jpeg_20409_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_0),
.A2(n_8),
.B1(n_23),
.B2(n_24),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_0),
.A2(n_23),
.B1(n_31),
.B2(n_37),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_1),
.A2(n_8),
.B1(n_24),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_1),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_3),
.B(n_35),
.Y(n_34)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_3),
.A2(n_34),
.B(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_3),
.B(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_3),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_3),
.A2(n_8),
.B(n_12),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_3),
.A2(n_31),
.B1(n_37),
.B2(n_99),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_3),
.A2(n_27),
.B1(n_109),
.B2(n_110),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_3),
.B(n_63),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_4),
.A2(n_31),
.B1(n_37),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_4),
.A2(n_32),
.B1(n_35),
.B2(n_54),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_4),
.A2(n_8),
.B1(n_24),
.B2(n_54),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_5),
.A2(n_32),
.B1(n_35),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_5),
.A2(n_31),
.B1(n_37),
.B2(n_46),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_5),
.A2(n_8),
.B1(n_24),
.B2(n_46),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_24),
.Y(n_25)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_7),
.A2(n_31),
.B1(n_37),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_7),
.A2(n_8),
.B1(n_24),
.B2(n_56),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_8),
.A2(n_9),
.B1(n_24),
.B2(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_8),
.A2(n_12),
.B1(n_24),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_11),
.A2(n_32),
.B1(n_35),
.B2(n_70),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_12),
.A2(n_31),
.B(n_50),
.C(n_51),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_12),
.B(n_31),
.Y(n_50)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_86),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_85),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_57),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_18),
.B(n_57),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_39),
.C(n_47),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_19),
.A2(n_20),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_21),
.B(n_30),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_25),
.B(n_26),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_22),
.B(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_24),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_25),
.B(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_25),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_25),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_27),
.B(n_99),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_28),
.Y(n_77)
);

AOI32xp33_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.A3(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_30)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_43)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_38),
.B(n_42),
.C(n_43),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_38),
.Y(n_42)
);

NAND2xp33_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_37),
.A2(n_52),
.B(n_99),
.C(n_100),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_39),
.A2(n_40),
.B1(n_47),
.B2(n_48),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_55),
.B(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_49),
.A2(n_51),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_49),
.A2(n_51),
.B1(n_53),
.B2(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_51),
.B(n_99),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_78),
.B2(n_79),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_66),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_75),
.B(n_76),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_75),
.A2(n_92),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

XOR2x2_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_129),
.B(n_134),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_117),
.B(n_128),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_105),
.B(n_116),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_96),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_96),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_110),
.B(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_102),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_101),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_111),
.B(n_115),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_108),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_118),
.B(n_119),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_125),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_124),
.C(n_125),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_131),
.Y(n_134)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);


endmodule