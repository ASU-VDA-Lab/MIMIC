module fake_jpeg_2084_n_485 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_485);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_485;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_48),
.B(n_53),
.Y(n_112)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_19),
.B(n_14),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx5_ASAP7_75t_SL g145 ( 
.A(n_61),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_15),
.B(n_14),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_68),
.B(n_90),
.Y(n_134)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_88),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_89),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_15),
.B(n_13),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_93),
.Y(n_140)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_96),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_94),
.B(n_95),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_40),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_36),
.B1(n_41),
.B2(n_42),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_99),
.A2(n_127),
.B1(n_132),
.B2(n_95),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_53),
.A2(n_38),
.B(n_25),
.C(n_42),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_102),
.B(n_21),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_106),
.A2(n_46),
.B1(n_45),
.B2(n_61),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_57),
.A2(n_26),
.B1(n_25),
.B2(n_39),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_117),
.A2(n_125),
.B1(n_147),
.B2(n_153),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_62),
.A2(n_26),
.B1(n_25),
.B2(n_39),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_36),
.B1(n_41),
.B2(n_44),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_89),
.A2(n_40),
.B1(n_20),
.B2(n_44),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_137),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_50),
.B(n_30),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_141),
.B(n_151),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_62),
.A2(n_26),
.B1(n_20),
.B2(n_44),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g149 ( 
.A1(n_54),
.A2(n_30),
.B1(n_20),
.B2(n_21),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_32),
.B1(n_24),
.B2(n_45),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_50),
.B(n_32),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_52),
.A2(n_30),
.B1(n_21),
.B2(n_24),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_83),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_157),
.A2(n_188),
.B(n_193),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_166),
.Y(n_205)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_105),
.Y(n_162)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_163),
.A2(n_110),
.B1(n_101),
.B2(n_138),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_168),
.Y(n_214)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_102),
.B(n_32),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_111),
.A2(n_45),
.B1(n_46),
.B2(n_24),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_175),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_206)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_183),
.Y(n_209)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_106),
.B(n_46),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_199),
.Y(n_201)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_121),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_103),
.B(n_75),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_186),
.Y(n_218)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_142),
.A2(n_94),
.B1(n_93),
.B2(n_90),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_187),
.A2(n_113),
.B1(n_138),
.B2(n_130),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_103),
.B(n_13),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_145),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_190),
.B(n_194),
.Y(n_226)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_98),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_135),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_104),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_108),
.Y(n_229)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_104),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_136),
.A2(n_82),
.B1(n_80),
.B2(n_77),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_198),
.A2(n_100),
.B1(n_101),
.B2(n_110),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_139),
.B(n_74),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_204),
.A2(n_207),
.B1(n_222),
.B2(n_230),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_164),
.A2(n_143),
.B1(n_150),
.B2(n_65),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_182),
.A2(n_149),
.B1(n_123),
.B2(n_148),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_215),
.A2(n_231),
.B1(n_170),
.B2(n_169),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_165),
.B(n_107),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_193),
.C(n_126),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_157),
.A2(n_173),
.B1(n_163),
.B2(n_158),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_109),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_225),
.Y(n_239)
);

OAI32xp33_ASAP7_75t_L g225 ( 
.A1(n_161),
.A2(n_109),
.A3(n_120),
.B1(n_152),
.B2(n_145),
.Y(n_225)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_198),
.B(n_120),
.CI(n_126),
.CON(n_227),
.SN(n_227)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_227),
.B(n_144),
.Y(n_260)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_235),
.Y(n_266)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_237),
.Y(n_294)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_200),
.A2(n_172),
.B(n_174),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_240),
.A2(n_241),
.B(n_249),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_218),
.A2(n_206),
.B(n_200),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_197),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_242),
.B(n_243),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_191),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_192),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_257),
.C(n_262),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_195),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_247),
.Y(n_281)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_246),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_201),
.B(n_224),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_218),
.A2(n_179),
.B(n_186),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_250),
.B(n_244),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_209),
.A2(n_201),
.B1(n_230),
.B2(n_227),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_251),
.A2(n_259),
.B1(n_227),
.B2(n_226),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_209),
.A2(n_133),
.B1(n_113),
.B2(n_130),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_252),
.A2(n_213),
.B1(n_196),
.B2(n_176),
.Y(n_287)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_133),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_254),
.Y(n_285)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_255),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_207),
.B(n_156),
.C(n_189),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_202),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_260),
.B(n_203),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_205),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_264),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_162),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_209),
.A2(n_204),
.B1(n_212),
.B2(n_211),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_205),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_265),
.A2(n_273),
.B1(n_293),
.B2(n_257),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_254),
.A2(n_227),
.B1(n_223),
.B2(n_219),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_267),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_251),
.A2(n_239),
.B1(n_256),
.B2(n_254),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_272),
.A2(n_278),
.B1(n_291),
.B2(n_252),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_256),
.A2(n_220),
.B1(n_223),
.B2(n_219),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_274),
.B(n_290),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_239),
.A2(n_220),
.B1(n_234),
.B2(n_232),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_264),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_292),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_234),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_282),
.B(n_255),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_244),
.B(n_232),
.C(n_233),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_250),
.C(n_253),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_259),
.B1(n_235),
.B2(n_237),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_289),
.B(n_148),
.Y(n_324)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_240),
.B(n_213),
.CI(n_202),
.CON(n_290),
.SN(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_254),
.A2(n_233),
.B1(n_208),
.B2(n_228),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_245),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_263),
.A2(n_171),
.B1(n_178),
.B2(n_180),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_295),
.A2(n_303),
.B1(n_308),
.B2(n_291),
.Y(n_325)
);

OAI32xp33_ASAP7_75t_L g296 ( 
.A1(n_272),
.A2(n_260),
.A3(n_257),
.B1(n_236),
.B2(n_243),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_296),
.A2(n_297),
.B(n_294),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_277),
.A2(n_241),
.B(n_285),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_277),
.A2(n_249),
.B(n_248),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_298),
.A2(n_311),
.B(n_290),
.Y(n_331)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_268),
.Y(n_299)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_288),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_300),
.B(n_321),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_302),
.A2(n_320),
.B1(n_273),
.B2(n_293),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_278),
.A2(n_262),
.B1(n_250),
.B2(n_249),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_304),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_275),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_305),
.A2(n_309),
.B1(n_316),
.B2(n_323),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_262),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_314),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_310),
.C(n_324),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_288),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_261),
.C(n_242),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_276),
.A2(n_235),
.B(n_238),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_268),
.Y(n_312)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_312),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_258),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_271),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_283),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_317),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_282),
.B(n_208),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_266),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_269),
.B(n_235),
.Y(n_319)
);

NAND3xp33_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_322),
.C(n_274),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_265),
.A2(n_255),
.B1(n_246),
.B2(n_228),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_269),
.B(n_184),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_144),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_325),
.B(n_353),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_326),
.A2(n_333),
.B1(n_348),
.B2(n_349),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_281),
.C(n_285),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_329),
.B(n_351),
.C(n_355),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_347),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_331),
.A2(n_317),
.B(n_115),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_321),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_332),
.B(n_342),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_320),
.A2(n_281),
.B1(n_290),
.B2(n_287),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_267),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_334),
.B(n_337),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_307),
.B(n_324),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_271),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_339),
.B(n_343),
.Y(n_372)
);

FAx1_ASAP7_75t_SL g340 ( 
.A(n_297),
.B(n_290),
.CI(n_284),
.CON(n_340),
.SN(n_340)
);

MAJx2_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_344),
.C(n_346),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_301),
.B(n_284),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_303),
.B(n_296),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_323),
.B(n_283),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_315),
.A2(n_270),
.B1(n_266),
.B2(n_294),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_295),
.A2(n_302),
.B1(n_309),
.B2(n_315),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_SL g350 ( 
.A(n_298),
.B(n_270),
.C(n_246),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_352),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_123),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_313),
.B(n_111),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_311),
.A2(n_63),
.B1(n_67),
.B2(n_66),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_305),
.B(n_108),
.C(n_60),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_336),
.Y(n_357)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_335),
.Y(n_358)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_358),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_345),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_361),
.B(n_366),
.Y(n_401)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_354),
.Y(n_362)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_362),
.Y(n_391)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_341),
.Y(n_364)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_364),
.Y(n_394)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_338),
.Y(n_365)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_365),
.Y(n_404)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_346),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_331),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_367),
.B(n_373),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_349),
.A2(n_313),
.B1(n_316),
.B2(n_312),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_369),
.A2(n_326),
.B1(n_343),
.B2(n_340),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_327),
.B(n_328),
.C(n_337),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_55),
.C(n_16),
.Y(n_396)
);

INVxp33_ASAP7_75t_SL g373 ( 
.A(n_347),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_374),
.B(n_376),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_344),
.A2(n_299),
.B(n_304),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_375),
.A2(n_377),
.B(n_355),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_348),
.Y(n_376)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_380),
.B(n_381),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_329),
.B(n_317),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_339),
.B(n_12),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_382),
.B(n_0),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_384),
.A2(n_385),
.B1(n_376),
.B2(n_377),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_363),
.A2(n_340),
.B1(n_334),
.B2(n_328),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_386),
.B(n_378),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_327),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_388),
.B(n_397),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_368),
.B(n_351),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_395),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_368),
.B(n_115),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_396),
.B(n_364),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_360),
.B(n_16),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_360),
.B(n_43),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_398),
.B(n_399),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_372),
.B(n_371),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_374),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_400),
.A2(n_362),
.B1(n_358),
.B2(n_380),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_0),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_402),
.B(n_403),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_375),
.B(n_10),
.C(n_1),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_0),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_383),
.Y(n_406)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_406),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_388),
.B(n_366),
.C(n_371),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_410),
.B(n_413),
.Y(n_437)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_412),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_389),
.B(n_367),
.C(n_365),
.Y(n_413)
);

BUFx24_ASAP7_75t_SL g414 ( 
.A(n_387),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_414),
.B(n_417),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_363),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_415),
.B(n_418),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_416),
.B(n_419),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_385),
.A2(n_356),
.B(n_357),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_393),
.B(n_359),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_401),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_420),
.B(n_421),
.Y(n_426)
);

BUFx24_ASAP7_75t_SL g421 ( 
.A(n_390),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_392),
.A2(n_361),
.B(n_369),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_422),
.A2(n_424),
.B1(n_425),
.B2(n_1),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_423),
.B(n_386),
.C(n_402),
.Y(n_428)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_430),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_412),
.A2(n_404),
.B(n_384),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_429),
.A2(n_433),
.B(n_442),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_418),
.A2(n_379),
.B1(n_400),
.B2(n_394),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_415),
.B(n_398),
.C(n_397),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_431),
.B(n_434),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_413),
.A2(n_379),
.B(n_395),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_408),
.B(n_396),
.C(n_405),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_425),
.A2(n_406),
.B1(n_407),
.B2(n_411),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_436),
.B(n_438),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_1),
.C(n_2),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_4),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_410),
.A2(n_1),
.B(n_3),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_R g443 ( 
.A(n_441),
.B(n_409),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_443),
.A2(n_452),
.B1(n_445),
.B2(n_426),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_432),
.B(n_411),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_445),
.Y(n_461)
);

OR2x6_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_3),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_437),
.A2(n_9),
.B(n_4),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_448),
.A2(n_6),
.B(n_7),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_436),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_450),
.B(n_453),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_440),
.B(n_3),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_451),
.B(n_455),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_435),
.B(n_4),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_4),
.Y(n_454)
);

NOR2xp67_ASAP7_75t_L g459 ( 
.A(n_454),
.B(n_438),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_5),
.C(n_6),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_456),
.B(n_5),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_447),
.A2(n_433),
.B(n_427),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_457),
.A2(n_460),
.B(n_6),
.Y(n_473)
);

AOI21x1_ASAP7_75t_L g469 ( 
.A1(n_458),
.A2(n_445),
.B(n_455),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_459),
.B(n_462),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_449),
.A2(n_442),
.B(n_430),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_434),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_465),
.B(n_466),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_456),
.B(n_431),
.C(n_426),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_467),
.Y(n_470)
);

O2A1O1Ixp33_ASAP7_75t_SL g475 ( 
.A1(n_469),
.A2(n_457),
.B(n_466),
.C(n_463),
.Y(n_475)
);

NOR2x1p5_ASAP7_75t_L g471 ( 
.A(n_462),
.B(n_445),
.Y(n_471)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_471),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_461),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_472),
.B(n_473),
.Y(n_478)
);

OAI21xp33_ASAP7_75t_L g480 ( 
.A1(n_475),
.A2(n_476),
.B(n_470),
.Y(n_480)
);

O2A1O1Ixp33_ASAP7_75t_SL g476 ( 
.A1(n_468),
.A2(n_464),
.B(n_8),
.C(n_9),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_478),
.B(n_474),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_479),
.B(n_480),
.C(n_481),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_477),
.A2(n_9),
.B(n_7),
.Y(n_481)
);

AO21x2_ASAP7_75t_L g483 ( 
.A1(n_482),
.A2(n_9),
.B(n_7),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_483),
.A2(n_7),
.B(n_8),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_484),
.Y(n_485)
);


endmodule