module fake_jpeg_10442_n_284 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NOR3xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_0),
.C(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_38),
.Y(n_49)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_30),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_45),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_26),
.B1(n_21),
.B2(n_23),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_39),
.B1(n_37),
.B2(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_17),
.B1(n_29),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_60),
.B1(n_57),
.B2(n_45),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_40),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

CKINVDCx9p33_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_61),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_20),
.B1(n_27),
.B2(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_30),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_70),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_76),
.B1(n_59),
.B2(n_46),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_37),
.B1(n_27),
.B2(n_20),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_43),
.B(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_69),
.B(n_15),
.Y(n_101)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_34),
.B1(n_37),
.B2(n_22),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_71),
.A2(n_75),
.B1(n_59),
.B2(n_46),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_37),
.B1(n_35),
.B2(n_22),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_41),
.B1(n_26),
.B2(n_28),
.Y(n_75)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_42),
.A2(n_25),
.A3(n_41),
.B1(n_26),
.B2(n_18),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_77),
.A2(n_53),
.B(n_52),
.C(n_28),
.Y(n_109)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_79),
.Y(n_107)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_83),
.Y(n_111)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_84),
.B(n_41),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_28),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_62),
.B(n_61),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_109),
.B(n_97),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_91),
.A2(n_97),
.B1(n_4),
.B2(n_5),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_101),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_64),
.A2(n_82),
.B1(n_72),
.B2(n_88),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_60),
.B(n_54),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_106),
.B(n_79),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_81),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_73),
.C(n_66),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_67),
.B1(n_89),
.B2(n_87),
.Y(n_118)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_104),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_66),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_108),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_70),
.A2(n_52),
.B(n_59),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_109),
.A2(n_89),
.B1(n_50),
.B2(n_58),
.Y(n_132)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_65),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_63),
.B(n_53),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_83),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_78),
.B(n_15),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_114),
.B(n_13),
.Y(n_126)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_117),
.B(n_119),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_91),
.B1(n_108),
.B2(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_120),
.B(n_124),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_136),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_122),
.B(n_123),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_67),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_128),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_114),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_131),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_141),
.B1(n_92),
.B2(n_93),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_3),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_133),
.A2(n_134),
.B(n_101),
.Y(n_167)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_65),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_3),
.Y(n_137)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_112),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_143),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_4),
.Y(n_142)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_144),
.B(n_152),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_145),
.A2(n_151),
.B1(n_156),
.B2(n_162),
.Y(n_192)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_98),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_160),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_109),
.Y(n_149)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_143),
.A2(n_102),
.B1(n_115),
.B2(n_103),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_121),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_110),
.Y(n_155)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

AO21x1_ASAP7_75t_SL g156 ( 
.A1(n_139),
.A2(n_115),
.B(n_6),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_5),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_138),
.B1(n_118),
.B2(n_141),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_170),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_167),
.B(n_133),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_6),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

AO21x1_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_6),
.B(n_7),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_169),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_142),
.Y(n_170)
);

AND2x6_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_8),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_128),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_182),
.C(n_183),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_155),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_177),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_150),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_146),
.B(n_165),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_178),
.A2(n_151),
.B(n_167),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_156),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_179),
.A2(n_169),
.B(n_172),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_153),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_125),
.C(n_140),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_133),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_125),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_195),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_147),
.B(n_136),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_197),
.Y(n_202)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_186),
.B(n_129),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_199),
.B(n_206),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_204),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_178),
.B(n_129),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_187),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_213),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_193),
.A2(n_191),
.B1(n_181),
.B2(n_144),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_209),
.A2(n_216),
.B1(n_218),
.B2(n_180),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_162),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_212),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_196),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_184),
.A2(n_160),
.B(n_171),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_214),
.B(n_217),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_182),
.A2(n_117),
.B(n_119),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_215),
.B(n_219),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_154),
.B1(n_145),
.B2(n_130),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_174),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_222),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_183),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_227),
.C(n_231),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_177),
.C(n_187),
.Y(n_227)
);

FAx1_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_175),
.CI(n_158),
.CON(n_229),
.SN(n_229)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_230),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_126),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_9),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_9),
.C(n_10),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_201),
.C(n_213),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_229),
.B(n_204),
.Y(n_239)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_198),
.Y(n_240)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g241 ( 
.A(n_229),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_242),
.Y(n_252)
);

INVxp67_ASAP7_75t_SL g242 ( 
.A(n_232),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_246),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_244),
.B(n_249),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_245),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_208),
.B1(n_202),
.B2(n_216),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_248),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_205),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_247),
.B(n_233),
.Y(n_250)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_250),
.Y(n_261)
);

OAI21x1_ASAP7_75t_SL g254 ( 
.A1(n_245),
.A2(n_209),
.B(n_203),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_9),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_233),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_258),
.B(n_230),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_227),
.C(n_220),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_258),
.Y(n_265)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_257),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_262),
.B(n_264),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_256),
.A2(n_225),
.B1(n_247),
.B2(n_238),
.Y(n_263)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_260),
.C(n_250),
.Y(n_271)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_253),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_266),
.A2(n_259),
.B(n_252),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_207),
.B1(n_235),
.B2(n_11),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_267),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_268),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_269),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_10),
.C(n_11),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_SL g275 ( 
.A1(n_274),
.A2(n_268),
.B(n_261),
.C(n_267),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_278),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_273),
.A2(n_255),
.B(n_11),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_272),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_280),
.B(n_276),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_281),
.A2(n_279),
.B(n_270),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_10),
.B(n_12),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_12),
.Y(n_284)
);


endmodule