module fake_jpeg_18063_n_248 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_38),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_22),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_28),
.B1(n_25),
.B2(n_18),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_45),
.A2(n_47),
.B1(n_57),
.B2(n_24),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_25),
.B1(n_18),
.B2(n_19),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_37),
.B1(n_41),
.B2(n_44),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_48),
.A2(n_19),
.B1(n_42),
.B2(n_36),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_53),
.B(n_62),
.Y(n_65)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_18),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_40),
.B(n_36),
.C(n_39),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_19),
.B1(n_23),
.B2(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_21),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_32),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_32),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_66),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_79),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_55),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_75),
.B(n_45),
.Y(n_108)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_40),
.C(n_36),
.Y(n_72)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_17),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_76),
.B(n_84),
.Y(n_100)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_81),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_40),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_49),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_42),
.B1(n_36),
.B2(n_22),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_85),
.B1(n_94),
.B2(n_61),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_17),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_57),
.B(n_31),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_49),
.Y(n_91)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_30),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_92),
.B(n_30),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_101),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_92),
.B1(n_93),
.B2(n_77),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_110),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_108),
.A2(n_111),
.B(n_115),
.Y(n_121)
);

AOI32xp33_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_51),
.A3(n_59),
.B1(n_58),
.B2(n_42),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_67),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_56),
.Y(n_111)
);

AOI22x1_ASAP7_75t_L g112 ( 
.A1(n_70),
.A2(n_48),
.B1(n_56),
.B2(n_58),
.Y(n_112)
);

OAI22x1_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_75),
.B1(n_83),
.B2(n_74),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_59),
.B1(n_24),
.B2(n_21),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_33),
.B1(n_59),
.B2(n_73),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_0),
.Y(n_115)
);

OR2x2_ASAP7_75t_SL g116 ( 
.A(n_67),
.B(n_26),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_68),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_133),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_119),
.B(n_110),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_124),
.B(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_100),
.B(n_65),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_131),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_129),
.A2(n_141),
.B1(n_144),
.B2(n_115),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_93),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_136),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_95),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_132),
.B(n_137),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_145),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_86),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_90),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_26),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_105),
.B(n_33),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_146),
.Y(n_151)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_143),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_30),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_83),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_118),
.C(n_108),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_165),
.C(n_4),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_141),
.A2(n_104),
.B1(n_112),
.B2(n_101),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_157),
.A2(n_167),
.B1(n_132),
.B2(n_142),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_121),
.A2(n_99),
.B(n_112),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_166),
.B(n_27),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_97),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_170),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_113),
.B1(n_99),
.B2(n_71),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_168),
.B1(n_132),
.B2(n_122),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_125),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_163),
.B(n_164),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_127),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_99),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_115),
.B1(n_88),
.B2(n_80),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_116),
.B1(n_88),
.B2(n_80),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_66),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_143),
.B1(n_144),
.B2(n_121),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_171),
.A2(n_174),
.B1(n_177),
.B2(n_180),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_130),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_173),
.A2(n_181),
.B(n_182),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_122),
.B(n_124),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_179),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_136),
.Y(n_176)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_149),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_1),
.B(n_3),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_27),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_184),
.Y(n_196)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_27),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_186),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_1),
.B(n_3),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_4),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_190),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_189),
.C(n_169),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_16),
.C(n_15),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_161),
.B1(n_162),
.B2(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_157),
.B1(n_166),
.B2(n_164),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_203),
.Y(n_208)
);

AOI321xp33_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_153),
.A3(n_169),
.B1(n_167),
.B2(n_152),
.C(n_163),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_198),
.B(n_195),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_188),
.C(n_177),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_194),
.B(n_181),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_156),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_200),
.C(n_205),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_156),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_178),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_179),
.A2(n_148),
.B1(n_5),
.B2(n_6),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_16),
.C(n_14),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_212),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_211),
.B(n_218),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_185),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_213),
.A2(n_14),
.B1(n_13),
.B2(n_6),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_189),
.C(n_178),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_217),
.C(n_205),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_175),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_197),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_201),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_187),
.C(n_190),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_184),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_13),
.C(n_5),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_199),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_223),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_222),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_191),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_208),
.Y(n_229)
);

AO22x1_ASAP7_75t_L g226 ( 
.A1(n_218),
.A2(n_194),
.B1(n_193),
.B2(n_186),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_228),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_216),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_232),
.Y(n_237)
);

NOR2xp67_ASAP7_75t_R g232 ( 
.A(n_226),
.B(n_210),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_235),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_234),
.A2(n_220),
.B1(n_219),
.B2(n_224),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_240),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_234),
.A2(n_224),
.B1(n_7),
.B2(n_9),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_238),
.A2(n_4),
.B1(n_7),
.B2(n_9),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_11),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_230),
.B(n_7),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_243),
.B(n_238),
.Y(n_244)
);

FAx1_ASAP7_75t_SL g246 ( 
.A(n_244),
.B(n_245),
.CI(n_10),
.CON(n_246),
.SN(n_246)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_239),
.C(n_10),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_246),
.A2(n_10),
.B(n_244),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_246),
.Y(n_248)
);


endmodule