module fake_netlist_1_11340_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVxp67_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
BUFx2_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
CKINVDCx16_ASAP7_75t_R g5 ( .A(n_4), .Y(n_5) );
OAI21x1_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_6) );
NAND2xp5_ASAP7_75t_L g7 ( .A(n_5), .B(n_3), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_5), .B(n_2), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
AOI221xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_8), .B1(n_6), .B2(n_2), .C(n_1), .Y(n_10) );
INVx1_ASAP7_75t_SL g11 ( .A(n_9), .Y(n_11) );
OR2x6_ASAP7_75t_L g12 ( .A(n_11), .B(n_6), .Y(n_12) );
AOI22xp33_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_0), .B1(n_10), .B2(n_9), .Y(n_13) );
endmodule