module real_aes_8229_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g554 ( .A1(n_0), .A2(n_172), .B(n_555), .C(n_558), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_1), .B(n_543), .Y(n_559) );
INVx1_ASAP7_75t_L g421 ( .A(n_2), .Y(n_421) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_3), .A2(n_107), .B1(n_414), .B2(n_415), .Y(n_106) );
INVx1_ASAP7_75t_L g415 ( .A(n_3), .Y(n_415) );
INVx1_ASAP7_75t_L g190 ( .A(n_4), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_5), .B(n_161), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_6), .A2(n_458), .B(n_537), .Y(n_536) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_7), .A2(n_137), .B(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_8), .A2(n_38), .B1(n_117), .B2(n_126), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_9), .B(n_137), .Y(n_201) );
AND2x6_ASAP7_75t_L g135 ( .A(n_10), .B(n_136), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_11), .A2(n_135), .B(n_461), .C(n_518), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_12), .B(n_39), .Y(n_422) );
INVx1_ASAP7_75t_L g133 ( .A(n_13), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_14), .B(n_124), .Y(n_144) );
INVx1_ASAP7_75t_L g182 ( .A(n_15), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_16), .B(n_161), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_17), .B(n_138), .Y(n_206) );
AO32x2_ASAP7_75t_L g169 ( .A1(n_18), .A2(n_134), .A3(n_137), .B1(n_170), .B2(n_174), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_19), .B(n_126), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_20), .B(n_138), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_21), .A2(n_54), .B1(n_117), .B2(n_126), .Y(n_173) );
AOI22xp33_ASAP7_75t_SL g123 ( .A1(n_22), .A2(n_81), .B1(n_124), .B2(n_126), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_23), .B(n_126), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_24), .A2(n_134), .B(n_461), .C(n_463), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_25), .A2(n_134), .B(n_461), .C(n_508), .Y(n_507) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_26), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_27), .B(n_129), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_28), .Y(n_427) );
OAI22xp5_ASAP7_75t_SL g745 ( .A1(n_29), .A2(n_746), .B1(n_749), .B2(n_750), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_29), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_30), .A2(n_458), .B(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_31), .B(n_129), .Y(n_167) );
INVx2_ASAP7_75t_L g119 ( .A(n_32), .Y(n_119) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_33), .A2(n_482), .B(n_491), .C(n_493), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_34), .B(n_126), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_35), .B(n_129), .Y(n_151) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_36), .A2(n_75), .B1(n_747), .B2(n_748), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_36), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_37), .B(n_146), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_40), .B(n_457), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_41), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_42), .B(n_161), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_43), .B(n_458), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_44), .A2(n_482), .B(n_491), .C(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_45), .A2(n_79), .B1(n_412), .B2(n_413), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_45), .Y(n_412) );
OAI22xp5_ASAP7_75t_SL g442 ( .A1(n_45), .A2(n_412), .B1(n_443), .B2(n_444), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_46), .B(n_126), .Y(n_196) );
INVx1_ASAP7_75t_L g556 ( .A(n_47), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g116 ( .A1(n_48), .A2(n_89), .B1(n_117), .B2(n_120), .Y(n_116) );
INVx1_ASAP7_75t_L g529 ( .A(n_49), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_50), .B(n_126), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_51), .B(n_126), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_52), .B(n_458), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_53), .B(n_188), .Y(n_200) );
AOI22xp33_ASAP7_75t_SL g210 ( .A1(n_55), .A2(n_59), .B1(n_124), .B2(n_126), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_56), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_57), .B(n_126), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_58), .B(n_126), .Y(n_225) );
INVx1_ASAP7_75t_L g136 ( .A(n_60), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_61), .B(n_458), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_62), .B(n_543), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_63), .A2(n_185), .B(n_188), .C(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_64), .B(n_126), .Y(n_191) );
INVx1_ASAP7_75t_L g132 ( .A(n_65), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_66), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_67), .B(n_161), .Y(n_495) );
AO32x2_ASAP7_75t_L g114 ( .A1(n_68), .A2(n_115), .A3(n_128), .B1(n_134), .B2(n_137), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_69), .B(n_127), .Y(n_519) );
INVx1_ASAP7_75t_L g224 ( .A(n_70), .Y(n_224) );
INVx1_ASAP7_75t_L g159 ( .A(n_71), .Y(n_159) );
CKINVDCx16_ASAP7_75t_R g553 ( .A(n_72), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_73), .B(n_465), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_74), .A2(n_461), .B(n_478), .C(n_482), .Y(n_477) );
INVx1_ASAP7_75t_L g748 ( .A(n_75), .Y(n_748) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_76), .B(n_124), .Y(n_160) );
CKINVDCx16_ASAP7_75t_R g538 ( .A(n_77), .Y(n_538) );
INVx1_ASAP7_75t_L g435 ( .A(n_78), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_79), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_80), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_82), .B(n_117), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_83), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_84), .B(n_124), .Y(n_164) );
INVx2_ASAP7_75t_L g130 ( .A(n_85), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_86), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_87), .B(n_121), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_88), .B(n_124), .Y(n_197) );
OR2x2_ASAP7_75t_L g418 ( .A(n_90), .B(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g447 ( .A(n_90), .B(n_420), .Y(n_447) );
INVx2_ASAP7_75t_L g744 ( .A(n_90), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_91), .A2(n_102), .B1(n_124), .B2(n_125), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_92), .B(n_458), .Y(n_489) );
INVx1_ASAP7_75t_L g494 ( .A(n_93), .Y(n_494) );
AOI222xp33_ASAP7_75t_L g440 ( .A1(n_94), .A2(n_441), .B1(n_745), .B2(n_751), .C1(n_756), .C2(n_757), .Y(n_440) );
INVxp67_ASAP7_75t_L g541 ( .A(n_95), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_96), .B(n_124), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_97), .B(n_435), .Y(n_434) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_98), .A2(n_104), .B1(n_428), .B2(n_436), .C1(n_439), .C2(n_760), .Y(n_103) );
AOI321xp33_ASAP7_75t_L g105 ( .A1(n_98), .A2(n_106), .A3(n_416), .B1(n_423), .B2(n_424), .C(n_426), .Y(n_105) );
INVx1_ASAP7_75t_L g423 ( .A(n_98), .Y(n_423) );
INVx1_ASAP7_75t_L g479 ( .A(n_99), .Y(n_479) );
INVx1_ASAP7_75t_L g515 ( .A(n_100), .Y(n_515) );
AND2x2_ASAP7_75t_L g531 ( .A(n_101), .B(n_129), .Y(n_531) );
INVxp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_106), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g414 ( .A(n_107), .Y(n_414) );
XOR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_411), .Y(n_107) );
INVx2_ASAP7_75t_L g443 ( .A(n_108), .Y(n_443) );
AND3x1_ASAP7_75t_L g108 ( .A(n_109), .B(n_331), .C(n_379), .Y(n_108) );
NOR4xp25_ASAP7_75t_L g109 ( .A(n_110), .B(n_259), .C(n_304), .D(n_318), .Y(n_109) );
OAI311xp33_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_175), .A3(n_202), .B1(n_212), .C1(n_227), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_139), .Y(n_111) );
OAI21xp33_ASAP7_75t_L g212 ( .A1(n_112), .A2(n_213), .B(n_215), .Y(n_212) );
AND2x2_ASAP7_75t_L g320 ( .A(n_112), .B(n_247), .Y(n_320) );
AND2x2_ASAP7_75t_L g377 ( .A(n_112), .B(n_263), .Y(n_377) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g270 ( .A(n_113), .B(n_168), .Y(n_270) );
AND2x2_ASAP7_75t_L g327 ( .A(n_113), .B(n_275), .Y(n_327) );
INVx1_ASAP7_75t_L g368 ( .A(n_113), .Y(n_368) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_114), .Y(n_236) );
AND2x2_ASAP7_75t_L g277 ( .A(n_114), .B(n_168), .Y(n_277) );
AND2x2_ASAP7_75t_L g281 ( .A(n_114), .B(n_169), .Y(n_281) );
INVx1_ASAP7_75t_L g293 ( .A(n_114), .Y(n_293) );
OAI22xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_121), .B1(n_123), .B2(n_127), .Y(n_115) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx3_ASAP7_75t_L g120 ( .A(n_118), .Y(n_120) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_118), .Y(n_126) );
AND2x6_ASAP7_75t_L g461 ( .A(n_118), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g125 ( .A(n_119), .Y(n_125) );
INVx1_ASAP7_75t_L g189 ( .A(n_119), .Y(n_189) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_120), .Y(n_496) );
INVx2_ASAP7_75t_L g558 ( .A(n_120), .Y(n_558) );
INVx2_ASAP7_75t_L g150 ( .A(n_121), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_121), .A2(n_171), .B1(n_172), .B2(n_173), .Y(n_170) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_121), .A2(n_172), .B1(n_209), .B2(n_210), .Y(n_208) );
INVx4_ASAP7_75t_L g557 ( .A(n_121), .Y(n_557) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx3_ASAP7_75t_L g127 ( .A(n_122), .Y(n_127) );
INVx1_ASAP7_75t_L g146 ( .A(n_122), .Y(n_146) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_122), .Y(n_166) );
AND2x2_ASAP7_75t_L g459 ( .A(n_122), .B(n_189), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_122), .Y(n_462) );
INVx2_ASAP7_75t_L g183 ( .A(n_124), .Y(n_183) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx3_ASAP7_75t_L g158 ( .A(n_126), .Y(n_158) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_126), .Y(n_481) );
INVx5_ASAP7_75t_L g161 ( .A(n_127), .Y(n_161) );
INVx1_ASAP7_75t_L g468 ( .A(n_128), .Y(n_468) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_129), .A2(n_141), .B(n_151), .Y(n_140) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_129), .A2(n_156), .B(n_167), .Y(n_155) );
INVx1_ASAP7_75t_L g471 ( .A(n_129), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_129), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_129), .A2(n_526), .B(n_527), .Y(n_525) );
AND2x2_ASAP7_75t_SL g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_L g138 ( .A(n_130), .B(n_131), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
NAND3xp33_ASAP7_75t_L g207 ( .A(n_134), .B(n_208), .C(n_211), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_134), .A2(n_220), .B(n_223), .Y(n_219) );
BUFx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI21xp5_ASAP7_75t_L g141 ( .A1(n_135), .A2(n_142), .B(n_147), .Y(n_141) );
OAI21xp5_ASAP7_75t_L g156 ( .A1(n_135), .A2(n_157), .B(n_162), .Y(n_156) );
OAI21xp5_ASAP7_75t_L g180 ( .A1(n_135), .A2(n_181), .B(n_186), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_135), .A2(n_195), .B(n_198), .Y(n_194) );
AND2x4_ASAP7_75t_L g458 ( .A(n_135), .B(n_459), .Y(n_458) );
INVx4_ASAP7_75t_SL g483 ( .A(n_135), .Y(n_483) );
NAND2x1p5_ASAP7_75t_L g516 ( .A(n_135), .B(n_459), .Y(n_516) );
OA21x2_ASAP7_75t_L g193 ( .A1(n_137), .A2(n_194), .B(n_201), .Y(n_193) );
INVx4_ASAP7_75t_L g211 ( .A(n_137), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_137), .A2(n_506), .B(n_507), .Y(n_505) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_137), .Y(n_535) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g174 ( .A(n_138), .Y(n_174) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_152), .Y(n_139) );
AND2x2_ASAP7_75t_L g214 ( .A(n_140), .B(n_168), .Y(n_214) );
INVx2_ASAP7_75t_L g248 ( .A(n_140), .Y(n_248) );
AND2x2_ASAP7_75t_L g263 ( .A(n_140), .B(n_169), .Y(n_263) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_140), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_140), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g283 ( .A(n_140), .B(n_246), .Y(n_283) );
INVx1_ASAP7_75t_L g295 ( .A(n_140), .Y(n_295) );
INVx1_ASAP7_75t_L g336 ( .A(n_140), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_140), .B(n_236), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_145), .Y(n_142) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_150), .Y(n_147) );
O2A1O1Ixp5_ASAP7_75t_L g223 ( .A1(n_150), .A2(n_187), .B(n_224), .C(n_225), .Y(n_223) );
NOR2xp67_ASAP7_75t_L g152 ( .A(n_153), .B(n_168), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g213 ( .A(n_154), .B(n_214), .Y(n_213) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_154), .Y(n_241) );
AND2x2_ASAP7_75t_SL g294 ( .A(n_154), .B(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g298 ( .A(n_154), .B(n_168), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_154), .B(n_293), .Y(n_356) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g246 ( .A(n_155), .Y(n_246) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_155), .Y(n_262) );
OR2x2_ASAP7_75t_L g335 ( .A(n_155), .B(n_336), .Y(n_335) );
O2A1O1Ixp5_ASAP7_75t_SL g157 ( .A1(n_158), .A2(n_159), .B(n_160), .C(n_161), .Y(n_157) );
INVx2_ASAP7_75t_L g172 ( .A(n_161), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_161), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_161), .A2(n_221), .B(n_222), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_161), .B(n_541), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_165), .Y(n_162) );
INVx1_ASAP7_75t_L g185 ( .A(n_165), .Y(n_185) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g465 ( .A(n_166), .Y(n_465) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx2_ASAP7_75t_L g242 ( .A(n_169), .Y(n_242) );
AND2x2_ASAP7_75t_L g247 ( .A(n_169), .B(n_248), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g186 ( .A1(n_172), .A2(n_187), .B(n_190), .C(n_191), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_172), .A2(n_199), .B(n_200), .Y(n_198) );
INVx2_ASAP7_75t_L g179 ( .A(n_174), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_174), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_175), .B(n_230), .Y(n_393) );
INVx1_ASAP7_75t_SL g175 ( .A(n_176), .Y(n_175) );
OR2x2_ASAP7_75t_L g363 ( .A(n_176), .B(n_204), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_193), .Y(n_176) );
AND2x2_ASAP7_75t_L g239 ( .A(n_177), .B(n_230), .Y(n_239) );
INVx2_ASAP7_75t_L g251 ( .A(n_177), .Y(n_251) );
AND2x2_ASAP7_75t_L g285 ( .A(n_177), .B(n_233), .Y(n_285) );
AND2x2_ASAP7_75t_L g352 ( .A(n_177), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_178), .B(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g232 ( .A(n_178), .B(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g272 ( .A(n_178), .B(n_193), .Y(n_272) );
AND2x2_ASAP7_75t_L g289 ( .A(n_178), .B(n_290), .Y(n_289) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_192), .Y(n_178) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_179), .A2(n_219), .B(n_226), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_184), .C(n_185), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_183), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_183), .A2(n_519), .B(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_185), .A2(n_479), .B(n_480), .C(n_481), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_187), .A2(n_464), .B(n_466), .Y(n_463) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g215 ( .A(n_193), .B(n_216), .Y(n_215) );
INVx3_ASAP7_75t_L g233 ( .A(n_193), .Y(n_233) );
AND2x2_ASAP7_75t_L g238 ( .A(n_193), .B(n_218), .Y(n_238) );
AND2x2_ASAP7_75t_L g311 ( .A(n_193), .B(n_290), .Y(n_311) );
AND2x2_ASAP7_75t_L g376 ( .A(n_193), .B(n_366), .Y(n_376) );
OAI311xp33_ASAP7_75t_L g259 ( .A1(n_202), .A2(n_260), .A3(n_264), .B1(n_266), .C1(n_286), .Y(n_259) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g271 ( .A(n_203), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g330 ( .A(n_203), .B(n_238), .Y(n_330) );
AND2x2_ASAP7_75t_L g404 ( .A(n_203), .B(n_285), .Y(n_404) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_204), .B(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g339 ( .A(n_204), .Y(n_339) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx3_ASAP7_75t_L g230 ( .A(n_205), .Y(n_230) );
NOR2x1_ASAP7_75t_L g302 ( .A(n_205), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g359 ( .A(n_205), .B(n_233), .Y(n_359) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
INVx1_ASAP7_75t_L g256 ( .A(n_206), .Y(n_256) );
AO21x1_ASAP7_75t_L g255 ( .A1(n_208), .A2(n_211), .B(n_256), .Y(n_255) );
AO21x2_ASAP7_75t_L g475 ( .A1(n_211), .A2(n_476), .B(n_485), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_211), .B(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_211), .B(n_498), .Y(n_497) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_211), .A2(n_514), .B(n_521), .Y(n_513) );
INVx3_ASAP7_75t_L g543 ( .A(n_211), .Y(n_543) );
AND2x2_ASAP7_75t_L g234 ( .A(n_214), .B(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g287 ( .A(n_214), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g367 ( .A(n_214), .B(n_368), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g266 ( .A1(n_215), .A2(n_247), .B1(n_267), .B2(n_271), .C(n_273), .Y(n_266) );
INVx1_ASAP7_75t_L g391 ( .A(n_216), .Y(n_391) );
OR2x2_ASAP7_75t_L g357 ( .A(n_217), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g252 ( .A(n_218), .B(n_233), .Y(n_252) );
OR2x2_ASAP7_75t_L g254 ( .A(n_218), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g279 ( .A(n_218), .Y(n_279) );
INVx2_ASAP7_75t_L g290 ( .A(n_218), .Y(n_290) );
AND2x2_ASAP7_75t_L g317 ( .A(n_218), .B(n_255), .Y(n_317) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_218), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_234), .B1(n_237), .B2(n_240), .C(n_243), .Y(n_227) );
INVx1_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
AND2x2_ASAP7_75t_L g328 ( .A(n_230), .B(n_238), .Y(n_328) );
AND2x2_ASAP7_75t_L g378 ( .A(n_230), .B(n_232), .Y(n_378) );
INVx2_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g265 ( .A(n_232), .B(n_236), .Y(n_265) );
AND2x2_ASAP7_75t_L g344 ( .A(n_232), .B(n_317), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_233), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g303 ( .A(n_233), .Y(n_303) );
OAI21xp33_ASAP7_75t_L g313 ( .A1(n_234), .A2(n_314), .B(n_316), .Y(n_313) );
OR2x2_ASAP7_75t_L g257 ( .A(n_235), .B(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g323 ( .A(n_235), .B(n_283), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_235), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g300 ( .A(n_236), .B(n_269), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_236), .B(n_383), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_237), .B(n_263), .Y(n_373) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AND2x2_ASAP7_75t_L g296 ( .A(n_238), .B(n_251), .Y(n_296) );
INVx1_ASAP7_75t_L g312 ( .A(n_239), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_249), .B1(n_253), .B2(n_257), .Y(n_243) );
INVx2_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g275 ( .A(n_246), .Y(n_275) );
INVx1_ASAP7_75t_L g288 ( .A(n_246), .Y(n_288) );
INVx1_ASAP7_75t_L g258 ( .A(n_247), .Y(n_258) );
AND2x2_ASAP7_75t_L g329 ( .A(n_247), .B(n_275), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_247), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_252), .Y(n_249) );
OR2x2_ASAP7_75t_L g253 ( .A(n_250), .B(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_250), .B(n_366), .Y(n_365) );
NOR2xp67_ASAP7_75t_L g397 ( .A(n_250), .B(n_398), .Y(n_397) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g400 ( .A(n_252), .B(n_352), .Y(n_400) );
INVx1_ASAP7_75t_SL g366 ( .A(n_254), .Y(n_366) );
AND2x2_ASAP7_75t_L g306 ( .A(n_255), .B(n_290), .Y(n_306) );
INVx1_ASAP7_75t_L g353 ( .A(n_255), .Y(n_353) );
OAI222xp33_ASAP7_75t_L g394 ( .A1(n_260), .A2(n_350), .B1(n_395), .B2(n_396), .C1(n_399), .C2(n_401), .Y(n_394) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx1_ASAP7_75t_L g315 ( .A(n_262), .Y(n_315) );
AND2x2_ASAP7_75t_L g326 ( .A(n_263), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_263), .B(n_368), .Y(n_395) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_265), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g370 ( .A(n_267), .Y(n_370) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_SL g308 ( .A(n_270), .Y(n_308) );
AND2x2_ASAP7_75t_L g387 ( .A(n_270), .B(n_348), .Y(n_387) );
AND2x2_ASAP7_75t_L g410 ( .A(n_270), .B(n_294), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_272), .B(n_306), .Y(n_305) );
OAI32xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_276), .A3(n_278), .B1(n_280), .B2(n_284), .Y(n_273) );
BUFx2_ASAP7_75t_L g348 ( .A(n_275), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_276), .B(n_294), .Y(n_375) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g314 ( .A(n_277), .B(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g382 ( .A(n_277), .B(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g371 ( .A(n_278), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x2_ASAP7_75t_L g342 ( .A(n_281), .B(n_315), .Y(n_342) );
INVx2_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
OAI221xp5_ASAP7_75t_SL g304 ( .A1(n_283), .A2(n_305), .B1(n_307), .B2(n_309), .C(n_313), .Y(n_304) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g316 ( .A(n_285), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g322 ( .A(n_285), .B(n_306), .Y(n_322) );
AOI221xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_289), .B1(n_291), .B2(n_296), .C(n_297), .Y(n_286) );
INVx1_ASAP7_75t_L g405 ( .A(n_287), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_288), .B(n_382), .Y(n_381) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_289), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_294), .B(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g360 ( .A(n_294), .Y(n_360) );
BUFx3_ASAP7_75t_L g383 ( .A(n_295), .Y(n_383) );
INVx1_ASAP7_75t_SL g324 ( .A(n_296), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_296), .B(n_338), .Y(n_337) );
AOI21xp33_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_299), .B(n_301), .Y(n_297) );
OAI221xp5_ASAP7_75t_L g402 ( .A1(n_298), .A2(n_399), .B1(n_403), .B2(n_405), .C(n_406), .Y(n_402) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g345 ( .A(n_303), .B(n_306), .Y(n_345) );
INVx1_ASAP7_75t_L g409 ( .A(n_303), .Y(n_409) );
INVx2_ASAP7_75t_L g398 ( .A(n_306), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_306), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g351 ( .A(n_311), .B(n_352), .Y(n_351) );
OAI221xp5_ASAP7_75t_SL g318 ( .A1(n_319), .A2(n_321), .B1(n_323), .B2(n_324), .C(n_325), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_328), .B1(n_329), .B2(n_330), .Y(n_325) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_327), .A2(n_389), .B1(n_390), .B2(n_392), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g406 ( .A1(n_330), .A2(n_407), .B(n_410), .Y(n_406) );
NOR4xp25_ASAP7_75t_SL g331 ( .A(n_332), .B(n_340), .C(n_349), .D(n_369), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_337), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .B1(n_346), .B2(n_347), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g385 ( .A(n_345), .Y(n_385) );
OAI221xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_354), .B1(n_357), .B2(n_360), .C(n_361), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g372 ( .A(n_352), .Y(n_372) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI21xp5_ASAP7_75t_SL g361 ( .A1(n_362), .A2(n_364), .B(n_367), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI211xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B(n_373), .C(n_374), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B1(n_377), .B2(n_378), .Y(n_374) );
CKINVDCx14_ASAP7_75t_R g384 ( .A(n_378), .Y(n_384) );
NOR3xp33_ASAP7_75t_L g379 ( .A(n_380), .B(n_394), .C(n_402), .Y(n_379) );
OAI221xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_384), .B1(n_385), .B2(n_386), .C(n_388), .Y(n_380) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
CKINVDCx16_ASAP7_75t_R g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2xp33_ASAP7_75t_L g761 ( .A(n_416), .B(n_762), .Y(n_761) );
INVx1_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g425 ( .A(n_418), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_418), .B(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g438 ( .A(n_418), .Y(n_438) );
NOR2x2_ASAP7_75t_L g759 ( .A(n_419), .B(n_744), .Y(n_759) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OR2x2_ASAP7_75t_L g743 ( .A(n_420), .B(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_433), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OA21x2_ASAP7_75t_L g437 ( .A1(n_432), .A2(n_433), .B(n_438), .Y(n_437) );
NOR2xp33_ASAP7_75t_SL g762 ( .A(n_432), .B(n_434), .Y(n_762) );
INVx1_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx3_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI22xp5_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_445), .B1(n_448), .B2(n_741), .Y(n_441) );
INVx1_ASAP7_75t_L g752 ( .A(n_442), .Y(n_752) );
INVx2_ASAP7_75t_L g444 ( .A(n_443), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g753 ( .A(n_446), .Y(n_753) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx2_ASAP7_75t_L g754 ( .A(n_449), .Y(n_754) );
AND3x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_645), .C(n_702), .Y(n_449) );
NOR3xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_590), .C(n_626), .Y(n_450) );
OAI211xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_499), .B(n_545), .C(n_577), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_472), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x4_ASAP7_75t_L g548 ( .A(n_454), .B(n_549), .Y(n_548) );
INVx5_ASAP7_75t_L g576 ( .A(n_454), .Y(n_576) );
AND2x2_ASAP7_75t_L g649 ( .A(n_454), .B(n_565), .Y(n_649) );
AND2x2_ASAP7_75t_L g687 ( .A(n_454), .B(n_593), .Y(n_687) );
AND2x2_ASAP7_75t_L g707 ( .A(n_454), .B(n_550), .Y(n_707) );
OR2x6_ASAP7_75t_L g454 ( .A(n_455), .B(n_469), .Y(n_454) );
AOI21xp5_ASAP7_75t_SL g455 ( .A1(n_456), .A2(n_460), .B(n_468), .Y(n_455) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx5_ASAP7_75t_L g492 ( .A(n_461), .Y(n_492) );
INVx2_ASAP7_75t_L g467 ( .A(n_465), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_467), .A2(n_494), .B(n_495), .C(n_496), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_467), .A2(n_496), .B(n_529), .C(n_530), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_472), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_487), .Y(n_472) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_473), .Y(n_588) );
AND2x2_ASAP7_75t_L g602 ( .A(n_473), .B(n_549), .Y(n_602) );
INVx1_ASAP7_75t_L g625 ( .A(n_473), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_473), .B(n_576), .Y(n_664) );
OR2x2_ASAP7_75t_L g701 ( .A(n_473), .B(n_547), .Y(n_701) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_474), .Y(n_637) );
AND2x2_ASAP7_75t_L g644 ( .A(n_474), .B(n_550), .Y(n_644) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g565 ( .A(n_475), .B(n_550), .Y(n_565) );
BUFx2_ASAP7_75t_L g593 ( .A(n_475), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_484), .Y(n_476) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g537 ( .A1(n_483), .A2(n_492), .B(n_538), .C(n_539), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_SL g552 ( .A1(n_483), .A2(n_492), .B(n_553), .C(n_554), .Y(n_552) );
INVx5_ASAP7_75t_L g547 ( .A(n_487), .Y(n_547) );
BUFx2_ASAP7_75t_L g569 ( .A(n_487), .Y(n_569) );
AND2x2_ASAP7_75t_L g726 ( .A(n_487), .B(n_580), .Y(n_726) );
OR2x6_ASAP7_75t_L g487 ( .A(n_488), .B(n_497), .Y(n_487) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_532), .Y(n_500) );
OAI221xp5_ASAP7_75t_L g626 ( .A1(n_501), .A2(n_627), .B1(n_634), .B2(n_635), .C(n_638), .Y(n_626) );
OR2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_511), .Y(n_501) );
AND2x2_ASAP7_75t_L g533 ( .A(n_502), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_502), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g561 ( .A(n_503), .B(n_512), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_503), .B(n_513), .Y(n_571) );
OR2x2_ASAP7_75t_L g582 ( .A(n_503), .B(n_534), .Y(n_582) );
AND2x2_ASAP7_75t_L g585 ( .A(n_503), .B(n_573), .Y(n_585) );
AND2x2_ASAP7_75t_L g601 ( .A(n_503), .B(n_523), .Y(n_601) );
OR2x2_ASAP7_75t_L g617 ( .A(n_503), .B(n_513), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_503), .B(n_534), .Y(n_679) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_504), .B(n_523), .Y(n_671) );
AND2x2_ASAP7_75t_L g674 ( .A(n_504), .B(n_513), .Y(n_674) );
OR2x2_ASAP7_75t_L g595 ( .A(n_511), .B(n_582), .Y(n_595) );
INVx2_ASAP7_75t_L g621 ( .A(n_511), .Y(n_621) );
OR2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_523), .Y(n_511) );
AND2x2_ASAP7_75t_L g544 ( .A(n_512), .B(n_524), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_512), .B(n_534), .Y(n_600) );
OR2x2_ASAP7_75t_L g611 ( .A(n_512), .B(n_524), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_512), .B(n_573), .Y(n_670) );
OAI221xp5_ASAP7_75t_L g703 ( .A1(n_512), .A2(n_704), .B1(n_706), .B2(n_708), .C(n_711), .Y(n_703) );
INVx5_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_513), .B(n_534), .Y(n_642) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_517), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_523), .B(n_573), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_523), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g589 ( .A(n_523), .B(n_561), .Y(n_589) );
OR2x2_ASAP7_75t_L g633 ( .A(n_523), .B(n_534), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_523), .B(n_585), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_523), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g698 ( .A(n_523), .B(n_699), .Y(n_698) );
INVx5_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_SL g562 ( .A(n_524), .B(n_533), .Y(n_562) );
O2A1O1Ixp33_ASAP7_75t_SL g566 ( .A1(n_524), .A2(n_567), .B(n_570), .C(n_574), .Y(n_566) );
OR2x2_ASAP7_75t_L g604 ( .A(n_524), .B(n_600), .Y(n_604) );
OR2x2_ASAP7_75t_L g640 ( .A(n_524), .B(n_582), .Y(n_640) );
OAI311xp33_ASAP7_75t_L g646 ( .A1(n_524), .A2(n_585), .A3(n_647), .B1(n_650), .C1(n_657), .Y(n_646) );
AND2x2_ASAP7_75t_L g697 ( .A(n_524), .B(n_534), .Y(n_697) );
AND2x2_ASAP7_75t_L g705 ( .A(n_524), .B(n_560), .Y(n_705) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_524), .Y(n_723) );
AND2x2_ASAP7_75t_L g740 ( .A(n_524), .B(n_561), .Y(n_740) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_531), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_544), .Y(n_532) );
AND2x2_ASAP7_75t_L g568 ( .A(n_533), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g724 ( .A(n_533), .Y(n_724) );
AND2x2_ASAP7_75t_L g560 ( .A(n_534), .B(n_561), .Y(n_560) );
INVx3_ASAP7_75t_L g573 ( .A(n_534), .Y(n_573) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_534), .Y(n_616) );
INVxp67_ASAP7_75t_L g655 ( .A(n_534), .Y(n_655) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B(n_542), .Y(n_534) );
OA21x2_ASAP7_75t_L g550 ( .A1(n_543), .A2(n_551), .B(n_559), .Y(n_550) );
AND2x2_ASAP7_75t_L g733 ( .A(n_544), .B(n_581), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_560), .B1(n_562), .B2(n_563), .C(n_566), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_547), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g586 ( .A(n_547), .B(n_576), .Y(n_586) );
AND2x2_ASAP7_75t_L g594 ( .A(n_547), .B(n_549), .Y(n_594) );
OR2x2_ASAP7_75t_L g606 ( .A(n_547), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g624 ( .A(n_547), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g648 ( .A(n_547), .B(n_649), .Y(n_648) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_547), .Y(n_668) );
AND2x2_ASAP7_75t_L g720 ( .A(n_547), .B(n_644), .Y(n_720) );
OAI31xp33_ASAP7_75t_L g728 ( .A1(n_547), .A2(n_597), .A3(n_696), .B(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_548), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g692 ( .A(n_548), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_548), .B(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g580 ( .A(n_549), .B(n_576), .Y(n_580) );
INVx1_ASAP7_75t_L g667 ( .A(n_549), .Y(n_667) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g717 ( .A(n_550), .B(n_576), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
INVx1_ASAP7_75t_SL g727 ( .A(n_560), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_561), .B(n_632), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_562), .A2(n_674), .B1(n_712), .B2(n_715), .Y(n_711) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g575 ( .A(n_565), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g634 ( .A(n_565), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_565), .B(n_586), .Y(n_739) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g709 ( .A(n_568), .B(n_710), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_569), .A2(n_628), .B(n_630), .Y(n_627) );
OR2x2_ASAP7_75t_L g635 ( .A(n_569), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g656 ( .A(n_569), .B(n_644), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_569), .B(n_667), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_569), .B(n_707), .Y(n_706) );
OAI221xp5_ASAP7_75t_SL g683 ( .A1(n_570), .A2(n_684), .B1(n_689), .B2(n_692), .C(n_693), .Y(n_683) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
OR2x2_ASAP7_75t_L g660 ( .A(n_571), .B(n_633), .Y(n_660) );
INVx1_ASAP7_75t_L g699 ( .A(n_571), .Y(n_699) );
INVx2_ASAP7_75t_L g675 ( .A(n_572), .Y(n_675) );
INVx1_ASAP7_75t_L g609 ( .A(n_573), .Y(n_609) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g614 ( .A(n_576), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_576), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g643 ( .A(n_576), .B(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g731 ( .A(n_576), .B(n_701), .Y(n_731) );
AOI222xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .B1(n_583), .B2(n_586), .C1(n_587), .C2(n_589), .Y(n_577) );
INVxp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g587 ( .A(n_580), .B(n_588), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_580), .A2(n_630), .B1(n_658), .B2(n_659), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_580), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
OAI21xp33_ASAP7_75t_SL g618 ( .A1(n_589), .A2(n_619), .B(n_622), .Y(n_618) );
OAI211xp5_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_595), .B(n_596), .C(n_618), .Y(n_590) );
INVxp67_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AOI221xp5_ASAP7_75t_L g596 ( .A1(n_594), .A2(n_597), .B1(n_602), .B2(n_603), .C(n_605), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_594), .B(n_682), .Y(n_681) );
INVxp67_ASAP7_75t_L g688 ( .A(n_594), .Y(n_688) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
AND2x2_ASAP7_75t_L g690 ( .A(n_599), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g607 ( .A(n_602), .Y(n_607) );
AND2x2_ASAP7_75t_L g613 ( .A(n_602), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_608), .B1(n_612), .B2(n_615), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_609), .B(n_621), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_610), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g710 ( .A(n_614), .Y(n_710) );
AND2x2_ASAP7_75t_L g729 ( .A(n_614), .B(n_644), .Y(n_729) );
OR2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_621), .B(n_678), .Y(n_737) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_624), .B(n_692), .Y(n_735) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g658 ( .A(n_636), .Y(n_658) );
BUFx2_ASAP7_75t_L g682 ( .A(n_637), .Y(n_682) );
OAI21xp5_ASAP7_75t_SL g638 ( .A1(n_639), .A2(n_641), .B(n_643), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NOR3xp33_ASAP7_75t_L g645 ( .A(n_646), .B(n_661), .C(n_683), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI21xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_653), .B(n_656), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
A2O1A1Ixp33_ASAP7_75t_SL g661 ( .A1(n_662), .A2(n_665), .B(n_669), .C(n_672), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_662), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NOR2xp67_ASAP7_75t_SL g666 ( .A(n_667), .B(n_668), .Y(n_666) );
OR2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_SL g691 ( .A(n_671), .Y(n_691) );
OAI21xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_676), .B(n_680), .Y(n_672) );
AND2x4_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
AND2x2_ASAP7_75t_L g696 ( .A(n_674), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B1(n_698), .B2(n_700), .Y(n_693) );
INVx2_ASAP7_75t_SL g714 ( .A(n_701), .Y(n_714) );
NOR3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_718), .C(n_730), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVxp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_714), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OAI221xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_721), .B1(n_725), .B2(n_727), .C(n_728), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_L g730 ( .A1(n_719), .A2(n_731), .B(n_732), .C(n_734), .Y(n_730) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B1(n_738), .B2(n_740), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g755 ( .A(n_742), .Y(n_755) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g756 ( .A(n_745), .Y(n_756) );
INVx1_ASAP7_75t_L g749 ( .A(n_746), .Y(n_749) );
OAI22xp5_ASAP7_75t_SL g751 ( .A1(n_752), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_751) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx3_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
endmodule