module fake_jpeg_21755_n_147 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_147);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_7),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_24),
.B(n_11),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_78),
.Y(n_91)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_78),
.B(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_47),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_56),
.B1(n_57),
.B2(n_50),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_62),
.B1(n_64),
.B2(n_51),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_52),
.B1(n_53),
.B2(n_49),
.Y(n_93)
);

BUFx8_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_71),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_99),
.C(n_54),
.Y(n_110)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_96),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_98),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_103),
.B1(n_72),
.B2(n_2),
.Y(n_116)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

CKINVDCx6p67_ASAP7_75t_R g129 ( 
.A(n_107),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_86),
.B1(n_90),
.B2(n_59),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_112),
.B1(n_113),
.B2(n_119),
.Y(n_127)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_21),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_110),
.B(n_117),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_68),
.A3(n_70),
.B1(n_60),
.B2(n_65),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_45),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_67),
.B1(n_66),
.B2(n_55),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_63),
.B1(n_2),
.B2(n_4),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_23),
.B1(n_39),
.B2(n_8),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_124),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_125),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_0),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_118),
.B(n_114),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_134),
.A2(n_128),
.B(n_116),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_136),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_129),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_133),
.B1(n_130),
.B2(n_129),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_131),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_121),
.B(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_113),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

AOI322xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_28),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_16),
.C2(n_17),
.Y(n_143)
);

AOI322xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_32),
.A3(n_20),
.B1(n_29),
.B2(n_30),
.C1(n_36),
.C2(n_33),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_34),
.C(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_6),
.Y(n_147)
);


endmodule