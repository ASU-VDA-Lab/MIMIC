module real_aes_3959_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_889;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_892;
wire n_528;
wire n_202;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_756;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_914;
wire n_203;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_155;
wire n_653;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_922;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_888;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g233 ( .A(n_0), .B(n_165), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_1), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_2), .A2(n_16), .B1(n_897), .B2(n_898), .Y(n_896) );
INVx1_ASAP7_75t_L g898 ( .A(n_2), .Y(n_898) );
O2A1O1Ixp33_ASAP7_75t_SL g169 ( .A1(n_3), .A2(n_129), .B(n_170), .C(n_172), .Y(n_169) );
OAI22xp33_ASAP7_75t_L g238 ( .A1(n_4), .A2(n_84), .B1(n_128), .B2(n_134), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_5), .A2(n_33), .B1(n_544), .B2(n_545), .Y(n_543) );
INVxp67_ASAP7_75t_L g504 ( .A(n_6), .Y(n_504) );
INVx1_ASAP7_75t_L g889 ( .A(n_6), .Y(n_889) );
INVx1_ASAP7_75t_L g892 ( .A(n_6), .Y(n_892) );
BUFx2_ASAP7_75t_L g920 ( .A(n_6), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_7), .A2(n_104), .B1(n_914), .B2(n_924), .Y(n_103) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_8), .A2(n_91), .B1(n_581), .B2(n_582), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_9), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g131 ( .A1(n_10), .A2(n_71), .B1(n_132), .B2(n_134), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_11), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_12), .A2(n_34), .B1(n_529), .B2(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g605 ( .A(n_13), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_14), .A2(n_63), .B1(n_126), .B2(n_128), .Y(n_125) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_15), .A2(n_70), .B(n_143), .Y(n_142) );
OA21x2_ASAP7_75t_L g145 ( .A1(n_15), .A2(n_70), .B(n_143), .Y(n_145) );
INVx1_ASAP7_75t_L g897 ( .A(n_16), .Y(n_897) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_17), .B(n_614), .Y(n_613) );
XOR2x2_ASAP7_75t_L g497 ( .A(n_18), .B(n_51), .Y(n_497) );
INVx1_ASAP7_75t_SL g603 ( .A(n_19), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_20), .B(n_140), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_21), .Y(n_262) );
BUFx3_ASAP7_75t_L g109 ( .A(n_22), .Y(n_109) );
BUFx8_ASAP7_75t_SL g913 ( .A(n_22), .Y(n_913) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_23), .A2(n_177), .B(n_178), .C(n_180), .Y(n_176) );
OAI22xp33_ASAP7_75t_SL g236 ( .A1(n_24), .A2(n_48), .B1(n_128), .B2(n_155), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_25), .A2(n_31), .B1(n_155), .B2(n_160), .Y(n_225) );
O2A1O1Ixp5_ASAP7_75t_L g620 ( .A1(n_26), .A2(n_533), .B(n_621), .C(n_624), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_27), .B(n_550), .Y(n_611) );
O2A1O1Ixp5_ASAP7_75t_L g192 ( .A1(n_28), .A2(n_129), .B(n_193), .C(n_195), .Y(n_192) );
INVx1_ASAP7_75t_L g509 ( .A(n_29), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_29), .B(n_83), .Y(n_923) );
INVx1_ASAP7_75t_SL g629 ( .A(n_30), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_32), .Y(n_112) );
AND2x2_ASAP7_75t_L g921 ( .A(n_35), .B(n_922), .Y(n_921) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_36), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_37), .B(n_210), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_38), .A2(n_42), .B1(n_549), .B2(n_551), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_39), .A2(n_69), .B1(n_551), .B2(n_569), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_40), .B(n_546), .Y(n_610) );
INVx2_ASAP7_75t_L g562 ( .A(n_41), .Y(n_562) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_43), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_44), .B(n_291), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_45), .Y(n_596) );
O2A1O1Ixp33_ASAP7_75t_L g600 ( .A1(n_46), .A2(n_180), .B(n_601), .C(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g678 ( .A(n_47), .Y(n_678) );
INVx2_ASAP7_75t_L g630 ( .A(n_49), .Y(n_630) );
INVx1_ASAP7_75t_L g143 ( .A(n_50), .Y(n_143) );
AND2x4_ASAP7_75t_L g138 ( .A(n_52), .B(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g183 ( .A(n_52), .B(n_139), .Y(n_183) );
INVx2_ASAP7_75t_L g570 ( .A(n_53), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_54), .B(n_511), .Y(n_510) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_55), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_56), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_57), .Y(n_202) );
INVx2_ASAP7_75t_L g161 ( .A(n_58), .Y(n_161) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_59), .A2(n_129), .B(n_264), .C(n_265), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_60), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g893 ( .A1(n_61), .A2(n_894), .B1(n_895), .B2(n_896), .Y(n_893) );
CKINVDCx5p33_ASAP7_75t_R g894 ( .A(n_61), .Y(n_894) );
INVx1_ASAP7_75t_SL g625 ( .A(n_62), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_64), .A2(n_80), .B1(n_171), .B2(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_65), .B(n_140), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_66), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_67), .Y(n_248) );
NAND2xp33_ASAP7_75t_R g144 ( .A(n_68), .B(n_145), .Y(n_144) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_68), .A2(n_102), .B1(n_210), .B2(n_347), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g905 ( .A(n_72), .Y(n_905) );
O2A1O1Ixp33_ASAP7_75t_L g571 ( .A1(n_73), .A2(n_180), .B(n_544), .C(n_572), .Y(n_571) );
OR2x6_ASAP7_75t_L g506 ( .A(n_74), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g918 ( .A(n_74), .Y(n_918) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_75), .Y(n_159) );
CKINVDCx16_ASAP7_75t_R g664 ( .A(n_76), .Y(n_664) );
INVx1_ASAP7_75t_L g674 ( .A(n_77), .Y(n_674) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_78), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_79), .B(n_529), .Y(n_615) );
NOR2xp67_ASAP7_75t_L g597 ( .A(n_81), .B(n_193), .Y(n_597) );
O2A1O1Ixp33_ASAP7_75t_L g565 ( .A1(n_82), .A2(n_129), .B(n_566), .C(n_568), .Y(n_565) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_82), .A2(n_129), .B(n_566), .C(n_568), .Y(n_654) );
INVx1_ASAP7_75t_L g508 ( .A(n_83), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_85), .A2(n_95), .B1(n_535), .B2(n_537), .Y(n_534) );
INVx1_ASAP7_75t_L g922 ( .A(n_86), .Y(n_922) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_87), .Y(n_127) );
BUFx5_ASAP7_75t_L g128 ( .A(n_87), .Y(n_128) );
INVx1_ASAP7_75t_L g133 ( .A(n_87), .Y(n_133) );
INVx2_ASAP7_75t_L g185 ( .A(n_88), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_89), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g268 ( .A(n_90), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_92), .Y(n_179) );
INVx2_ASAP7_75t_SL g139 ( .A(n_93), .Y(n_139) );
INVx1_ASAP7_75t_L g200 ( .A(n_94), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_96), .B(n_145), .Y(n_675) );
INVx1_ASAP7_75t_SL g557 ( .A(n_97), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_98), .B(n_574), .Y(n_632) );
INVx2_ASAP7_75t_L g205 ( .A(n_99), .Y(n_205) );
AND2x2_ASAP7_75t_L g539 ( .A(n_100), .B(n_152), .Y(n_539) );
OAI21xp33_ASAP7_75t_SL g260 ( .A1(n_101), .A2(n_128), .B(n_261), .Y(n_260) );
INVxp67_ASAP7_75t_SL g163 ( .A(n_102), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_102), .B(n_210), .Y(n_209) );
AO21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_110), .B(n_513), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
BUFx8_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
CKINVDCx6p67_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_113), .B(n_498), .C(n_510), .Y(n_110) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_111), .A2(n_113), .B(n_499), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
XNOR2x1_ASAP7_75t_L g113 ( .A(n_114), .B(n_497), .Y(n_113) );
OAI22x1_ASAP7_75t_L g515 ( .A1(n_114), .A2(n_516), .B1(n_888), .B2(n_890), .Y(n_515) );
AO22x2_ASAP7_75t_L g899 ( .A1(n_114), .A2(n_516), .B1(n_900), .B2(n_901), .Y(n_899) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_394), .Y(n_114) );
NOR3xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_305), .C(n_353), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_250), .Y(n_116) );
OAI21xp33_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_186), .B(n_217), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_118), .A2(n_465), .B(n_467), .Y(n_464) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OR2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_146), .Y(n_119) );
OR2x2_ASAP7_75t_L g392 ( .A(n_120), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_120), .B(n_425), .Y(n_424) );
INVx2_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g273 ( .A(n_122), .Y(n_273) );
INVx2_ASAP7_75t_L g304 ( .A(n_122), .Y(n_304) );
AND2x2_ASAP7_75t_L g325 ( .A(n_122), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g444 ( .A(n_122), .B(n_148), .Y(n_444) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_144), .Y(n_122) );
AND2x2_ASAP7_75t_L g345 ( .A(n_123), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_136), .Y(n_123) );
AOI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_129), .B1(n_131), .B2(n_135), .Y(n_124) );
AOI22xp5_ASAP7_75t_L g158 ( .A1(n_126), .A2(n_159), .B1(n_160), .B2(n_161), .Y(n_158) );
INVx1_ASAP7_75t_L g177 ( .A(n_126), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_126), .A2(n_128), .B1(n_247), .B2(n_248), .Y(n_246) );
INVx2_ASAP7_75t_L g530 ( .A(n_126), .Y(n_530) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_126), .Y(n_601) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g134 ( .A(n_127), .Y(n_134) );
INVx6_ASAP7_75t_L g155 ( .A(n_127), .Y(n_155) );
INVx3_ASAP7_75t_L g194 ( .A(n_127), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_128), .A2(n_155), .B1(n_156), .B2(n_157), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_128), .B(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_128), .B(n_202), .Y(n_201) );
AOI22xp33_ASAP7_75t_SL g243 ( .A1(n_128), .A2(n_155), .B1(n_244), .B2(n_245), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_128), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g529 ( .A(n_128), .Y(n_529) );
INVx2_ASAP7_75t_L g537 ( .A(n_128), .Y(n_537) );
INVx2_ASAP7_75t_L g550 ( .A(n_128), .Y(n_550) );
INVx1_ASAP7_75t_L g567 ( .A(n_128), .Y(n_567) );
INVx2_ASAP7_75t_L g581 ( .A(n_128), .Y(n_581) );
NAND2xp33_ASAP7_75t_L g595 ( .A(n_128), .B(n_596), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g153 ( .A1(n_129), .A2(n_135), .B1(n_154), .B2(n_158), .Y(n_153) );
INVx1_ASAP7_75t_L g216 ( .A(n_129), .Y(n_216) );
OAI221xp5_ASAP7_75t_L g242 ( .A1(n_129), .A2(n_138), .B1(n_180), .B2(n_243), .C(n_246), .Y(n_242) );
INVx2_ASAP7_75t_SL g586 ( .A(n_129), .Y(n_586) );
INVx1_ASAP7_75t_L g598 ( .A(n_129), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_129), .B(n_674), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_129), .B(n_678), .Y(n_677) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx4_ASAP7_75t_L g135 ( .A(n_130), .Y(n_135) );
INVx3_ASAP7_75t_L g180 ( .A(n_130), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_130), .B(n_200), .Y(n_199) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_130), .Y(n_224) );
INVx1_ASAP7_75t_L g228 ( .A(n_130), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_130), .B(n_236), .Y(n_235) );
INVxp67_ASAP7_75t_L g584 ( .A(n_130), .Y(n_584) );
INVx2_ASAP7_75t_L g171 ( .A(n_132), .Y(n_171) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g160 ( .A(n_133), .Y(n_160) );
INVx2_ASAP7_75t_L g569 ( .A(n_134), .Y(n_569) );
INVx1_ASAP7_75t_L g669 ( .A(n_134), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g197 ( .A1(n_135), .A2(n_198), .B1(n_199), .B2(n_201), .Y(n_197) );
INVx2_ASAP7_75t_L g213 ( .A(n_135), .Y(n_213) );
O2A1O1Ixp5_ASAP7_75t_SL g663 ( .A1(n_135), .A2(n_664), .B(n_665), .C(n_668), .Y(n_663) );
NOR2xp67_ASAP7_75t_L g136 ( .A(n_137), .B(n_140), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_137), .B(n_291), .Y(n_631) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_138), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_138), .B(n_166), .Y(n_239) );
AND2x2_ASAP7_75t_L g538 ( .A(n_138), .B(n_290), .Y(n_538) );
INVx3_ASAP7_75t_L g555 ( .A(n_138), .Y(n_555) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx3_ASAP7_75t_L g203 ( .A(n_141), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_141), .B(n_268), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_141), .B(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx4_ASAP7_75t_L g166 ( .A(n_142), .Y(n_166) );
BUFx3_ASAP7_75t_L g291 ( .A(n_142), .Y(n_291) );
BUFx3_ASAP7_75t_L g152 ( .A(n_145), .Y(n_152) );
INVx1_ASAP7_75t_L g206 ( .A(n_145), .Y(n_206) );
INVx1_ASAP7_75t_L g258 ( .A(n_145), .Y(n_258) );
INVx2_ASAP7_75t_L g348 ( .A(n_145), .Y(n_348) );
INVx1_ASAP7_75t_L g563 ( .A(n_145), .Y(n_563) );
INVx2_ASAP7_75t_SL g146 ( .A(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_147), .B(n_277), .Y(n_397) );
AND2x2_ASAP7_75t_L g484 ( .A(n_147), .B(n_428), .Y(n_484) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_167), .Y(n_147) );
INVx1_ASAP7_75t_L g301 ( .A(n_148), .Y(n_301) );
OAI21x1_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_153), .B(n_162), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_150), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_150), .B(n_290), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_151), .B(n_183), .Y(n_222) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g214 ( .A(n_154), .Y(n_214) );
INVx2_ASAP7_75t_L g173 ( .A(n_155), .Y(n_173) );
INVx2_ASAP7_75t_SL g227 ( .A(n_155), .Y(n_227) );
INVx1_ASAP7_75t_L g614 ( .A(n_155), .Y(n_614) );
INVx2_ASAP7_75t_L g623 ( .A(n_155), .Y(n_623) );
INVx1_ASAP7_75t_L g667 ( .A(n_155), .Y(n_667) );
INVx1_ASAP7_75t_L g215 ( .A(n_158), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_160), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_160), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g536 ( .A(n_160), .Y(n_536) );
INVx2_ASAP7_75t_L g551 ( .A(n_160), .Y(n_551) );
OR2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
INVx2_ASAP7_75t_L g241 ( .A(n_164), .Y(n_241) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_SL g181 ( .A(n_165), .B(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_SL g184 ( .A(n_166), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g210 ( .A(n_166), .Y(n_210) );
OR2x2_ASAP7_75t_L g207 ( .A(n_167), .B(n_208), .Y(n_207) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_167), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_167), .B(n_190), .Y(n_282) );
INVx2_ASAP7_75t_L g303 ( .A(n_167), .Y(n_303) );
INVx1_ASAP7_75t_L g342 ( .A(n_167), .Y(n_342) );
INVx1_ASAP7_75t_L g383 ( .A(n_167), .Y(n_383) );
AND2x2_ASAP7_75t_L g418 ( .A(n_167), .B(n_208), .Y(n_418) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_167), .Y(n_473) );
AO31x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_175), .A3(n_181), .B(n_184), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx3_ASAP7_75t_L g544 ( .A(n_171), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_173), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_177), .A2(n_628), .B1(n_629), .B2(n_630), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_180), .A2(n_238), .B(n_239), .Y(n_237) );
INVx3_ASAP7_75t_L g531 ( .A(n_180), .Y(n_531) );
NOR3xp33_ASAP7_75t_L g191 ( .A(n_182), .B(n_192), .C(n_197), .Y(n_191) );
AOI221xp5_ASAP7_75t_L g212 ( .A1(n_182), .A2(n_213), .B1(n_214), .B2(n_215), .C(n_216), .Y(n_212) );
NOR4xp25_ASAP7_75t_L g564 ( .A(n_182), .B(n_565), .C(n_571), .D(n_574), .Y(n_564) );
NOR2x1_ASAP7_75t_SL g592 ( .A(n_182), .B(n_241), .Y(n_592) );
INVx4_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g257 ( .A(n_183), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
OR2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_207), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g272 ( .A(n_190), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g311 ( .A(n_190), .B(n_303), .Y(n_311) );
INVx2_ASAP7_75t_L g326 ( .A(n_190), .Y(n_326) );
INVx2_ASAP7_75t_L g352 ( .A(n_190), .Y(n_352) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_203), .B(n_204), .Y(n_190) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g198 ( .A(n_194), .Y(n_198) );
INVx1_ASAP7_75t_L g264 ( .A(n_194), .Y(n_264) );
INVx2_ASAP7_75t_L g546 ( .A(n_194), .Y(n_546) );
INVx2_ASAP7_75t_L g582 ( .A(n_194), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_203), .B(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g680 ( .A(n_203), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_207), .Y(n_308) );
OR2x2_ASAP7_75t_L g323 ( .A(n_207), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g400 ( .A(n_207), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_208), .B(n_352), .Y(n_351) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_208), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_208), .B(n_408), .Y(n_434) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_211), .Y(n_208) );
INVx2_ASAP7_75t_L g553 ( .A(n_210), .Y(n_553) );
AND2x2_ASAP7_75t_L g344 ( .A(n_211), .B(n_345), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_213), .A2(n_260), .B(n_263), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_213), .A2(n_610), .B(n_611), .Y(n_609) );
AOI322xp5_ASAP7_75t_L g426 ( .A1(n_217), .A2(n_366), .A3(n_404), .B1(n_427), .B2(n_429), .C1(n_430), .C2(n_431), .Y(n_426) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_230), .Y(n_217) );
AND2x2_ASAP7_75t_L g431 ( .A(n_218), .B(n_411), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_218), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g482 ( .A(n_218), .B(n_374), .Y(n_482) );
INVx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_219), .B(n_279), .Y(n_297) );
AND2x2_ASAP7_75t_L g358 ( .A(n_219), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_219), .B(n_320), .Y(n_402) );
AND2x4_ASAP7_75t_L g439 ( .A(n_219), .B(n_230), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_219), .B(n_361), .Y(n_480) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g269 ( .A(n_220), .B(n_240), .Y(n_269) );
INVx1_ASAP7_75t_L g318 ( .A(n_220), .Y(n_318) );
AND2x2_ASAP7_75t_L g462 ( .A(n_220), .B(n_295), .Y(n_462) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g280 ( .A(n_221), .Y(n_280) );
OAI21x1_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_229), .Y(n_221) );
INVx1_ASAP7_75t_L g289 ( .A(n_223), .Y(n_289) );
OA22x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B1(n_226), .B2(n_228), .Y(n_223) );
INVx4_ASAP7_75t_L g533 ( .A(n_224), .Y(n_533) );
INVx1_ASAP7_75t_L g292 ( .A(n_229), .Y(n_292) );
INVx1_ASAP7_75t_SL g387 ( .A(n_230), .Y(n_387) );
AND2x4_ASAP7_75t_L g230 ( .A(n_231), .B(n_240), .Y(n_230) );
AND2x2_ASAP7_75t_L g279 ( .A(n_231), .B(n_255), .Y(n_279) );
INVx1_ASAP7_75t_L g320 ( .A(n_231), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_231), .B(n_254), .Y(n_496) );
INVx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g295 ( .A(n_232), .Y(n_295) );
INVx1_ASAP7_75t_L g337 ( .A(n_232), .Y(n_337) );
AND2x2_ASAP7_75t_L g361 ( .A(n_232), .B(n_240), .Y(n_361) );
AND2x2_ASAP7_75t_L g411 ( .A(n_232), .B(n_255), .Y(n_411) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_232), .Y(n_415) );
AND2x4_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
OR2x2_ASAP7_75t_L g287 ( .A(n_240), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g317 ( .A(n_240), .B(n_318), .Y(n_317) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_249), .Y(n_240) );
OA21x2_ASAP7_75t_L g332 ( .A1(n_241), .A2(n_242), .B(n_249), .Y(n_332) );
AOI221xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_270), .B1(n_277), .B2(n_281), .C(n_283), .Y(n_250) );
INVxp67_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_269), .Y(n_252) );
AND2x2_ASAP7_75t_L g457 ( .A(n_253), .B(n_317), .Y(n_457) );
BUFx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g471 ( .A(n_254), .B(n_352), .Y(n_471) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g294 ( .A(n_255), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g315 ( .A(n_255), .Y(n_315) );
AND2x2_ASAP7_75t_L g338 ( .A(n_255), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g360 ( .A(n_255), .Y(n_360) );
BUFx2_ASAP7_75t_L g448 ( .A(n_255), .Y(n_448) );
INVx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AOI21x1_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_259), .B(n_267), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_269), .A2(n_293), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g460 ( .A(n_269), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_270), .A2(n_307), .B1(n_312), .B2(n_319), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_274), .Y(n_270) );
OR2x2_ASAP7_75t_L g368 ( .A(n_271), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
AND2x4_ASAP7_75t_L g399 ( .A(n_272), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g417 ( .A(n_272), .B(n_418), .Y(n_417) );
INVxp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g491 ( .A(n_276), .B(n_407), .Y(n_491) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_SL g403 ( .A(n_278), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g379 ( .A(n_280), .B(n_360), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_280), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g466 ( .A(n_280), .Y(n_466) );
OR2x2_ASAP7_75t_L g495 ( .A(n_280), .B(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_L g463 ( .A(n_281), .B(n_444), .Y(n_463) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AOI21xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_296), .B(n_298), .Y(n_283) );
INVx2_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_293), .Y(n_285) );
AND2x2_ASAP7_75t_L g319 ( .A(n_286), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g421 ( .A(n_286), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g330 ( .A(n_288), .B(n_331), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_290), .B(n_292), .Y(n_288) );
INVx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g374 ( .A(n_295), .B(n_331), .Y(n_374) );
OAI21xp33_ASAP7_75t_L g492 ( .A1(n_296), .A2(n_381), .B(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_302), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g474 ( .A(n_300), .B(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g349 ( .A(n_302), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g433 ( .A(n_302), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g370 ( .A(n_303), .Y(n_370) );
INVx1_ASAP7_75t_L g409 ( .A(n_304), .Y(n_409) );
AND2x4_ASAP7_75t_L g428 ( .A(n_304), .B(n_352), .Y(n_428) );
INVx1_ASAP7_75t_SL g475 ( .A(n_304), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_321), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g443 ( .A(n_311), .B(n_444), .Y(n_443) );
NOR2x1_ASAP7_75t_L g312 ( .A(n_313), .B(n_316), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g328 ( .A(n_314), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g427 ( .A(n_314), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_315), .B(n_339), .Y(n_489) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_319), .B(n_340), .Y(n_375) );
AND2x2_ASAP7_75t_L g366 ( .A(n_320), .B(n_330), .Y(n_366) );
AOI222xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_327), .B1(n_333), .B2(n_335), .C1(n_340), .C2(n_349), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OAI21xp33_ASAP7_75t_L g372 ( .A1(n_323), .A2(n_373), .B(n_375), .Y(n_372) );
OAI221xp5_ASAP7_75t_L g440 ( .A1(n_323), .A2(n_441), .B1(n_442), .B2(n_445), .C(n_449), .Y(n_440) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx2_ASAP7_75t_L g355 ( .A(n_325), .Y(n_355) );
AND2x2_ASAP7_75t_L g384 ( .A(n_326), .B(n_344), .Y(n_384) );
INVx1_ASAP7_75t_L g408 ( .A(n_326), .Y(n_408) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_326), .Y(n_437) );
OAI21xp5_ASAP7_75t_L g420 ( .A1(n_327), .A2(n_421), .B(n_423), .Y(n_420) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g451 ( .A(n_330), .B(n_422), .Y(n_451) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g339 ( .A(n_332), .Y(n_339) );
INVxp67_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_338), .Y(n_365) );
INVx2_ASAP7_75t_L g416 ( .A(n_339), .Y(n_416) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
OR2x2_ASAP7_75t_L g472 ( .A(n_343), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g438 ( .A(n_344), .Y(n_438) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_348), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g574 ( .A(n_348), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_349), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g393 ( .A(n_351), .B(n_370), .Y(n_393) );
NAND4xp25_ASAP7_75t_L g353 ( .A(n_354), .B(n_362), .C(n_371), .D(n_376), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
A2O1A1Ixp33_ASAP7_75t_L g449 ( .A1(n_355), .A2(n_450), .B(n_451), .C(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g390 ( .A(n_360), .Y(n_390) );
INVx1_ASAP7_75t_L g422 ( .A(n_360), .Y(n_422) );
OAI21xp5_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_366), .B(n_367), .Y(n_362) );
INVxp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVxp33_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2x1p5_ASAP7_75t_L g453 ( .A(n_374), .B(n_448), .Y(n_453) );
AND2x4_ASAP7_75t_L g465 ( .A(n_374), .B(n_466), .Y(n_465) );
NAND2x1p5_ASAP7_75t_L g476 ( .A(n_374), .B(n_389), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_380), .B1(n_385), .B2(n_391), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2x1p5_ASAP7_75t_SL g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVx2_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g450 ( .A(n_383), .Y(n_450) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_384), .Y(n_430) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
OR2x2_ASAP7_75t_L g441 ( .A(n_388), .B(n_414), .Y(n_441) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g429 ( .A(n_393), .Y(n_429) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_454), .Y(n_394) );
NOR3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_419), .C(n_440), .Y(n_395) );
NAND3xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .C(n_410), .Y(n_396) );
AOI22x1_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B1(n_403), .B2(n_405), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
OAI21xp33_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_412), .B(n_417), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_416), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g488 ( .A(n_415), .Y(n_488) );
INVx1_ASAP7_75t_L g468 ( .A(n_416), .Y(n_468) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_418), .Y(n_425) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_426), .C(n_432), .Y(n_419) );
INVx1_ASAP7_75t_L g461 ( .A(n_422), .Y(n_461) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_435), .B(n_439), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_433), .A2(n_451), .B1(n_486), .B2(n_490), .Y(n_485) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVxp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NOR3xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_477), .C(n_492), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_464), .Y(n_455) );
OAI31xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .A3(n_462), .B(n_463), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B1(n_474), .B2(n_476), .Y(n_467) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NOR2x1_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_481), .B(n_483), .C(n_485), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
BUFx12f_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx10_ASAP7_75t_L g512 ( .A(n_502), .Y(n_512) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
OR2x6_ASAP7_75t_L g888 ( .A(n_505), .B(n_889), .Y(n_888) );
INVx8_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g891 ( .A(n_506), .B(n_892), .Y(n_891) );
OR2x6_ASAP7_75t_L g909 ( .A(n_506), .B(n_892), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_510), .A2(n_514), .B(n_910), .Y(n_513) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_893), .B1(n_899), .B2(n_903), .C(n_904), .Y(n_514) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_800), .Y(n_517) );
NAND3xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_720), .C(n_764), .Y(n_518) );
NOR3xp33_ASAP7_75t_L g519 ( .A(n_520), .B(n_690), .C(n_708), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_644), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_588), .B1(n_633), .B2(n_641), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g776 ( .A(n_523), .Y(n_776) );
OR2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_558), .Y(n_523) );
NOR2x1p5_ASAP7_75t_L g791 ( .A(n_524), .B(n_696), .Y(n_791) );
NAND2x1_ASAP7_75t_L g524 ( .A(n_525), .B(n_540), .Y(n_524) );
INVx2_ASAP7_75t_L g636 ( .A(n_525), .Y(n_636) );
INVx2_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g700 ( .A(n_526), .Y(n_700) );
AO31x2_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_532), .A3(n_538), .B(n_539), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_531), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_531), .A2(n_548), .B(n_552), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_533), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g672 ( .A(n_537), .Y(n_672) );
NOR2x1_ASAP7_75t_L g701 ( .A(n_540), .B(n_650), .Y(n_701) );
INVx1_ASAP7_75t_L g751 ( .A(n_540), .Y(n_751) );
AND2x2_ASAP7_75t_L g811 ( .A(n_540), .B(n_638), .Y(n_811) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g649 ( .A(n_541), .Y(n_649) );
AOI21x1_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_547), .B(n_556), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_544), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
AOI21x1_ASAP7_75t_L g638 ( .A1(n_553), .A2(n_639), .B(n_640), .Y(n_638) );
OAI21x1_ASAP7_75t_L g608 ( .A1(n_554), .A2(n_609), .B(n_612), .Y(n_608) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OAI21x1_ASAP7_75t_L g679 ( .A1(n_555), .A2(n_675), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g768 ( .A(n_559), .B(n_699), .Y(n_768) );
NOR2x1_ASAP7_75t_L g559 ( .A(n_560), .B(n_575), .Y(n_559) );
AND2x2_ASAP7_75t_L g724 ( .A(n_560), .B(n_700), .Y(n_724) );
INVx1_ASAP7_75t_L g790 ( .A(n_560), .Y(n_790) );
AND2x4_ASAP7_75t_L g798 ( .A(n_560), .B(n_636), .Y(n_798) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_560), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_560), .B(n_853), .Y(n_852) );
OR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_564), .Y(n_560) );
INVxp67_ASAP7_75t_SL g656 ( .A(n_561), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVx1_ASAP7_75t_L g577 ( .A(n_563), .Y(n_577) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_569), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g628 ( .A(n_569), .Y(n_628) );
INVxp67_ASAP7_75t_SL g655 ( .A(n_571), .Y(n_655) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_576), .Y(n_696) );
AND2x2_ASAP7_75t_L g719 ( .A(n_576), .B(n_648), .Y(n_719) );
INVx1_ASAP7_75t_L g847 ( .A(n_576), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_576), .B(n_700), .Y(n_850) );
OA21x2_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B(n_587), .Y(n_576) );
OAI21x1_ASAP7_75t_L g607 ( .A1(n_577), .A2(n_608), .B(n_616), .Y(n_607) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_579), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_583), .B1(n_585), .B2(n_586), .Y(n_579) );
OAI21xp5_ASAP7_75t_SL g626 ( .A1(n_583), .A2(n_627), .B(n_631), .Y(n_626) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g640 ( .A(n_587), .Y(n_640) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_606), .Y(n_588) );
OR2x6_ASAP7_75t_L g706 ( .A(n_589), .B(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g818 ( .A(n_589), .B(n_728), .Y(n_818) );
INVx2_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g759 ( .A(n_590), .B(n_760), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_590), .B(n_787), .Y(n_786) );
AND2x4_ASAP7_75t_L g807 ( .A(n_590), .B(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g642 ( .A(n_591), .Y(n_642) );
OR2x2_ASAP7_75t_L g660 ( .A(n_591), .B(n_661), .Y(n_660) );
OR2x2_ASAP7_75t_L g714 ( .A(n_591), .B(n_715), .Y(n_714) );
AND2x4_ASAP7_75t_L g733 ( .A(n_591), .B(n_661), .Y(n_733) );
AND2x2_ASAP7_75t_L g783 ( .A(n_591), .B(n_715), .Y(n_783) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_591), .Y(n_861) );
AO31x2_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .A3(n_599), .B(n_604), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_597), .B(n_598), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_598), .A2(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_617), .Y(n_606) );
AND2x2_ASAP7_75t_L g643 ( .A(n_607), .B(n_618), .Y(n_643) );
OR2x2_ASAP7_75t_L g766 ( .A(n_607), .B(n_714), .Y(n_766) );
AND2x2_ASAP7_75t_L g808 ( .A(n_607), .B(n_662), .Y(n_808) );
OAI21x1_ASAP7_75t_L g684 ( .A1(n_608), .A2(n_616), .B(n_680), .Y(n_684) );
AND2x2_ASAP7_75t_L g682 ( .A(n_617), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g858 ( .A(n_617), .B(n_642), .Y(n_858) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_618), .B(n_737), .Y(n_736) );
INVx3_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g689 ( .A(n_619), .Y(n_689) );
INVx1_ASAP7_75t_L g747 ( .A(n_619), .Y(n_747) );
OA21x2_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_626), .B(n_632), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g869 ( .A(n_634), .B(n_701), .Y(n_869) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
BUFx2_ASAP7_75t_SL g646 ( .A(n_636), .Y(n_646) );
INVx1_ASAP7_75t_L g712 ( .A(n_636), .Y(n_712) );
AND2x2_ASAP7_75t_L g752 ( .A(n_636), .B(n_650), .Y(n_752) );
AND2x2_ASAP7_75t_L g774 ( .A(n_637), .B(n_763), .Y(n_774) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g754 ( .A(n_638), .B(n_648), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_641), .B(n_793), .Y(n_792) );
INVxp33_ASAP7_75t_L g799 ( .A(n_641), .Y(n_799) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
INVx1_ASAP7_75t_L g737 ( .A(n_642), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_642), .Y(n_740) );
OR2x2_ASAP7_75t_L g819 ( .A(n_642), .B(n_820), .Y(n_819) );
AND2x2_ASAP7_75t_L g868 ( .A(n_642), .B(n_687), .Y(n_868) );
INVx1_ASAP7_75t_L g760 ( .A(n_643), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_657), .Y(n_644) );
INVx1_ASAP7_75t_L g729 ( .A(n_645), .Y(n_729) );
AND2x4_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
NAND2x1p5_ASAP7_75t_L g743 ( .A(n_647), .B(n_696), .Y(n_743) );
INVx3_ASAP7_75t_L g845 ( .A(n_647), .Y(n_845) );
AND2x4_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g763 ( .A(n_649), .Y(n_763) );
INVxp67_ASAP7_75t_SL g886 ( .A(n_650), .Y(n_886) );
OA21x2_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B(n_656), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI21xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_681), .B(n_685), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g834 ( .A(n_660), .Y(n_834) );
OR2x2_ASAP7_75t_L g865 ( .A(n_660), .B(n_837), .Y(n_865) );
AND2x2_ASAP7_75t_L g688 ( .A(n_661), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_661), .B(n_687), .Y(n_728) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g821 ( .A(n_662), .B(n_683), .Y(n_821) );
OAI21x1_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_670), .B(n_679), .Y(n_662) );
OAI21xp5_ASAP7_75t_L g715 ( .A1(n_663), .A2(n_670), .B(n_679), .Y(n_715) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_666), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND3x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_675), .C(n_676), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g758 ( .A(n_682), .B(n_733), .Y(n_758) );
INVxp67_ASAP7_75t_L g771 ( .A(n_682), .Y(n_771) );
INVx2_ASAP7_75t_L g687 ( .A(n_683), .Y(n_687) );
AND2x2_ASAP7_75t_L g741 ( .A(n_683), .B(n_689), .Y(n_741) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g777 ( .A(n_685), .Y(n_777) );
NAND2x1p5_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
INVx2_ASAP7_75t_L g787 ( .A(n_686), .Y(n_787) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
BUFx2_ASAP7_75t_SL g707 ( .A(n_687), .Y(n_707) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_687), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_688), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g755 ( .A(n_688), .Y(n_755) );
INVx2_ASAP7_75t_SL g705 ( .A(n_689), .Y(n_705) );
BUFx2_ASAP7_75t_L g810 ( .A(n_689), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_702), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x4_ASAP7_75t_L g692 ( .A(n_693), .B(n_697), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_695), .B(n_699), .Y(n_779) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g842 ( .A(n_696), .Y(n_842) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_701), .Y(n_698) );
BUFx3_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
NOR2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_706), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g713 ( .A(n_705), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g782 ( .A(n_705), .Y(n_782) );
AND2x2_ASAP7_75t_L g862 ( .A(n_705), .B(n_821), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_705), .B(n_783), .Y(n_866) );
NOR3xp33_ASAP7_75t_L g885 ( .A(n_705), .B(n_711), .C(n_886), .Y(n_885) );
AND2x2_ASAP7_75t_L g824 ( .A(n_706), .B(n_770), .Y(n_824) );
INVx1_ASAP7_75t_L g732 ( .A(n_707), .Y(n_732) );
O2A1O1Ixp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_713), .B(n_716), .C(n_718), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND2x1p5_ASAP7_75t_L g828 ( .A(n_711), .B(n_829), .Y(n_828) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
OR2x2_ASAP7_75t_L g753 ( .A(n_712), .B(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g773 ( .A(n_712), .B(n_774), .Y(n_773) );
OR2x2_ASAP7_75t_L g796 ( .A(n_714), .B(n_782), .Y(n_796) );
INVx1_ASAP7_75t_L g874 ( .A(n_714), .Y(n_874) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_715), .Y(n_770) );
OAI221xp5_ASAP7_75t_L g856 ( .A1(n_718), .A2(n_828), .B1(n_857), .B2(n_859), .C(n_863), .Y(n_856) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g723 ( .A(n_719), .B(n_724), .Y(n_723) );
NOR4xp25_ASAP7_75t_L g720 ( .A(n_721), .B(n_734), .C(n_744), .D(n_756), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_725), .B1(n_729), .B2(n_730), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_722), .A2(n_735), .B1(n_738), .B2(n_742), .Y(n_734) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AOI21xp33_ASAP7_75t_SL g803 ( .A1(n_723), .A2(n_804), .B(n_805), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_724), .B(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g780 ( .A(n_724), .Y(n_780) );
AND2x2_ASAP7_75t_L g841 ( .A(n_724), .B(n_842), .Y(n_841) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g836 ( .A(n_727), .B(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI211xp5_ASAP7_75t_L g838 ( .A1(n_730), .A2(n_839), .B(n_840), .C(n_843), .Y(n_838) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_733), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g814 ( .A(n_733), .B(n_787), .Y(n_814) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_741), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AND2x4_ASAP7_75t_L g854 ( .A(n_740), .B(n_808), .Y(n_854) );
INVx1_ASAP7_75t_L g879 ( .A(n_741), .Y(n_879) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g829 ( .A(n_743), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_748), .B1(n_753), .B2(n_755), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_746), .B(n_877), .Y(n_876) );
BUFx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_R g837 ( .A(n_747), .Y(n_837) );
OAI22xp33_ASAP7_75t_L g795 ( .A1(n_748), .A2(n_796), .B1(n_797), .B2(n_799), .Y(n_795) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_752), .Y(n_749) );
NOR2xp33_ASAP7_75t_SL g887 ( .A(n_750), .B(n_846), .Y(n_887) );
INVxp67_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AND2x2_ASAP7_75t_L g881 ( .A(n_751), .B(n_768), .Y(n_881) );
AND2x4_ASAP7_75t_L g826 ( .A(n_752), .B(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g871 ( .A(n_753), .Y(n_871) );
INVx2_ASAP7_75t_L g827 ( .A(n_754), .Y(n_827) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_759), .B(n_761), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OAI221xp5_ASAP7_75t_L g823 ( .A1(n_759), .A2(n_824), .B1(n_825), .B2(n_828), .C(n_830), .Y(n_823) );
AND2x2_ASAP7_75t_L g835 ( .A(n_762), .B(n_790), .Y(n_835) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_763), .Y(n_816) );
INVx1_ASAP7_75t_L g853 ( .A(n_763), .Y(n_853) );
NOR3xp33_ASAP7_75t_L g764 ( .A(n_765), .B(n_784), .C(n_795), .Y(n_764) );
OAI221xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_767), .B1(n_769), .B2(n_772), .C(n_775), .Y(n_765) );
INVx1_ASAP7_75t_L g870 ( .A(n_766), .Y(n_870) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
OR2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g880 ( .A1(n_770), .A2(n_881), .B1(n_882), .B2(n_883), .Y(n_880) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_774), .B(n_789), .Y(n_794) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_777), .B1(n_778), .B2(n_781), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
AND2x2_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
NAND2xp5_ASAP7_75t_SL g784 ( .A(n_785), .B(n_792), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_788), .Y(n_785) );
AND2x2_ASAP7_75t_L g788 ( .A(n_789), .B(n_791), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_791), .Y(n_831) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx2_ASAP7_75t_L g804 ( .A(n_796), .Y(n_804) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AND2x2_ASAP7_75t_L g815 ( .A(n_798), .B(n_816), .Y(n_815) );
AND2x4_ASAP7_75t_L g822 ( .A(n_798), .B(n_811), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_801), .B(n_855), .Y(n_800) );
NOR3xp33_ASAP7_75t_L g801 ( .A(n_802), .B(n_823), .C(n_838), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_813), .Y(n_802) );
NOR3xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_809), .C(n_812), .Y(n_805) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
OAI21xp33_ASAP7_75t_L g840 ( .A1(n_807), .A2(n_815), .B(n_841), .Y(n_840) );
AND2x2_ASAP7_75t_L g882 ( .A(n_808), .B(n_837), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
INVx1_ASAP7_75t_L g833 ( .A(n_810), .Y(n_833) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_815), .B1(n_817), .B2(n_822), .Y(n_813) );
NAND2xp5_ASAP7_75t_SL g817 ( .A(n_818), .B(n_819), .Y(n_817) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_826), .A2(n_874), .B1(n_875), .B2(n_878), .Y(n_873) );
AOI22xp33_ASAP7_75t_SL g830 ( .A1(n_831), .A2(n_832), .B1(n_835), .B2(n_836), .Y(n_830) );
INVx1_ASAP7_75t_L g839 ( .A(n_831), .Y(n_839) );
AND2x2_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
OAI21xp5_ASAP7_75t_SL g843 ( .A1(n_844), .A2(n_848), .B(n_854), .Y(n_843) );
NOR2x1_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
AND2x2_ASAP7_75t_L g848 ( .A(n_849), .B(n_851), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
NOR2xp33_ASAP7_75t_L g877 ( .A(n_850), .B(n_852), .Y(n_877) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_872), .Y(n_855) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
AND2x2_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .Y(n_860) );
AOI22xp33_ASAP7_75t_SL g863 ( .A1(n_864), .A2(n_869), .B1(n_870), .B2(n_871), .Y(n_863) );
NAND3xp33_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .C(n_867), .Y(n_864) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_873), .B(n_880), .Y(n_872) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_885), .B(n_887), .Y(n_884) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_888), .Y(n_900) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
BUFx8_ASAP7_75t_L g902 ( .A(n_891), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_893), .Y(n_903) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
BUFx2_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
NOR2xp33_ASAP7_75t_L g904 ( .A(n_905), .B(n_906), .Y(n_904) );
BUFx2_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
BUFx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
BUFx3_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
CKINVDCx20_ASAP7_75t_R g910 ( .A(n_911), .Y(n_910) );
CKINVDCx20_ASAP7_75t_R g911 ( .A(n_912), .Y(n_911) );
CKINVDCx20_ASAP7_75t_R g912 ( .A(n_913), .Y(n_912) );
CKINVDCx5p33_ASAP7_75t_R g914 ( .A(n_915), .Y(n_914) );
BUFx24_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
BUFx2_ASAP7_75t_L g926 ( .A(n_916), .Y(n_926) );
OR2x2_ASAP7_75t_SL g916 ( .A(n_917), .B(n_923), .Y(n_916) );
NAND3xp33_ASAP7_75t_L g917 ( .A(n_918), .B(n_919), .C(n_921), .Y(n_917) );
CKINVDCx5p33_ASAP7_75t_R g919 ( .A(n_920), .Y(n_919) );
CKINVDCx5p33_ASAP7_75t_R g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
endmodule