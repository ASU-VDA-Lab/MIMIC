module fake_jpeg_5332_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

HAxp5_ASAP7_75t_SL g33 ( 
.A(n_32),
.B(n_0),
.CON(n_33),
.SN(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_39),
.Y(n_47)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_28),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_23),
.B1(n_30),
.B2(n_32),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_52),
.B1(n_34),
.B2(n_16),
.Y(n_62)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_44),
.Y(n_79)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_29),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_35),
.Y(n_63)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_53),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_23),
.B1(n_30),
.B2(n_29),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_26),
.B1(n_24),
.B2(n_17),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_23),
.B1(n_32),
.B2(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_36),
.B1(n_35),
.B2(n_21),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_57),
.A2(n_65),
.B1(n_81),
.B2(n_16),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_40),
.C(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_60),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_54),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_63),
.B(n_73),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_77),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_55),
.A2(n_36),
.B1(n_17),
.B2(n_24),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_75),
.Y(n_98)
);

BUFx2_ASAP7_75t_SL g67 ( 
.A(n_45),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_67),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_80),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_32),
.B(n_39),
.C(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_72),
.Y(n_99)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_76),
.Y(n_104)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_41),
.B(n_26),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_82),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_28),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_28),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_86),
.Y(n_108)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_100),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_95),
.Y(n_116)
);

BUFx4f_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_45),
.Y(n_95)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_SL g119 ( 
.A1(n_101),
.A2(n_77),
.B(n_66),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_1),
.B(n_2),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_27),
.B(n_25),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_44),
.B1(n_16),
.B2(n_38),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_72),
.B1(n_78),
.B2(n_39),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_27),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_38),
.Y(n_128)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_85),
.Y(n_124)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_111),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_63),
.B(n_44),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_82),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_80),
.C(n_68),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_122),
.C(n_87),
.Y(n_140)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_121),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_73),
.B1(n_59),
.B2(n_62),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_117),
.A2(n_132),
.B1(n_137),
.B2(n_100),
.Y(n_143)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_59),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_118),
.A2(n_31),
.B(n_22),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_119),
.A2(n_127),
.B1(n_133),
.B2(n_22),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_71),
.B(n_68),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_120),
.A2(n_31),
.B(n_22),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_39),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_124),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_86),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_128),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_31),
.Y(n_129)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_138),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_98),
.B(n_15),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_131),
.B(n_134),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_104),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_96),
.A2(n_39),
.B1(n_38),
.B2(n_61),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_31),
.Y(n_136)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_111),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_88),
.B(n_92),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_139),
.A2(n_141),
.B(n_148),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_144),
.C(n_153),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_93),
.B(n_99),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_147),
.B1(n_149),
.B2(n_151),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_101),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_113),
.A2(n_106),
.B1(n_110),
.B2(n_97),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_90),
.B(n_103),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_106),
.B(n_90),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_113),
.A2(n_106),
.B1(n_94),
.B2(n_56),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_116),
.A2(n_114),
.B1(n_138),
.B2(n_130),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_152),
.A2(n_131),
.B1(n_135),
.B2(n_137),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_39),
.C(n_94),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_157),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_27),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_25),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_160),
.Y(n_176)
);

AND2x4_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_94),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_149),
.C(n_141),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_132),
.B(n_15),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_164),
.Y(n_167)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_113),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_20),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_142),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_159),
.A2(n_133),
.B1(n_123),
.B2(n_126),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_181),
.B1(n_182),
.B2(n_161),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_134),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_177),
.C(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_146),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_178),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_127),
.C(n_115),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_159),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g197 ( 
.A(n_179),
.B(n_165),
.CI(n_163),
.CON(n_197),
.SN(n_197)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_144),
.C(n_157),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_159),
.A2(n_135),
.B1(n_91),
.B2(n_22),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_91),
.C(n_20),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_155),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g187 ( 
.A(n_164),
.Y(n_187)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_139),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_193),
.C(n_194),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_181),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_189),
.B(n_204),
.Y(n_216)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_148),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_158),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_202),
.C(n_180),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_199),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_161),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_185),
.B(n_169),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_184),
.B1(n_178),
.B2(n_170),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_188),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_198),
.A2(n_185),
.B1(n_172),
.B2(n_179),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_208),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_203),
.B(n_145),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_204),
.A2(n_183),
.B1(n_177),
.B2(n_169),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_209),
.B(n_196),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_217),
.C(n_200),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_191),
.A2(n_142),
.B1(n_176),
.B2(n_162),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_197),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_215),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_176),
.B1(n_162),
.B2(n_160),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_195),
.B(n_2),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_2),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_215),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_220),
.C(n_221),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_200),
.C(n_202),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_222),
.B(n_226),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_225),
.C(n_227),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_91),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_20),
.C(n_5),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_20),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_218),
.C(n_213),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_216),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_237),
.Y(n_242)
);

BUFx4f_ASAP7_75t_SL g231 ( 
.A(n_219),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_231),
.B(n_236),
.Y(n_240)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_222),
.B(n_211),
.Y(n_234)
);

NOR2xp67_ASAP7_75t_SL g244 ( 
.A(n_234),
.B(n_8),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_212),
.Y(n_236)
);

NOR2x1p5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_229),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_239),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_206),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_3),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_241),
.B(n_243),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_232),
.A2(n_3),
.B1(n_5),
.B2(n_8),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_8),
.C(n_9),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_244),
.Y(n_247)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_247),
.Y(n_252)
);

AOI322xp5_ASAP7_75t_L g250 ( 
.A1(n_248),
.A2(n_240),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_10),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_9),
.C(n_10),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_249),
.A2(n_10),
.B(n_11),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_251),
.C(n_246),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_254),
.C(n_11),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_245),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_12),
.B1(n_13),
.B2(n_248),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_12),
.Y(n_257)
);


endmodule