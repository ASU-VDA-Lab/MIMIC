module fake_jpeg_31735_n_249 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_38),
.Y(n_42)
);

CKINVDCx6p67_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_17),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_53),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_17),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_16),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_59),
.Y(n_67)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_18),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_62),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_18),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_25),
.B(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_35),
.Y(n_85)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_38),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_39),
.B1(n_30),
.B2(n_36),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_68),
.B1(n_76),
.B2(n_79),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_54),
.A2(n_39),
.B1(n_61),
.B2(n_40),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_32),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_78),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_31),
.B1(n_21),
.B2(n_33),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_32),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_50),
.A2(n_40),
.B1(n_36),
.B2(n_31),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_55),
.A2(n_33),
.B1(n_31),
.B2(n_21),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_80),
.A2(n_69),
.B1(n_81),
.B2(n_77),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_21),
.B1(n_29),
.B2(n_26),
.Y(n_84)
);

OAI32xp33_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_96),
.A3(n_76),
.B1(n_80),
.B2(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_90),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_29),
.B1(n_26),
.B2(n_23),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_34),
.B1(n_4),
.B2(n_6),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_46),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_42),
.B(n_23),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_44),
.A2(n_34),
.B1(n_38),
.B2(n_5),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_34),
.B1(n_4),
.B2(n_5),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_42),
.B(n_15),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_2),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_34),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_108),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_47),
.B(n_43),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_109),
.B1(n_112),
.B2(n_127),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_71),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_104),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_114),
.Y(n_134)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_105),
.Y(n_152)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_34),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_110),
.A2(n_111),
.B1(n_118),
.B2(n_120),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_7),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_121),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_96),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_66),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_12),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_67),
.B(n_12),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_72),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_125),
.C(n_103),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_68),
.A2(n_75),
.B(n_65),
.C(n_96),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_81),
.B(n_95),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_69),
.B1(n_93),
.B2(n_95),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_130),
.A2(n_147),
.B1(n_150),
.B2(n_131),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_74),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_116),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_113),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_137),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_74),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_141),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_98),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_121),
.C(n_108),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_126),
.C(n_115),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_144),
.A2(n_151),
.B(n_146),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_100),
.A2(n_127),
.B1(n_103),
.B2(n_124),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_110),
.A2(n_97),
.B1(n_111),
.B2(n_104),
.Y(n_150)
);

NOR2x1_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_154),
.B(n_163),
.Y(n_186)
);

AOI22x1_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_144),
.B1(n_147),
.B2(n_130),
.Y(n_155)
);

OA21x2_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_139),
.B(n_152),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_104),
.C(n_123),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_162),
.C(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_153),
.Y(n_157)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

AOI322xp5_ASAP7_75t_SL g161 ( 
.A1(n_148),
.A2(n_114),
.A3(n_120),
.B1(n_101),
.B2(n_125),
.C1(n_128),
.C2(n_113),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_161),
.B(n_166),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_106),
.C(n_125),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_165),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_105),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_132),
.C(n_149),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_172),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_129),
.A2(n_132),
.B(n_149),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_140),
.B(n_135),
.Y(n_185)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_173),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_133),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_148),
.C(n_146),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_175),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_137),
.Y(n_176)
);

XOR2x2_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_156),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_177),
.A2(n_192),
.B1(n_180),
.B2(n_178),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_164),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_178),
.B(n_180),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_165),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_160),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_182),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_177),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_152),
.B1(n_140),
.B2(n_135),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_188),
.A2(n_157),
.B1(n_159),
.B2(n_162),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_183),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_173),
.A2(n_167),
.B1(n_155),
.B2(n_170),
.Y(n_192)
);

OAI32xp33_ASAP7_75t_L g193 ( 
.A1(n_155),
.A2(n_169),
.A3(n_175),
.B1(n_154),
.B2(n_158),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_171),
.Y(n_194)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_194),
.Y(n_200)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_187),
.B(n_167),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_199),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_207),
.B1(n_177),
.B2(n_194),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_174),
.C(n_176),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_195),
.C(n_183),
.Y(n_211)
);

OAI321xp33_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_168),
.A3(n_189),
.B1(n_181),
.B2(n_192),
.C(n_186),
.Y(n_204)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_205),
.A2(n_208),
.B(n_184),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_206),
.A2(n_210),
.B(n_189),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_185),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_212),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_216),
.A2(n_207),
.B(n_196),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_181),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_217),
.B(n_219),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_220),
.A2(n_210),
.B1(n_202),
.B2(n_197),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_182),
.B(n_206),
.C(n_201),
.Y(n_221)
);

AOI31xp67_ASAP7_75t_L g230 ( 
.A1(n_221),
.A2(n_200),
.A3(n_220),
.B(n_216),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_219),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_198),
.Y(n_225)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_225),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_205),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_227),
.Y(n_235)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_221),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_230),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_225),
.B(n_215),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_224),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_230),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_223),
.A2(n_217),
.B(n_211),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_236),
.B(n_237),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_212),
.C(n_200),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_239),
.B(n_241),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_242),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_231),
.B(n_222),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_226),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_237),
.C(n_233),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_245),
.A2(n_235),
.B(n_234),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_244),
.C(n_228),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_247),
.Y(n_249)
);


endmodule