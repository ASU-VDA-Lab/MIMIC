module fake_jpeg_28450_n_403 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_403);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_403;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_41),
.B(n_48),
.Y(n_86)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_44),
.Y(n_100)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_14),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_51),
.B(n_58),
.Y(n_106)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_23),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_16),
.B(n_14),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_60),
.B(n_70),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_34),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_64),
.B(n_23),
.Y(n_122)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_16),
.B(n_13),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_31),
.B1(n_32),
.B2(n_29),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_72),
.A2(n_80),
.B1(n_84),
.B2(n_94),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_73),
.B(n_89),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_34),
.B(n_38),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_L g162 ( 
.A1(n_77),
.A2(n_49),
.B(n_1),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_39),
.B1(n_33),
.B2(n_32),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_52),
.A2(n_31),
.B1(n_35),
.B2(n_19),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_31),
.B1(n_35),
.B2(n_19),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_65),
.B(n_22),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_87),
.B(n_102),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_22),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_40),
.A2(n_30),
.B1(n_26),
.B2(n_38),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_50),
.A2(n_26),
.B1(n_30),
.B2(n_39),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_110),
.Y(n_137)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_41),
.B(n_13),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

INVx5_ASAP7_75t_SL g109 ( 
.A(n_44),
.Y(n_109)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_57),
.A2(n_39),
.B1(n_27),
.B2(n_21),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_54),
.Y(n_111)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_42),
.Y(n_112)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_112),
.Y(n_172)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_122),
.Y(n_128)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_67),
.A2(n_29),
.B1(n_27),
.B2(n_21),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_119),
.A2(n_69),
.B1(n_20),
.B2(n_29),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_57),
.A2(n_27),
.B1(n_21),
.B2(n_28),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_61),
.Y(n_146)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_124),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_59),
.B1(n_47),
.B2(n_63),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_125),
.A2(n_148),
.B1(n_157),
.B2(n_117),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_64),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_132),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_58),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_134),
.Y(n_216)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_138),
.Y(n_196)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx4_ASAP7_75t_SL g207 ( 
.A(n_139),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_90),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_145),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_79),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_142),
.B(n_147),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_51),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_91),
.C(n_108),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_29),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_146),
.B(n_162),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_71),
.B(n_0),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_100),
.A2(n_69),
.B1(n_20),
.B2(n_28),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_37),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_156),
.Y(n_187)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_74),
.Y(n_153)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_155),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_75),
.B(n_37),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_121),
.A2(n_20),
.B1(n_37),
.B2(n_28),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_119),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_159),
.B(n_160),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_72),
.Y(n_160)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_76),
.B(n_105),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_169),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_93),
.B(n_0),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_140),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_118),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_74),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_85),
.B(n_1),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_173),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_95),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_123),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_10),
.Y(n_210)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_81),
.Y(n_176)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_159),
.A2(n_108),
.B(n_91),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_177),
.A2(n_180),
.B(n_186),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_183),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_179),
.B(n_192),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_88),
.B(n_81),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_85),
.C(n_88),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_184),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_136),
.A2(n_80),
.B1(n_104),
.B2(n_99),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_186),
.A2(n_191),
.B1(n_203),
.B2(n_129),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_117),
.B1(n_104),
.B2(n_3),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_188),
.A2(n_205),
.B1(n_208),
.B2(n_220),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_12),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_149),
.B(n_2),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_197),
.B(n_133),
.Y(n_245)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_135),
.Y(n_198)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_128),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_164),
.B(n_142),
.C(n_166),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_137),
.B(n_4),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_221),
.Y(n_233)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_131),
.Y(n_202)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_146),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_137),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_144),
.A2(n_11),
.B1(n_8),
.B2(n_9),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_210),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_164),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_211),
.B(n_212),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_134),
.B(n_6),
.Y(n_212)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_144),
.A2(n_10),
.B1(n_6),
.B2(n_8),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_175),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_151),
.Y(n_222)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_134),
.B(n_154),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_139),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_154),
.B1(n_175),
.B2(n_172),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_224),
.A2(n_248),
.B1(n_232),
.B2(n_257),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_226),
.A2(n_230),
.B(n_206),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_227),
.B(n_238),
.Y(n_292)
);

NAND3xp33_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_182),
.C(n_190),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_240),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_179),
.B(n_168),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_239),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_152),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_192),
.B(n_168),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_152),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_177),
.A2(n_155),
.B(n_138),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_196),
.B(n_195),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_164),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_249),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_180),
.A2(n_127),
.B1(n_161),
.B2(n_133),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_245),
.B(n_250),
.Y(n_284)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_247),
.Y(n_293)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_181),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_248),
.B(n_257),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_127),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_187),
.B(n_163),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_176),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_251),
.B(n_256),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_259),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_254),
.A2(n_255),
.B1(n_258),
.B2(n_193),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_214),
.A2(n_126),
.B1(n_129),
.B2(n_153),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_178),
.B(n_201),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_181),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_188),
.A2(n_191),
.B1(n_203),
.B2(n_198),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_216),
.B(n_170),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_200),
.B(n_126),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_213),
.C(n_209),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_208),
.A2(n_166),
.B1(n_220),
.B2(n_211),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_263),
.B1(n_207),
.B2(n_218),
.Y(n_280)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_262),
.B(n_264),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_202),
.A2(n_219),
.B1(n_222),
.B2(n_189),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_216),
.B(n_196),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_215),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_265),
.B(n_272),
.C(n_289),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_267),
.A2(n_271),
.B(n_288),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_236),
.A2(n_209),
.B1(n_195),
.B2(n_206),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_269),
.A2(n_278),
.B(n_270),
.Y(n_323)
);

OA21x2_ASAP7_75t_L g270 ( 
.A1(n_226),
.A2(n_194),
.B(n_207),
.Y(n_270)
);

OA21x2_ASAP7_75t_L g310 ( 
.A1(n_270),
.A2(n_267),
.B(n_277),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_245),
.B(n_264),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_194),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_273),
.A2(n_277),
.B(n_246),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_279),
.Y(n_301)
);

AOI221xp5_ASAP7_75t_L g276 ( 
.A1(n_233),
.A2(n_218),
.B1(n_207),
.B2(n_213),
.C(n_193),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g309 ( 
.A(n_276),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_241),
.A2(n_230),
.B(n_242),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_236),
.A2(n_251),
.B1(n_225),
.B2(n_252),
.Y(n_278)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_251),
.C(n_229),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_286),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_229),
.B(n_193),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_287),
.B(n_296),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_255),
.A2(n_256),
.B(n_260),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_237),
.B(n_193),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_258),
.A2(n_254),
.B1(n_247),
.B2(n_233),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_291),
.A2(n_298),
.B1(n_232),
.B2(n_246),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_280),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_234),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_295),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_239),
.B(n_235),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_235),
.B(n_244),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_297),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_225),
.A2(n_253),
.B1(n_263),
.B2(n_244),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_302),
.A2(n_303),
.B1(n_306),
.B2(n_316),
.Y(n_331)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_297),
.Y(n_304)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_304),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_298),
.A2(n_252),
.B1(n_262),
.B2(n_278),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_282),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_307),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_275),
.A2(n_295),
.B1(n_269),
.B2(n_270),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_308),
.A2(n_315),
.B1(n_317),
.B2(n_319),
.Y(n_338)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_282),
.Y(n_313)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_313),
.Y(n_333)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_314),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_266),
.B(n_284),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_293),
.A2(n_291),
.B1(n_275),
.B2(n_281),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_283),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_283),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_318),
.Y(n_339)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_293),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_320),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_287),
.B(n_285),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_292),
.B(n_288),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_265),
.B(n_272),
.C(n_290),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_326),
.C(n_274),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_279),
.B(n_290),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_279),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_327),
.B(n_330),
.C(n_332),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_312),
.A2(n_281),
.B1(n_270),
.B2(n_273),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_328),
.A2(n_336),
.B1(n_348),
.B2(n_315),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_290),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_289),
.C(n_268),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_334),
.B(n_335),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_268),
.C(n_292),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_312),
.A2(n_286),
.B1(n_323),
.B2(n_300),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_303),
.A2(n_316),
.B1(n_306),
.B2(n_302),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_337),
.A2(n_317),
.B1(n_310),
.B2(n_299),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_301),
.B(n_326),
.C(n_300),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_342),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_305),
.Y(n_342)
);

BUFx12f_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_343),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_304),
.B(n_313),
.C(n_305),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_342),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_314),
.A2(n_307),
.B1(n_318),
.B2(n_321),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_349),
.A2(n_350),
.B1(n_343),
.B2(n_330),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_331),
.A2(n_299),
.B1(n_310),
.B2(n_319),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_352),
.A2(n_365),
.B1(n_358),
.B2(n_356),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_335),
.B(n_309),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_357),
.Y(n_373)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_333),
.Y(n_356)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_356),
.Y(n_370)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_348),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_329),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_359),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_338),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_346),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_362),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_339),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_360),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_344),
.A2(n_337),
.B1(n_331),
.B2(n_339),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_364),
.A2(n_366),
.B1(n_343),
.B2(n_359),
.Y(n_371)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_347),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_340),
.A2(n_345),
.B1(n_336),
.B2(n_328),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_332),
.C(n_341),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_367),
.B(n_369),
.C(n_376),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_368),
.A2(n_371),
.B1(n_373),
.B2(n_380),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_334),
.C(n_327),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_355),
.A2(n_357),
.B(n_351),
.Y(n_372)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_372),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_374),
.B(n_375),
.Y(n_381)
);

BUFx24_ASAP7_75t_SL g375 ( 
.A(n_365),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_354),
.B(n_352),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_362),
.C(n_350),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_379),
.B(n_380),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_360),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_385),
.B(n_386),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_379),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_378),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_387),
.B(n_388),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_383),
.A2(n_367),
.B(n_369),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_389),
.A2(n_393),
.B(n_386),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_368),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_392),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_385),
.A2(n_376),
.B(n_370),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_394),
.B(n_395),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_390),
.B(n_391),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_396),
.A2(n_393),
.B(n_382),
.Y(n_397)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_397),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_398),
.B(n_381),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_399),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_401),
.B(n_400),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_402),
.B(n_382),
.Y(n_403)
);


endmodule