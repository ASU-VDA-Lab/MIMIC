module fake_jpeg_101_n_97 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_97);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_97;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_24),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_32),
.C(n_2),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_1),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_29),
.B(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_47),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_32),
.B1(n_28),
.B2(n_33),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_36),
.B1(n_38),
.B2(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_1),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_56),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_50),
.B(n_2),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_64),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_43),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_13),
.C(n_22),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_12),
.C(n_20),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_3),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_74),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_79),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_75),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_69),
.B(n_3),
.Y(n_81)
);

AOI221xp5_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.C(n_9),
.Y(n_85)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_83),
.Y(n_87)
);

NOR3xp33_ASAP7_75t_SL g89 ( 
.A(n_85),
.B(n_76),
.C(n_81),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_82),
.A2(n_4),
.B(n_10),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_11),
.C(n_15),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_90),
.B(n_88),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_87),
.Y(n_93)
);

OAI221xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_84),
.B1(n_77),
.B2(n_18),
.C(n_23),
.Y(n_94)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_94),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_16),
.Y(n_97)
);


endmodule