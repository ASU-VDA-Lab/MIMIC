module fake_jpeg_16280_n_391 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_391);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_391;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_38),
.B(n_40),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_52),
.Y(n_96)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_28),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_28),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_53),
.B(n_54),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_27),
.B(n_13),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_65),
.Y(n_98)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_1),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_19),
.B1(n_21),
.B2(n_27),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_81),
.B(n_15),
.Y(n_164)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_17),
.C(n_33),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_36),
.Y(n_120)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_89),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_46),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_48),
.A2(n_25),
.B1(n_36),
.B2(n_31),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_32),
.B1(n_31),
.B2(n_25),
.Y(n_125)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_93),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_103),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_55),
.A2(n_34),
.B1(n_29),
.B2(n_35),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_32),
.B1(n_31),
.B2(n_37),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_108),
.Y(n_130)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_40),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_17),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_21),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_110),
.B(n_115),
.Y(n_135)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_21),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_38),
.B(n_19),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_116),
.B(n_29),
.Y(n_152)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_45),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_36),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_119),
.B(n_149),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_120),
.A2(n_125),
.B1(n_147),
.B2(n_80),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_74),
.A2(n_19),
.B1(n_34),
.B2(n_35),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_121),
.A2(n_109),
.B1(n_80),
.B2(n_13),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_86),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_138),
.Y(n_172)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_132),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_133),
.A2(n_101),
.B1(n_70),
.B2(n_105),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_91),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_160),
.B1(n_161),
.B2(n_119),
.Y(n_170)
);

OR2x2_ASAP7_75t_SL g137 ( 
.A(n_98),
.B(n_37),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_SL g210 ( 
.A1(n_137),
.A2(n_164),
.B(n_5),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_92),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_68),
.B(n_71),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_139),
.B(n_2),
.C(n_4),
.Y(n_200)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_77),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_144),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_67),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_94),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_151),
.Y(n_185)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_146),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_75),
.A2(n_29),
.B1(n_22),
.B2(n_15),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_148),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_33),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_96),
.B(n_33),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_166),
.Y(n_190)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_152),
.B(n_154),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_103),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_159),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_111),
.B(n_22),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_77),
.B(n_102),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_76),
.A2(n_82),
.B1(n_100),
.B2(n_105),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_101),
.A2(n_22),
.B1(n_15),
.B2(n_16),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_73),
.B(n_33),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_74),
.B(n_2),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_150),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_83),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_12),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_170),
.A2(n_177),
.B1(n_189),
.B2(n_187),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_162),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_171),
.B(n_173),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_SL g217 ( 
.A1(n_174),
.A2(n_186),
.B(n_177),
.C(n_189),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_179),
.B(n_181),
.Y(n_238)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_149),
.B(n_33),
.CI(n_17),
.CON(n_181),
.SN(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_183),
.Y(n_240)
);

OAI32xp33_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_16),
.A3(n_33),
.B1(n_94),
.B2(n_11),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_186),
.B(n_192),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_188),
.B(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_191),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_120),
.B(n_16),
.C(n_10),
.Y(n_192)
);

AOI32xp33_ASAP7_75t_L g193 ( 
.A1(n_120),
.A2(n_90),
.A3(n_83),
.B1(n_12),
.B2(n_11),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_200),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_90),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_133),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_195),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_118),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_197),
.Y(n_222)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_207),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_166),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_201),
.A2(n_205),
.B1(n_130),
.B2(n_128),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_4),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_203),
.A2(n_211),
.B(n_7),
.Y(n_249)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_122),
.Y(n_204)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

AO22x1_ASAP7_75t_SL g205 ( 
.A1(n_136),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_126),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_158),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_213),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_200),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_167),
.B(n_160),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_141),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_131),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_214),
.B(n_185),
.Y(n_253)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_8),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_216),
.B(n_252),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_217),
.A2(n_176),
.B1(n_204),
.B2(n_215),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_190),
.B(n_139),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_218),
.A2(n_221),
.B(n_248),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_219),
.A2(n_209),
.B1(n_199),
.B2(n_202),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_170),
.A2(n_156),
.B1(n_141),
.B2(n_128),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_220),
.A2(n_232),
.B1(n_245),
.B2(n_254),
.Y(n_268)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_139),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_229),
.Y(n_263)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_246),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_135),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_123),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_199),
.Y(n_274)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_182),
.A2(n_156),
.B1(n_155),
.B2(n_151),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_233),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_155),
.B1(n_123),
.B2(n_145),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_242),
.B1(n_244),
.B2(n_247),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_176),
.A2(n_129),
.B1(n_146),
.B2(n_142),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_211),
.A2(n_137),
.B1(n_122),
.B2(n_131),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_205),
.A2(n_132),
.B1(n_148),
.B2(n_7),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_179),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_SL g248 ( 
.A1(n_205),
.A2(n_7),
.B(n_8),
.C(n_165),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_249),
.A2(n_203),
.B(n_201),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_251),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_172),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_179),
.A2(n_181),
.B1(n_192),
.B2(n_203),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_184),
.B(n_206),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_255),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_256),
.A2(n_249),
.B(n_221),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_281),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_239),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_261),
.B(n_264),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_240),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_175),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_273),
.C(n_237),
.Y(n_297)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_225),
.Y(n_266)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_266),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_267),
.A2(n_288),
.B1(n_258),
.B2(n_276),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_221),
.A2(n_169),
.B(n_206),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_248),
.B(n_247),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_272),
.A2(n_277),
.B1(n_283),
.B2(n_286),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_229),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_284),
.Y(n_292)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_241),
.Y(n_275)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_275),
.Y(n_309)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_231),
.Y(n_276)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_276),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_223),
.A2(n_202),
.B1(n_217),
.B2(n_218),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_278),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_227),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_279),
.B(n_282),
.Y(n_303)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_228),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_217),
.A2(n_218),
.B1(n_221),
.B2(n_220),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_230),
.B(n_216),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_250),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_285),
.B(n_288),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_217),
.A2(n_236),
.B1(n_237),
.B2(n_244),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_224),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_234),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_293),
.A2(n_257),
.B(n_289),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_294),
.A2(n_296),
.B(n_308),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_263),
.B(n_232),
.Y(n_295)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_295),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_235),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_297),
.B(n_290),
.Y(n_334)
);

XOR2x2_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_256),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_298),
.A2(n_280),
.B(n_258),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_224),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_299),
.B(n_317),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_235),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_313),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_222),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_311),
.C(n_312),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_248),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_265),
.B(n_243),
.C(n_245),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_226),
.C(n_246),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_274),
.B(n_248),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_272),
.A2(n_286),
.B1(n_287),
.B2(n_284),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_314),
.A2(n_315),
.B1(n_316),
.B2(n_280),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_270),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_289),
.B(n_262),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_257),
.B(n_266),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_318),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_319),
.A2(n_301),
.B(n_307),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_298),
.A2(n_268),
.B1(n_259),
.B2(n_282),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_320),
.A2(n_323),
.B1(n_332),
.B2(n_338),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_321),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_322),
.A2(n_330),
.B1(n_328),
.B2(n_325),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_308),
.A2(n_268),
.B1(n_259),
.B2(n_271),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_260),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_331),
.C(n_334),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_327),
.A2(n_329),
.B(n_335),
.Y(n_356)
);

MAJx2_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_291),
.C(n_306),
.Y(n_329)
);

AO22x1_ASAP7_75t_L g330 ( 
.A1(n_313),
.A2(n_293),
.B1(n_294),
.B2(n_292),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_319),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_312),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_308),
.A2(n_278),
.B1(n_290),
.B2(n_305),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_296),
.A2(n_295),
.B(n_292),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_296),
.A2(n_318),
.B1(n_315),
.B2(n_302),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_303),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_339),
.B(n_309),
.C(n_304),
.Y(n_342)
);

AO21x1_ASAP7_75t_L g340 ( 
.A1(n_302),
.A2(n_309),
.B(n_310),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_340),
.B(n_307),
.Y(n_346)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_337),
.Y(n_341)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_341),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_342),
.B(n_350),
.C(n_345),
.Y(n_366)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_343),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_346),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_347),
.A2(n_354),
.B1(n_355),
.B2(n_353),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_336),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_352),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_334),
.C(n_324),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_332),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_351),
.B(n_353),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_340),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_335),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_338),
.A2(n_323),
.B1(n_325),
.B2(n_320),
.Y(n_355)
);

OAI21x1_ASAP7_75t_L g357 ( 
.A1(n_326),
.A2(n_339),
.B(n_329),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_357),
.Y(n_365)
);

AOI21x1_ASAP7_75t_L g358 ( 
.A1(n_346),
.A2(n_324),
.B(n_347),
.Y(n_358)
);

O2A1O1Ixp33_ASAP7_75t_L g371 ( 
.A1(n_358),
.A2(n_357),
.B(n_342),
.C(n_356),
.Y(n_371)
);

AO221x1_ASAP7_75t_L g361 ( 
.A1(n_344),
.A2(n_343),
.B1(n_352),
.B2(n_354),
.C(n_351),
.Y(n_361)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_361),
.Y(n_376)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_363),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_366),
.B(n_356),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_342),
.B(n_350),
.C(n_345),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_367),
.B(n_350),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_355),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_368),
.B(n_349),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_370),
.B(n_373),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_371),
.B(n_374),
.Y(n_379)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_359),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_375),
.B(n_366),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_375),
.B(n_367),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_365),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_380),
.A2(n_365),
.B1(n_358),
.B2(n_362),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_379),
.B(n_376),
.C(n_370),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_381),
.B(n_382),
.Y(n_385)
);

NOR3xp33_ASAP7_75t_L g384 ( 
.A(n_383),
.B(n_369),
.C(n_377),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_384),
.B(n_381),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_386),
.A2(n_385),
.B(n_377),
.Y(n_387)
);

OAI221xp5_ASAP7_75t_L g388 ( 
.A1(n_387),
.A2(n_369),
.B1(n_372),
.B2(n_344),
.C(n_364),
.Y(n_388)
);

O2A1O1Ixp33_ASAP7_75t_SL g389 ( 
.A1(n_388),
.A2(n_360),
.B(n_341),
.C(n_372),
.Y(n_389)
);

FAx1_ASAP7_75t_SL g390 ( 
.A(n_389),
.B(n_363),
.CI(n_349),
.CON(n_390),
.SN(n_390)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_390),
.B(n_368),
.Y(n_391)
);


endmodule