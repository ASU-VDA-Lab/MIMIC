module fake_jpeg_28324_n_146 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_146);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_19),
.B(n_5),
.Y(n_20)
);

OAI21xp33_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_21),
.B(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_0),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_0),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_11),
.C(n_16),
.Y(n_33)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_34),
.B1(n_35),
.B2(n_24),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_23),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_24),
.A2(n_17),
.B1(n_18),
.B2(n_13),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_24),
.A2(n_17),
.B1(n_18),
.B2(n_13),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_23),
.B1(n_27),
.B2(n_26),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_35),
.B1(n_34),
.B2(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_23),
.B1(n_27),
.B2(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_47),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_25),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_25),
.Y(n_47)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_23),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_63),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_64),
.B1(n_56),
.B2(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_50),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_41),
.B1(n_47),
.B2(n_27),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_65),
.B(n_69),
.Y(n_72)
);

AOI32xp33_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_41),
.A3(n_20),
.B1(n_22),
.B2(n_30),
.Y(n_67)
);

AOI221xp5_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_54),
.B1(n_53),
.B2(n_48),
.C(n_50),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_41),
.B(n_20),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_49),
.B(n_14),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_70),
.B(n_13),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_76),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_74),
.B(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_70),
.B(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_81),
.B1(n_26),
.B2(n_36),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_80),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_60),
.B1(n_66),
.B2(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_48),
.B1(n_55),
.B2(n_36),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_52),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_26),
.B1(n_29),
.B2(n_52),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_66),
.C(n_58),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_22),
.C(n_11),
.Y(n_107)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_90),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_89),
.A2(n_91),
.B(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_14),
.C(n_10),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_46),
.B1(n_45),
.B2(n_58),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_18),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_97),
.A2(n_102),
.B(n_16),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_30),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_100),
.B1(n_106),
.B2(n_107),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_11),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_30),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_86),
.B(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_45),
.B1(n_16),
.B2(n_29),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_SL g109 ( 
.A1(n_101),
.A2(n_89),
.B(n_93),
.C(n_88),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_112),
.B1(n_98),
.B2(n_108),
.Y(n_119)
);

OAI21x1_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_94),
.B(n_96),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_111),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_93),
.B1(n_29),
.B2(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_116),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_30),
.A3(n_15),
.B1(n_14),
.B2(n_10),
.C1(n_12),
.C2(n_22),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_117),
.B(n_107),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_121),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_97),
.C(n_105),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_29),
.B1(n_16),
.B2(n_15),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_22),
.C(n_15),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_109),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_109),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_120),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_0),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_112),
.B(n_10),
.C(n_12),
.Y(n_128)
);

OAI321xp33_ASAP7_75t_L g135 ( 
.A1(n_128),
.A2(n_5),
.A3(n_8),
.B1(n_7),
.B2(n_4),
.C(n_9),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_133),
.B(n_134),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_130),
.A2(n_124),
.B1(n_12),
.B2(n_6),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_4),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_4),
.B(n_6),
.Y(n_139)
);

AOI322xp5_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_138),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_137),
.C2(n_132),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_R g138 ( 
.A1(n_133),
.A2(n_129),
.B(n_130),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_139),
.A2(n_1),
.B(n_2),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_1),
.B(n_2),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_SL g145 ( 
.A1(n_144),
.A2(n_143),
.B(n_1),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_3),
.Y(n_146)
);


endmodule