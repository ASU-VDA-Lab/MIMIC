module real_aes_8430_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g187 ( .A1(n_0), .A2(n_188), .B(n_189), .C(n_193), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_1), .B(n_183), .Y(n_194) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_2), .B(n_90), .C(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g444 ( .A(n_2), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_3), .B(n_148), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_4), .A2(n_129), .B(n_479), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_5), .A2(n_134), .B(n_139), .C(n_515), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_6), .A2(n_129), .B(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_7), .B(n_183), .Y(n_485) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_8), .A2(n_162), .B(n_212), .Y(n_211) );
AND2x6_ASAP7_75t_L g134 ( .A(n_9), .B(n_135), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_10), .A2(n_134), .B(n_139), .C(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g540 ( .A(n_11), .Y(n_540) );
INVx1_ASAP7_75t_L g106 ( .A(n_12), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_12), .B(n_39), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_13), .B(n_192), .Y(n_517) );
INVx1_ASAP7_75t_L g158 ( .A(n_14), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_15), .B(n_148), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_16), .A2(n_149), .B(n_525), .C(n_527), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_17), .B(n_183), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_18), .B(n_176), .Y(n_569) );
A2O1A1Ixp33_ASAP7_75t_L g169 ( .A1(n_19), .A2(n_139), .B(n_170), .C(n_175), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_20), .A2(n_191), .B(n_206), .C(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_21), .B(n_192), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_22), .A2(n_76), .B1(n_734), .B2(n_735), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_22), .Y(n_735) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_23), .B(n_192), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g466 ( .A(n_24), .Y(n_466) );
INVx1_ASAP7_75t_L g491 ( .A(n_25), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_26), .A2(n_139), .B(n_175), .C(n_215), .Y(n_214) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_27), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_28), .Y(n_513) );
INVx1_ASAP7_75t_L g567 ( .A(n_29), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_30), .A2(n_129), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g132 ( .A(n_31), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g136 ( .A1(n_32), .A2(n_137), .B(n_142), .C(n_152), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_33), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_34), .A2(n_191), .B(n_482), .C(n_484), .Y(n_481) );
INVxp67_ASAP7_75t_L g568 ( .A(n_35), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_36), .B(n_217), .Y(n_216) );
CKINVDCx14_ASAP7_75t_R g480 ( .A(n_37), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_38), .A2(n_139), .B(n_175), .C(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_39), .B(n_106), .Y(n_105) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_40), .A2(n_193), .B(n_538), .C(n_539), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_41), .B(n_168), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_42), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_43), .B(n_148), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_44), .B(n_129), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_45), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_46), .Y(n_564) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_47), .A2(n_137), .B(n_152), .C(n_226), .Y(n_225) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_48), .A2(n_87), .B1(n_119), .B2(n_120), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_48), .Y(n_120) );
INVx1_ASAP7_75t_L g190 ( .A(n_49), .Y(n_190) );
INVx1_ASAP7_75t_L g227 ( .A(n_50), .Y(n_227) );
INVx1_ASAP7_75t_L g503 ( .A(n_51), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_52), .B(n_129), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_53), .Y(n_179) );
CKINVDCx14_ASAP7_75t_R g536 ( .A(n_54), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_55), .Y(n_447) );
INVx1_ASAP7_75t_L g135 ( .A(n_56), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_57), .B(n_129), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_58), .B(n_183), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_59), .A2(n_174), .B(n_237), .C(n_239), .Y(n_236) );
INVx1_ASAP7_75t_L g157 ( .A(n_60), .Y(n_157) );
INVx1_ASAP7_75t_SL g483 ( .A(n_61), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_62), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_63), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_64), .B(n_183), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_65), .B(n_149), .Y(n_203) );
INVx1_ASAP7_75t_L g469 ( .A(n_66), .Y(n_469) );
CKINVDCx16_ASAP7_75t_R g186 ( .A(n_67), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_68), .B(n_145), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_69), .A2(n_139), .B(n_152), .C(n_263), .Y(n_262) );
CKINVDCx16_ASAP7_75t_R g235 ( .A(n_70), .Y(n_235) );
INVx1_ASAP7_75t_L g110 ( .A(n_71), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_72), .A2(n_129), .B(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_73), .A2(n_102), .B1(n_111), .B2(n_746), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_74), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_75), .A2(n_129), .B(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_76), .Y(n_734) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_77), .A2(n_168), .B(n_563), .Y(n_562) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_78), .Y(n_488) );
INVx1_ASAP7_75t_L g523 ( .A(n_79), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_80), .B(n_144), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_81), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_82), .A2(n_129), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g526 ( .A(n_83), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_84), .Y(n_745) );
INVx2_ASAP7_75t_L g155 ( .A(n_85), .Y(n_155) );
INVx1_ASAP7_75t_L g516 ( .A(n_86), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_87), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_88), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_89), .B(n_192), .Y(n_204) );
OR2x2_ASAP7_75t_L g441 ( .A(n_90), .B(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g452 ( .A(n_90), .B(n_443), .Y(n_452) );
INVx2_ASAP7_75t_L g456 ( .A(n_90), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_91), .A2(n_139), .B(n_152), .C(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_92), .B(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g143 ( .A(n_93), .Y(n_143) );
INVxp67_ASAP7_75t_L g240 ( .A(n_94), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_95), .B(n_162), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_96), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g199 ( .A(n_97), .Y(n_199) );
INVx1_ASAP7_75t_L g264 ( .A(n_98), .Y(n_264) );
INVx2_ASAP7_75t_L g506 ( .A(n_99), .Y(n_506) );
AND2x2_ASAP7_75t_L g229 ( .A(n_100), .B(n_154), .Y(n_229) );
CKINVDCx6p67_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_103), .Y(n_747) );
CKINVDCx9p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
OAI21x1_ASAP7_75t_SL g111 ( .A1(n_112), .A2(n_116), .B(n_448), .Y(n_111) );
OAI21xp5_ASAP7_75t_SL g448 ( .A1(n_112), .A2(n_446), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_439), .B(n_446), .Y(n_116) );
XOR2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_121), .Y(n_117) );
INVx2_ASAP7_75t_L g453 ( .A(n_121), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_121), .A2(n_737), .B1(n_740), .B2(n_741), .Y(n_736) );
OR3x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_353), .C(n_396), .Y(n_121) );
NAND5xp2_ASAP7_75t_L g122 ( .A(n_123), .B(n_280), .C(n_310), .D(n_327), .E(n_342), .Y(n_122) );
AOI221xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_195), .B1(n_242), .B2(n_248), .C(n_252), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_164), .Y(n_124) );
OR2x2_ASAP7_75t_L g257 ( .A(n_125), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g297 ( .A(n_125), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g315 ( .A(n_125), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_125), .B(n_250), .Y(n_332) );
OR2x2_ASAP7_75t_L g344 ( .A(n_125), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_125), .B(n_303), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_125), .B(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_125), .B(n_281), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_125), .B(n_289), .Y(n_395) );
AND2x2_ASAP7_75t_L g427 ( .A(n_125), .B(n_181), .Y(n_427) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_125), .Y(n_435) );
INVx5_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_126), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g254 ( .A(n_126), .B(n_230), .Y(n_254) );
BUFx2_ASAP7_75t_L g277 ( .A(n_126), .Y(n_277) );
AND2x2_ASAP7_75t_L g306 ( .A(n_126), .B(n_165), .Y(n_306) );
AND2x2_ASAP7_75t_L g361 ( .A(n_126), .B(n_258), .Y(n_361) );
OR2x6_ASAP7_75t_L g126 ( .A(n_127), .B(n_159), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_136), .B(n_154), .Y(n_127) );
BUFx2_ASAP7_75t_L g168 ( .A(n_129), .Y(n_168) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_134), .Y(n_129) );
NAND2x1p5_ASAP7_75t_L g200 ( .A(n_130), .B(n_134), .Y(n_200) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
INVx1_ASAP7_75t_L g174 ( .A(n_131), .Y(n_174) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
INVx1_ASAP7_75t_L g207 ( .A(n_132), .Y(n_207) );
INVx1_ASAP7_75t_L g141 ( .A(n_133), .Y(n_141) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_133), .Y(n_146) );
INVx3_ASAP7_75t_L g149 ( .A(n_133), .Y(n_149) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_133), .Y(n_192) );
INVx1_ASAP7_75t_L g217 ( .A(n_133), .Y(n_217) );
INVx4_ASAP7_75t_SL g153 ( .A(n_134), .Y(n_153) );
BUFx3_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
O2A1O1Ixp33_ASAP7_75t_SL g185 ( .A1(n_138), .A2(n_153), .B(n_186), .C(n_187), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g234 ( .A1(n_138), .A2(n_153), .B(n_235), .C(n_236), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_138), .A2(n_153), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g502 ( .A1(n_138), .A2(n_153), .B(n_503), .C(n_504), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_SL g522 ( .A1(n_138), .A2(n_153), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_SL g535 ( .A1(n_138), .A2(n_153), .B(n_536), .C(n_537), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_SL g563 ( .A1(n_138), .A2(n_153), .B(n_564), .C(n_565), .Y(n_563) );
INVx5_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
BUFx3_ASAP7_75t_L g151 ( .A(n_140), .Y(n_151) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_140), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_147), .C(n_150), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_144), .A2(n_150), .B(n_227), .C(n_228), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_144), .A2(n_469), .B(n_470), .C(n_471), .Y(n_468) );
O2A1O1Ixp5_ASAP7_75t_L g515 ( .A1(n_144), .A2(n_471), .B(n_516), .C(n_517), .Y(n_515) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx4_ASAP7_75t_L g238 ( .A(n_146), .Y(n_238) );
INVx2_ASAP7_75t_L g188 ( .A(n_148), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_148), .B(n_240), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_148), .A2(n_173), .B(n_491), .C(n_492), .Y(n_490) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_148), .A2(n_238), .B1(n_567), .B2(n_568), .Y(n_566) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_149), .B(n_540), .Y(n_539) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g193 ( .A(n_151), .Y(n_193) );
INVx1_ASAP7_75t_L g527 ( .A(n_151), .Y(n_527) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g177 ( .A(n_154), .Y(n_177) );
INVx1_ASAP7_75t_L g180 ( .A(n_154), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_154), .A2(n_224), .B(n_225), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_154), .A2(n_200), .B(n_488), .C(n_489), .Y(n_487) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_154), .A2(n_534), .B(n_541), .Y(n_533) );
AND2x2_ASAP7_75t_SL g154 ( .A(n_155), .B(n_156), .Y(n_154) );
AND2x2_ASAP7_75t_L g163 ( .A(n_155), .B(n_156), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
INVx3_ASAP7_75t_L g183 ( .A(n_161), .Y(n_183) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_161), .A2(n_198), .B(n_208), .Y(n_197) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_161), .A2(n_261), .B(n_269), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_161), .B(n_270), .Y(n_269) );
AO21x2_ASAP7_75t_L g464 ( .A1(n_161), .A2(n_465), .B(n_472), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_161), .B(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_161), .B(n_519), .Y(n_518) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_162), .A2(n_213), .B(n_214), .Y(n_212) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_162), .Y(n_232) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g210 ( .A(n_163), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_164), .B(n_315), .Y(n_324) );
OAI32xp33_ASAP7_75t_L g338 ( .A1(n_164), .A2(n_274), .A3(n_339), .B1(n_340), .B2(n_341), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_164), .B(n_340), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_164), .B(n_257), .Y(n_381) );
INVx1_ASAP7_75t_SL g410 ( .A(n_164), .Y(n_410) );
NAND4xp25_ASAP7_75t_L g419 ( .A(n_164), .B(n_197), .C(n_361), .D(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g164 ( .A(n_165), .B(n_181), .Y(n_164) );
INVx5_ASAP7_75t_L g251 ( .A(n_165), .Y(n_251) );
AND2x2_ASAP7_75t_L g281 ( .A(n_165), .B(n_182), .Y(n_281) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_165), .Y(n_360) );
AND2x2_ASAP7_75t_L g430 ( .A(n_165), .B(n_377), .Y(n_430) );
OR2x6_ASAP7_75t_L g165 ( .A(n_166), .B(n_178), .Y(n_165) );
AOI21xp5_ASAP7_75t_SL g166 ( .A1(n_167), .A2(n_169), .B(n_176), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_173), .Y(n_170) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_174), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_177), .B(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_180), .A2(n_512), .B(n_518), .Y(n_511) );
AND2x4_ASAP7_75t_L g303 ( .A(n_181), .B(n_251), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_181), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g337 ( .A(n_181), .B(n_258), .Y(n_337) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g250 ( .A(n_182), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g289 ( .A(n_182), .B(n_260), .Y(n_289) );
AND2x2_ASAP7_75t_L g298 ( .A(n_182), .B(n_259), .Y(n_298) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_194), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_191), .B(n_483), .Y(n_482) );
INVx4_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g538 ( .A(n_192), .Y(n_538) );
INVx2_ASAP7_75t_L g471 ( .A(n_193), .Y(n_471) );
AOI222xp33_ASAP7_75t_L g366 ( .A1(n_195), .A2(n_367), .B1(n_369), .B2(n_371), .C1(n_374), .C2(n_375), .Y(n_366) );
AND2x4_ASAP7_75t_L g195 ( .A(n_196), .B(n_219), .Y(n_195) );
AND2x2_ASAP7_75t_L g299 ( .A(n_196), .B(n_300), .Y(n_299) );
NAND3xp33_ASAP7_75t_L g416 ( .A(n_196), .B(n_277), .C(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_211), .Y(n_196) );
INVx5_ASAP7_75t_SL g247 ( .A(n_197), .Y(n_247) );
OAI322xp33_ASAP7_75t_L g252 ( .A1(n_197), .A2(n_253), .A3(n_255), .B1(n_256), .B2(n_271), .C1(n_274), .C2(n_276), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_197), .B(n_245), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_197), .B(n_231), .Y(n_425) );
OAI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_201), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_200), .A2(n_466), .B(n_467), .Y(n_465) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_200), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_205), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_205), .A2(n_216), .B(n_218), .Y(n_215) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
INVx2_ASAP7_75t_L g561 ( .A(n_210), .Y(n_561) );
INVx2_ASAP7_75t_L g245 ( .A(n_211), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_211), .B(n_221), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_219), .B(n_284), .Y(n_339) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
OR2x2_ASAP7_75t_L g318 ( .A(n_220), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_230), .Y(n_220) );
OR2x2_ASAP7_75t_L g246 ( .A(n_221), .B(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_221), .B(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g286 ( .A(n_221), .B(n_231), .Y(n_286) );
AND2x2_ASAP7_75t_L g309 ( .A(n_221), .B(n_245), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_221), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g325 ( .A(n_221), .B(n_284), .Y(n_325) );
AND2x2_ASAP7_75t_L g333 ( .A(n_221), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_221), .B(n_293), .Y(n_383) );
INVx5_ASAP7_75t_SL g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g273 ( .A(n_222), .B(n_247), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_222), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g300 ( .A(n_222), .B(n_231), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_222), .B(n_347), .Y(n_388) );
OR2x2_ASAP7_75t_L g404 ( .A(n_222), .B(n_348), .Y(n_404) );
AND2x2_ASAP7_75t_SL g411 ( .A(n_222), .B(n_365), .Y(n_411) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_222), .Y(n_418) );
OR2x6_ASAP7_75t_L g222 ( .A(n_223), .B(n_229), .Y(n_222) );
AND2x2_ASAP7_75t_L g272 ( .A(n_230), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g322 ( .A(n_230), .B(n_245), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_230), .B(n_247), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_230), .B(n_284), .Y(n_406) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_231), .B(n_247), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_231), .B(n_245), .Y(n_294) );
OR2x2_ASAP7_75t_L g348 ( .A(n_231), .B(n_245), .Y(n_348) );
AND2x2_ASAP7_75t_L g365 ( .A(n_231), .B(n_244), .Y(n_365) );
INVxp67_ASAP7_75t_L g387 ( .A(n_231), .Y(n_387) );
AND2x2_ASAP7_75t_L g414 ( .A(n_231), .B(n_284), .Y(n_414) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_231), .Y(n_421) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_241), .Y(n_231) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_232), .A2(n_478), .B(n_485), .Y(n_477) );
OA21x2_ASAP7_75t_L g500 ( .A1(n_232), .A2(n_501), .B(n_507), .Y(n_500) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_232), .A2(n_521), .B(n_528), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_237), .A2(n_264), .B(n_265), .C(n_266), .Y(n_263) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_238), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_238), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_246), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_244), .B(n_295), .Y(n_368) );
INVx1_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g284 ( .A(n_245), .B(n_247), .Y(n_284) );
OR2x2_ASAP7_75t_L g351 ( .A(n_245), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g295 ( .A(n_246), .Y(n_295) );
OR2x2_ASAP7_75t_L g356 ( .A(n_246), .B(n_348), .Y(n_356) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g255 ( .A(n_250), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_250), .B(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g256 ( .A(n_251), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_251), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_251), .B(n_258), .Y(n_291) );
INVx2_ASAP7_75t_L g336 ( .A(n_251), .Y(n_336) );
AND2x2_ASAP7_75t_L g349 ( .A(n_251), .B(n_289), .Y(n_349) );
AND2x2_ASAP7_75t_L g374 ( .A(n_251), .B(n_298), .Y(n_374) );
INVx1_ASAP7_75t_L g326 ( .A(n_256), .Y(n_326) );
INVx2_ASAP7_75t_SL g313 ( .A(n_257), .Y(n_313) );
INVx1_ASAP7_75t_L g316 ( .A(n_258), .Y(n_316) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_259), .Y(n_279) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx2_ASAP7_75t_L g377 ( .A(n_260), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_268), .Y(n_261) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx3_ASAP7_75t_L g484 ( .A(n_267), .Y(n_484) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g346 ( .A(n_273), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g352 ( .A(n_273), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_273), .A2(n_355), .B1(n_357), .B2(n_362), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_273), .B(n_365), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_274), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g308 ( .A(n_275), .Y(n_308) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
OR2x2_ASAP7_75t_L g290 ( .A(n_277), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_277), .B(n_281), .Y(n_341) );
AND2x2_ASAP7_75t_L g364 ( .A(n_277), .B(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g340 ( .A(n_279), .Y(n_340) );
AOI211xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B(n_287), .C(n_301), .Y(n_280) );
INVx1_ASAP7_75t_L g304 ( .A(n_281), .Y(n_304) );
OAI221xp5_ASAP7_75t_SL g412 ( .A1(n_281), .A2(n_413), .B1(n_415), .B2(n_416), .C(n_419), .Y(n_412) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g431 ( .A(n_284), .Y(n_431) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g380 ( .A(n_286), .B(n_319), .Y(n_380) );
A2O1A1Ixp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_290), .B(n_292), .C(n_296), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
OAI32xp33_ASAP7_75t_L g405 ( .A1(n_294), .A2(n_295), .A3(n_358), .B1(n_395), .B2(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
AND2x2_ASAP7_75t_L g437 ( .A(n_297), .B(n_336), .Y(n_437) );
AND2x2_ASAP7_75t_L g384 ( .A(n_298), .B(n_336), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_298), .B(n_306), .Y(n_402) );
AOI31xp33_ASAP7_75t_SL g301 ( .A1(n_302), .A2(n_304), .A3(n_305), .B(n_307), .Y(n_301) );
INVxp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_303), .B(n_315), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_303), .B(n_313), .Y(n_400) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_303), .A2(n_333), .B1(n_423), .B2(n_426), .C(n_428), .Y(n_422) );
CKINVDCx16_ASAP7_75t_R g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
AND2x2_ASAP7_75t_L g328 ( .A(n_308), .B(n_329), .Y(n_328) );
AOI222xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_317), .B1(n_320), .B2(n_323), .C1(n_325), .C2(n_326), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_312), .B(n_314), .Y(n_311) );
INVx1_ASAP7_75t_L g393 ( .A(n_312), .Y(n_393) );
INVx1_ASAP7_75t_L g415 ( .A(n_315), .Y(n_415) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_318), .A2(n_429), .B1(n_431), .B2(n_432), .Y(n_428) );
INVx1_ASAP7_75t_L g334 ( .A(n_319), .Y(n_334) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_331), .B1(n_333), .B2(n_335), .C(n_338), .Y(n_327) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g372 ( .A(n_330), .B(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g424 ( .A(n_330), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g399 ( .A(n_335), .Y(n_399) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx1_ASAP7_75t_L g363 ( .A(n_336), .Y(n_363) );
INVx1_ASAP7_75t_L g345 ( .A(n_337), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_340), .B(n_427), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_346), .B1(n_349), .B2(n_350), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g436 ( .A(n_349), .Y(n_436) );
INVxp33_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_351), .B(n_395), .Y(n_394) );
OAI32xp33_ASAP7_75t_L g385 ( .A1(n_352), .A2(n_386), .A3(n_387), .B1(n_388), .B2(n_389), .Y(n_385) );
NAND4xp25_ASAP7_75t_L g353 ( .A(n_354), .B(n_366), .C(n_378), .D(n_390), .Y(n_353) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
NAND2xp33_ASAP7_75t_SL g357 ( .A(n_358), .B(n_359), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_361), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
CKINVDCx16_ASAP7_75t_R g371 ( .A(n_372), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_375), .A2(n_391), .B1(n_408), .B2(n_411), .C(n_412), .Y(n_407) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g426 ( .A(n_377), .B(n_427), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .B1(n_382), .B2(n_384), .C(n_385), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_387), .B(n_418), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B(n_394), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND4xp25_ASAP7_75t_L g396 ( .A(n_397), .B(n_407), .C(n_422), .D(n_433), .Y(n_396) );
O2A1O1Ixp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_401), .B(n_403), .C(n_405), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g438 ( .A(n_425), .Y(n_438) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI21xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_437), .B(n_438), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_SL g446 ( .A(n_441), .B(n_447), .Y(n_446) );
NOR2x2_ASAP7_75t_L g744 ( .A(n_442), .B(n_456), .Y(n_744) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g455 ( .A(n_443), .B(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
OAI222xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_733), .B1(n_736), .B2(n_742), .C1(n_743), .C2(n_745), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_453), .B1(n_454), .B2(n_457), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g739 ( .A(n_452), .Y(n_739) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx6_ASAP7_75t_L g740 ( .A(n_455), .Y(n_740) );
INVx3_ASAP7_75t_L g741 ( .A(n_457), .Y(n_741) );
AND2x2_ASAP7_75t_SL g457 ( .A(n_458), .B(n_688), .Y(n_457) );
NOR4xp25_ASAP7_75t_L g458 ( .A(n_459), .B(n_625), .C(n_659), .D(n_675), .Y(n_458) );
NAND4xp25_ASAP7_75t_SL g459 ( .A(n_460), .B(n_554), .C(n_589), .D(n_605), .Y(n_459) );
AOI222xp33_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_495), .B1(n_529), .B2(n_542), .C1(n_547), .C2(n_553), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AOI31xp33_ASAP7_75t_L g721 ( .A1(n_462), .A2(n_722), .A3(n_723), .B(n_725), .Y(n_721) );
OR2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_474), .Y(n_462) );
AND2x2_ASAP7_75t_L g696 ( .A(n_463), .B(n_476), .Y(n_696) );
BUFx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_SL g546 ( .A(n_464), .Y(n_546) );
AND2x2_ASAP7_75t_L g553 ( .A(n_464), .B(n_486), .Y(n_553) );
AND2x2_ASAP7_75t_L g610 ( .A(n_464), .B(n_477), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_474), .B(n_640), .Y(n_639) );
INVx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_475), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_475), .B(n_557), .Y(n_600) );
AND2x2_ASAP7_75t_L g693 ( .A(n_475), .B(n_633), .Y(n_693) );
OAI321xp33_ASAP7_75t_L g727 ( .A1(n_475), .A2(n_546), .A3(n_700), .B1(n_728), .B2(n_730), .C(n_731), .Y(n_727) );
NAND4xp25_ASAP7_75t_L g731 ( .A(n_475), .B(n_532), .C(n_640), .D(n_732), .Y(n_731) );
AND2x4_ASAP7_75t_L g475 ( .A(n_476), .B(n_486), .Y(n_475) );
AND2x2_ASAP7_75t_L g595 ( .A(n_476), .B(n_544), .Y(n_595) );
AND2x2_ASAP7_75t_L g614 ( .A(n_476), .B(n_546), .Y(n_614) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g545 ( .A(n_477), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g570 ( .A(n_477), .B(n_486), .Y(n_570) );
AND2x2_ASAP7_75t_L g656 ( .A(n_477), .B(n_544), .Y(n_656) );
INVx3_ASAP7_75t_SL g544 ( .A(n_486), .Y(n_544) );
AND2x2_ASAP7_75t_L g588 ( .A(n_486), .B(n_575), .Y(n_588) );
OR2x2_ASAP7_75t_L g621 ( .A(n_486), .B(n_546), .Y(n_621) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_486), .Y(n_628) );
AND2x2_ASAP7_75t_L g657 ( .A(n_486), .B(n_545), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_486), .B(n_630), .Y(n_672) );
AND2x2_ASAP7_75t_L g704 ( .A(n_486), .B(n_696), .Y(n_704) );
AND2x2_ASAP7_75t_L g713 ( .A(n_486), .B(n_558), .Y(n_713) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_493), .Y(n_486) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_508), .Y(n_496) );
INVx1_ASAP7_75t_SL g681 ( .A(n_497), .Y(n_681) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g549 ( .A(n_498), .B(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g531 ( .A(n_499), .B(n_510), .Y(n_531) );
AND2x2_ASAP7_75t_L g617 ( .A(n_499), .B(n_533), .Y(n_617) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g587 ( .A(n_500), .B(n_520), .Y(n_587) );
OR2x2_ASAP7_75t_L g598 ( .A(n_500), .B(n_533), .Y(n_598) );
AND2x2_ASAP7_75t_L g624 ( .A(n_500), .B(n_533), .Y(n_624) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_500), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_508), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_508), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g597 ( .A(n_509), .B(n_598), .Y(n_597) );
AOI322xp5_ASAP7_75t_L g683 ( .A1(n_509), .A2(n_587), .A3(n_593), .B1(n_624), .B2(n_674), .C1(n_684), .C2(n_686), .Y(n_683) );
OR2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_520), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_510), .B(n_532), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_510), .B(n_533), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_510), .B(n_550), .Y(n_604) );
AND2x2_ASAP7_75t_L g658 ( .A(n_510), .B(n_624), .Y(n_658) );
INVx1_ASAP7_75t_L g662 ( .A(n_510), .Y(n_662) );
AND2x2_ASAP7_75t_L g674 ( .A(n_510), .B(n_520), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_510), .B(n_549), .Y(n_706) );
INVx4_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g571 ( .A(n_511), .B(n_520), .Y(n_571) );
BUFx3_ASAP7_75t_L g585 ( .A(n_511), .Y(n_585) );
AND3x2_ASAP7_75t_L g667 ( .A(n_511), .B(n_647), .C(n_668), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g530 ( .A(n_520), .B(n_531), .C(n_532), .Y(n_530) );
INVx1_ASAP7_75t_SL g550 ( .A(n_520), .Y(n_550) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_520), .Y(n_652) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g646 ( .A(n_531), .B(n_647), .Y(n_646) );
INVxp67_ASAP7_75t_L g653 ( .A(n_531), .Y(n_653) );
AND2x2_ASAP7_75t_L g691 ( .A(n_532), .B(n_669), .Y(n_691) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx3_ASAP7_75t_L g572 ( .A(n_533), .Y(n_572) );
AND2x2_ASAP7_75t_L g647 ( .A(n_533), .B(n_550), .Y(n_647) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
OR2x2_ASAP7_75t_L g591 ( .A(n_544), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g710 ( .A(n_544), .B(n_610), .Y(n_710) );
AND2x2_ASAP7_75t_L g724 ( .A(n_544), .B(n_546), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_545), .B(n_558), .Y(n_665) );
AND2x2_ASAP7_75t_L g712 ( .A(n_545), .B(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g575 ( .A(n_546), .B(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g592 ( .A(n_546), .B(n_558), .Y(n_592) );
INVx1_ASAP7_75t_L g602 ( .A(n_546), .Y(n_602) );
AND2x2_ASAP7_75t_L g633 ( .A(n_546), .B(n_558), .Y(n_633) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OAI221xp5_ASAP7_75t_L g675 ( .A1(n_548), .A2(n_676), .B1(n_680), .B2(n_682), .C(n_683), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_549), .B(n_551), .Y(n_548) );
AND2x2_ASAP7_75t_L g579 ( .A(n_549), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_552), .B(n_586), .Y(n_729) );
AOI322xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_571), .A3(n_572), .B1(n_573), .B2(n_579), .C1(n_581), .C2(n_588), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_570), .Y(n_556) );
NAND2x1p5_ASAP7_75t_L g609 ( .A(n_557), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_557), .B(n_620), .Y(n_619) );
O2A1O1Ixp33_ASAP7_75t_L g643 ( .A1(n_557), .A2(n_570), .B(n_644), .C(n_645), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_557), .B(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_557), .B(n_614), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_557), .B(n_696), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_557), .B(n_724), .Y(n_723) );
BUFx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_558), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_558), .B(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g685 ( .A(n_558), .B(n_572), .Y(n_685) );
OA21x2_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_562), .B(n_569), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AO21x2_ASAP7_75t_L g576 ( .A1(n_560), .A2(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g577 ( .A(n_562), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_569), .Y(n_578) );
INVx1_ASAP7_75t_L g660 ( .A(n_570), .Y(n_660) );
OAI31xp33_ASAP7_75t_L g670 ( .A1(n_570), .A2(n_595), .A3(n_671), .B(n_673), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_570), .B(n_576), .Y(n_722) );
INVx1_ASAP7_75t_SL g583 ( .A(n_571), .Y(n_583) );
AND2x2_ASAP7_75t_L g616 ( .A(n_571), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g697 ( .A(n_571), .B(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g582 ( .A(n_572), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g607 ( .A(n_572), .Y(n_607) );
AND2x2_ASAP7_75t_L g634 ( .A(n_572), .B(n_587), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_572), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g726 ( .A(n_572), .B(n_674), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_574), .B(n_644), .Y(n_717) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g613 ( .A(n_576), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g631 ( .A(n_576), .Y(n_631) );
NAND2xp33_ASAP7_75t_SL g581 ( .A(n_582), .B(n_584), .Y(n_581) );
OAI211xp5_ASAP7_75t_SL g625 ( .A1(n_583), .A2(n_626), .B(n_632), .C(n_648), .Y(n_625) );
OR2x2_ASAP7_75t_L g700 ( .A(n_583), .B(n_681), .Y(n_700) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
CKINVDCx16_ASAP7_75t_R g637 ( .A(n_585), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_585), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g606 ( .A(n_587), .B(n_607), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_593), .B(n_596), .C(n_599), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_SL g640 ( .A(n_592), .Y(n_640) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_595), .B(n_633), .Y(n_638) );
INVx1_ASAP7_75t_L g644 ( .A(n_595), .Y(n_644) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g603 ( .A(n_598), .B(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g636 ( .A(n_598), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g698 ( .A(n_598), .Y(n_698) );
AOI21xp33_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_601), .B(n_603), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_601), .A2(n_612), .B(n_615), .Y(n_611) );
AOI211xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_608), .B(n_611), .C(n_618), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_606), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_609), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_SL g622 ( .A(n_610), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g677 ( .A1(n_612), .A2(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_617), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g642 ( .A(n_617), .Y(n_642) );
AOI21xp33_ASAP7_75t_SL g618 ( .A1(n_619), .A2(n_622), .B(n_623), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g673 ( .A(n_624), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_630), .B(n_656), .Y(n_682) );
AND2x2_ASAP7_75t_L g695 ( .A(n_630), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g709 ( .A(n_630), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g719 ( .A(n_630), .B(n_657), .Y(n_719) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI211xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B(n_635), .C(n_643), .Y(n_632) );
INVx1_ASAP7_75t_L g679 ( .A(n_633), .Y(n_679) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .B1(n_639), .B2(n_641), .Y(n_635) );
OR2x2_ASAP7_75t_L g641 ( .A(n_637), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_637), .B(n_698), .Y(n_720) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g714 ( .A(n_647), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_654), .B1(n_657), .B2(n_658), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g732 ( .A(n_652), .Y(n_732) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g678 ( .A(n_656), .Y(n_678) );
OAI211xp5_ASAP7_75t_SL g659 ( .A1(n_660), .A2(n_661), .B(n_663), .C(n_670), .Y(n_659) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVxp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVxp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_678), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NOR5xp2_ASAP7_75t_L g688 ( .A(n_689), .B(n_707), .C(n_715), .D(n_721), .E(n_727), .Y(n_688) );
OAI211xp5_ASAP7_75t_SL g689 ( .A1(n_690), .A2(n_692), .B(n_694), .C(n_701), .Y(n_689) );
INVxp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_697), .B(n_699), .Y(n_694) );
OAI21xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_704), .B(n_705), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_704), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI21xp33_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_711), .B(n_714), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g730 ( .A(n_710), .Y(n_730) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_718), .B(n_720), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
CKINVDCx16_ASAP7_75t_R g742 ( .A(n_733), .Y(n_742) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx3_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
endmodule