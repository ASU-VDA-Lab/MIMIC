module fake_jpeg_30308_n_104 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_9),
.B(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_50),
.Y(n_54)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_48),
.Y(n_60)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_0),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_17),
.C(n_31),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_0),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_59),
.B(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_42),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_41),
.B1(n_40),
.B2(n_39),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_75),
.B(n_74),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_18),
.B1(n_30),
.B2(n_29),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_72),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_14),
.B1(n_27),
.B2(n_26),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_12),
.B1(n_23),
.B2(n_22),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_8),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_76),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_1),
.Y(n_76)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_16),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_6),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_4),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_84),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_85),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_5),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_32),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_78),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_96),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_78),
.B1(n_79),
.B2(n_20),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_97),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_95),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_90),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_92),
.Y(n_102)
);

BUFx24_ASAP7_75t_SL g103 ( 
.A(n_102),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_21),
.Y(n_104)
);


endmodule