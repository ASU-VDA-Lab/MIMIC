module fake_jpeg_27379_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_5),
.B(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_36),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_0),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_13),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_44),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_21),
.B1(n_25),
.B2(n_22),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_30),
.B1(n_31),
.B2(n_28),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_22),
.B1(n_21),
.B2(n_25),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_30),
.B1(n_20),
.B2(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_14),
.Y(n_44)
);

AND2x4_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_22),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_33),
.B(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_50),
.Y(n_78)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_23),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_63),
.Y(n_70)
);

MAJx2_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_33),
.C(n_36),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_65),
.C(n_61),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_16),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_47),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_37),
.B(n_33),
.Y(n_67)
);

OA21x2_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_75),
.B(n_52),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_65),
.Y(n_86)
);

OA22x2_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_33),
.B1(n_40),
.B2(n_32),
.Y(n_75)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_44),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_58),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_16),
.C(n_15),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_19),
.C(n_24),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_48),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_81),
.B(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_90),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_92),
.C(n_94),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_55),
.B1(n_51),
.B2(n_63),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_91),
.B(n_93),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_73),
.A2(n_51),
.B1(n_62),
.B2(n_59),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_77),
.B1(n_75),
.B2(n_82),
.Y(n_104)
);

NOR2xp67_ASAP7_75t_SL g93 ( 
.A(n_70),
.B(n_18),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_64),
.C(n_56),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_67),
.C(n_71),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_15),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_91),
.A2(n_74),
.B(n_78),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_102),
.B(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_101),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_74),
.B(n_68),
.Y(n_102)
);

A2O1A1O1Ixp25_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_75),
.B(n_68),
.C(n_27),
.D(n_18),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_96),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_1),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_101),
.A2(n_19),
.B1(n_92),
.B2(n_66),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_109),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_76),
.C(n_66),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_76),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_98),
.B(n_105),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_112),
.C(n_114),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_106),
.B1(n_27),
.B2(n_17),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_17),
.B1(n_12),
.B2(n_11),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_123),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_115),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_110),
.C(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_125),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_120),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_115),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_129),
.Y(n_130)
);

AOI322xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_118),
.A3(n_9),
.B1(n_8),
.B2(n_4),
.C1(n_1),
.C2(n_6),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.C(n_2),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_5),
.C1(n_8),
.C2(n_128),
.Y(n_132)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_133),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_2),
.C(n_5),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_134),
.Y(n_136)
);


endmodule