module fake_ariane_581_n_2775 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_598, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_238, n_365, n_429, n_455, n_588, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_2775);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_588;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_2775;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_1298;
wire n_737;
wire n_2653;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_1761;
wire n_829;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2233;
wire n_2370;
wire n_2663;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2620;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1253;
wire n_1468;
wire n_762;
wire n_1661;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_2745;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_2628;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2662;
wire n_1259;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2599;
wire n_727;
wire n_699;
wire n_2075;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_957;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_845;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2525;
wire n_1815;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2613;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_683;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1588;
wire n_1148;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_723;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2275;
wire n_2205;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_447),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_152),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_549),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_590),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_305),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_270),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_297),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_18),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_498),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_263),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_235),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_230),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_351),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_567),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_273),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_41),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_572),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_282),
.Y(n_623)
);

BUFx10_ASAP7_75t_L g624 ( 
.A(n_222),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_449),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_212),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_505),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_290),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_101),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_501),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_571),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_497),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_77),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_414),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_411),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_492),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_579),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_439),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_504),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_584),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_237),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_582),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_64),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_404),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_503),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_509),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_482),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_292),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_576),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_435),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_188),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_264),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_442),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_133),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_458),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_574),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_131),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_339),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_312),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_603),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_275),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_477),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_56),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_577),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_95),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_87),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_139),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_44),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_294),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_472),
.Y(n_670)
);

BUFx8_ASAP7_75t_SL g671 ( 
.A(n_527),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_563),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_499),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_561),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_233),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_484),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_256),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_300),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_320),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_177),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_505),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_493),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_104),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_416),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_479),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_338),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_322),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_192),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_365),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_382),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_288),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_80),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_526),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_437),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_460),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_136),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_445),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_512),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_502),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_498),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_347),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_510),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_414),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_588),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_464),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_359),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_281),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_65),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_431),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_149),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_377),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_566),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_231),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_283),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_112),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_318),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_500),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_190),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_8),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_288),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_417),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_234),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_205),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_605),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_431),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_511),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_89),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_249),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_165),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_488),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_167),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_171),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_508),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_363),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_242),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_294),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_321),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_490),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_591),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_550),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_436),
.Y(n_741)
);

INVx1_ASAP7_75t_SL g742 ( 
.A(n_105),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_75),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_282),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_78),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_514),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_224),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_544),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_49),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_286),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_23),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_569),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_424),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_72),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_333),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_314),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_35),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_1),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_425),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_119),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_478),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_304),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_266),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_270),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_120),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_352),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_211),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_228),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_390),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_441),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_125),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_436),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_146),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_280),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_525),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_0),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_102),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_390),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_365),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_366),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_166),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_20),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_487),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_587),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_181),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_322),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_597),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_97),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_305),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_272),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_26),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_374),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_0),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_31),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_470),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_104),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_445),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_44),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_149),
.Y(n_799)
);

BUFx10_ASAP7_75t_L g800 ( 
.A(n_362),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_496),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_60),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_137),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_494),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_138),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_114),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_509),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_140),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_53),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_86),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_554),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_10),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_492),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_131),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_135),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_233),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_271),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_203),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_292),
.Y(n_819)
);

INVx1_ASAP7_75t_SL g820 ( 
.A(n_83),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_334),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_461),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_507),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_235),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_331),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_218),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_18),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_260),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_276),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_364),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_310),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_188),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_103),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_332),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_506),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_5),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_133),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_125),
.Y(n_838)
);

BUFx10_ASAP7_75t_L g839 ( 
.A(n_424),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_317),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_118),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_495),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_158),
.Y(n_843)
);

BUFx5_ASAP7_75t_L g844 ( 
.A(n_29),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_513),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_480),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_48),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_306),
.Y(n_848)
);

CKINVDCx14_ASAP7_75t_R g849 ( 
.A(n_450),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_844),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_844),
.Y(n_851)
);

CKINVDCx20_ASAP7_75t_R g852 ( 
.A(n_629),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_629),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_643),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_620),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_615),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_615),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_617),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_617),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_641),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_646),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_844),
.Y(n_862)
);

CKINVDCx16_ASAP7_75t_R g863 ( 
.A(n_849),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_844),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_844),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_608),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_844),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_844),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_693),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_628),
.Y(n_870)
);

CKINVDCx16_ASAP7_75t_R g871 ( 
.A(n_624),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_628),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_628),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_628),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_669),
.B(n_1),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_734),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_641),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_612),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_746),
.Y(n_879)
);

INVxp33_ASAP7_75t_SL g880 ( 
.A(n_650),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_628),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_638),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_638),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_638),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_631),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_631),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_638),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_659),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_643),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_659),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_673),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_673),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_638),
.Y(n_893)
);

INVxp33_ASAP7_75t_L g894 ( 
.A(n_680),
.Y(n_894)
);

CKINVDCx16_ASAP7_75t_R g895 ( 
.A(n_624),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_681),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_681),
.Y(n_897)
);

INVxp67_ASAP7_75t_SL g898 ( 
.A(n_707),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_707),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_764),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_796),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_619),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_796),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_748),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_806),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_752),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_806),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_611),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_613),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_637),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_618),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_625),
.Y(n_912)
);

CKINVDCx16_ASAP7_75t_R g913 ( 
.A(n_624),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_626),
.Y(n_914)
);

NOR2xp67_ASAP7_75t_L g915 ( 
.A(n_675),
.B(n_2),
.Y(n_915)
);

INVxp67_ASAP7_75t_SL g916 ( 
.A(n_645),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_633),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_644),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_647),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_648),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_645),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_652),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_668),
.Y(n_923)
);

INVxp33_ASAP7_75t_L g924 ( 
.A(n_770),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_800),
.B(n_2),
.Y(n_925)
);

CKINVDCx16_ASAP7_75t_R g926 ( 
.A(n_800),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_684),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_691),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_652),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_692),
.Y(n_930)
);

INVxp67_ASAP7_75t_SL g931 ( 
.A(n_645),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_695),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_696),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_697),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_700),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_702),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_703),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_706),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_708),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_645),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_645),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_658),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_658),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_658),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_752),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_658),
.Y(n_946)
);

INVxp67_ASAP7_75t_SL g947 ( 
.A(n_683),
.Y(n_947)
);

INVxp33_ASAP7_75t_SL g948 ( 
.A(n_622),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_683),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_748),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_683),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_711),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_916),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_948),
.B(n_672),
.Y(n_954)
);

INVx5_ASAP7_75t_L g955 ( 
.A(n_904),
.Y(n_955)
);

BUFx12f_ASAP7_75t_L g956 ( 
.A(n_885),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_902),
.B(n_675),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_877),
.B(n_712),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_898),
.B(n_811),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_904),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_931),
.B(n_609),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_948),
.B(n_915),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_856),
.B(n_857),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_904),
.Y(n_964)
);

CKINVDCx6p67_ASAP7_75t_R g965 ( 
.A(n_863),
.Y(n_965)
);

BUFx8_ASAP7_75t_L g966 ( 
.A(n_925),
.Y(n_966)
);

BUFx12f_ASAP7_75t_L g967 ( 
.A(n_885),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_947),
.B(n_609),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_922),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_902),
.B(n_649),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_SL g971 ( 
.A(n_871),
.B(n_671),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_910),
.B(n_790),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_850),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_910),
.B(n_649),
.Y(n_974)
);

BUFx12f_ASAP7_75t_L g975 ( 
.A(n_886),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_879),
.B(n_640),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_879),
.B(n_640),
.Y(n_977)
);

INVx5_ASAP7_75t_L g978 ( 
.A(n_904),
.Y(n_978)
);

INVx5_ASAP7_75t_L g979 ( 
.A(n_904),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_886),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_866),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_925),
.B(n_790),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_950),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_906),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_874),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_874),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_858),
.B(n_800),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_866),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_906),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_850),
.Y(n_990)
);

INVx5_ASAP7_75t_L g991 ( 
.A(n_950),
.Y(n_991)
);

BUFx12f_ASAP7_75t_L g992 ( 
.A(n_945),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_875),
.B(n_848),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_875),
.B(n_848),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_859),
.B(n_663),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_945),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_851),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_SL g998 ( 
.A(n_895),
.B(n_666),
.Y(n_998)
);

INVx5_ASAP7_75t_L g999 ( 
.A(n_950),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_860),
.B(n_888),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_SL g1001 ( 
.A(n_913),
.B(n_666),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_950),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_950),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_890),
.B(n_663),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_869),
.B(n_642),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_891),
.B(n_656),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_869),
.B(n_642),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_893),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_893),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_892),
.B(n_701),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_896),
.B(n_660),
.Y(n_1011)
);

INVx5_ASAP7_75t_L g1012 ( 
.A(n_921),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_941),
.Y(n_1013)
);

INVxp67_ASAP7_75t_L g1014 ( 
.A(n_878),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_897),
.B(n_664),
.Y(n_1015)
);

INVx2_ASAP7_75t_SL g1016 ( 
.A(n_899),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_901),
.B(n_674),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_SL g1018 ( 
.A(n_926),
.B(n_729),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_851),
.Y(n_1019)
);

NAND2x1_ASAP7_75t_L g1020 ( 
.A(n_990),
.B(n_921),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_1008),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_973),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_973),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_997),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_997),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_985),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1019),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_953),
.B(n_862),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_985),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_986),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_986),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1013),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_982),
.B(n_894),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_954),
.B(n_862),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_1008),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_987),
.B(n_864),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_1006),
.A2(n_865),
.B(n_864),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_1008),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_987),
.B(n_903),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_976),
.B(n_865),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1013),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_961),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1008),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_1008),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_977),
.B(n_867),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_968),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_982),
.A2(n_880),
.B1(n_729),
.B2(n_689),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1009),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_1009),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_1009),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1009),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1009),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_960),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1012),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_960),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1012),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1012),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_982),
.B(n_924),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1012),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_1005),
.B(n_880),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1012),
.Y(n_1061)
);

INVx5_ASAP7_75t_L g1062 ( 
.A(n_960),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_969),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_970),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_960),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_960),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_SL g1067 ( 
.A(n_971),
.B(n_677),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_964),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_974),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_964),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_964),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_993),
.B(n_867),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_964),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_964),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_963),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_983),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_963),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_965),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_983),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1000),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1016),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1016),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_993),
.B(n_994),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_957),
.B(n_972),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_983),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_983),
.Y(n_1086)
);

AND3x2_ASAP7_75t_L g1087 ( 
.A(n_998),
.B(n_861),
.C(n_855),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_983),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_1007),
.B(n_962),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1002),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1002),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_981),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_1002),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_957),
.B(n_905),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_993),
.B(n_907),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1002),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_981),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1002),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1003),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1003),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1003),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1003),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1003),
.Y(n_1103)
);

AND2x6_ASAP7_75t_L g1104 ( 
.A(n_994),
.B(n_748),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_955),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_955),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_955),
.Y(n_1107)
);

NAND2xp33_ASAP7_75t_L g1108 ( 
.A(n_988),
.B(n_683),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1034),
.B(n_988),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1029),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_1044),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_1104),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1033),
.B(n_957),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_1092),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1026),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1026),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_1089),
.B(n_962),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1064),
.B(n_994),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_1092),
.B(n_1014),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1060),
.A2(n_1011),
.B1(n_1017),
.B2(n_1015),
.Y(n_1120)
);

INVxp67_ASAP7_75t_SL g1121 ( 
.A(n_1063),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1030),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1029),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1031),
.Y(n_1124)
);

BUFx8_ASAP7_75t_SL g1125 ( 
.A(n_1078),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1033),
.B(n_972),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1031),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_1064),
.B(n_989),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1030),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1027),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1081),
.B(n_972),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_1097),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1069),
.B(n_1080),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1032),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1041),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1041),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1032),
.Y(n_1137)
);

NAND3xp33_ASAP7_75t_L g1138 ( 
.A(n_1080),
.B(n_984),
.C(n_980),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1069),
.B(n_958),
.Y(n_1139)
);

NAND2xp33_ASAP7_75t_R g1140 ( 
.A(n_1087),
.B(n_965),
.Y(n_1140)
);

INVx4_ASAP7_75t_L g1141 ( 
.A(n_1021),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1027),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1022),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1042),
.B(n_959),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1022),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1024),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1024),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1023),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1081),
.B(n_966),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1023),
.Y(n_1150)
);

AND2x6_ASAP7_75t_L g1151 ( 
.A(n_1084),
.B(n_748),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1025),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_1025),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1082),
.B(n_996),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1075),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1075),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1043),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1077),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_1058),
.Y(n_1159)
);

INVx4_ASAP7_75t_L g1160 ( 
.A(n_1021),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1042),
.B(n_966),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_1104),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1082),
.B(n_966),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1021),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1042),
.B(n_876),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1077),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1043),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1028),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1072),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1020),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1047),
.B(n_900),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1048),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1020),
.Y(n_1173)
);

INVx2_ASAP7_75t_SL g1174 ( 
.A(n_1104),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1104),
.A2(n_689),
.B1(n_728),
.B2(n_677),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1084),
.B(n_1001),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1104),
.A2(n_754),
.B1(n_818),
.B2(n_728),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_1047),
.B(n_1004),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1048),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1039),
.B(n_1018),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1039),
.B(n_956),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1094),
.Y(n_1182)
);

INVxp67_ASAP7_75t_L g1183 ( 
.A(n_1058),
.Y(n_1183)
);

AO21x2_ASAP7_75t_L g1184 ( 
.A1(n_1037),
.A2(n_872),
.B(n_870),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1050),
.Y(n_1185)
);

CKINVDCx6p67_ASAP7_75t_R g1186 ( 
.A(n_1104),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1050),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1066),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1051),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1066),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1036),
.B(n_956),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1068),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1095),
.B(n_995),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_1039),
.B(n_967),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1044),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1039),
.B(n_967),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1083),
.B(n_975),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1040),
.B(n_975),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1068),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1094),
.B(n_995),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1071),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1104),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1046),
.B(n_995),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1071),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1079),
.Y(n_1205)
);

INVx8_ASAP7_75t_L g1206 ( 
.A(n_1095),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1044),
.Y(n_1207)
);

AO21x2_ASAP7_75t_L g1208 ( 
.A1(n_1037),
.A2(n_872),
.B(n_870),
.Y(n_1208)
);

INVxp67_ASAP7_75t_SL g1209 ( 
.A(n_1021),
.Y(n_1209)
);

INVxp67_ASAP7_75t_R g1210 ( 
.A(n_1067),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1046),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1046),
.B(n_1004),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1079),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1095),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1051),
.Y(n_1215)
);

NAND2xp33_ASAP7_75t_L g1216 ( 
.A(n_1045),
.B(n_683),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1095),
.Y(n_1217)
);

CKINVDCx6p67_ASAP7_75t_R g1218 ( 
.A(n_1062),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1088),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1021),
.B(n_992),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1108),
.A2(n_818),
.B1(n_824),
.B2(n_754),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1088),
.Y(n_1222)
);

INVx4_ASAP7_75t_L g1223 ( 
.A(n_1021),
.Y(n_1223)
);

NAND3xp33_ASAP7_75t_L g1224 ( 
.A(n_1052),
.B(n_627),
.C(n_606),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1090),
.Y(n_1225)
);

NAND2xp33_ASAP7_75t_L g1226 ( 
.A(n_1053),
.B(n_771),
.Y(n_1226)
);

AND2x6_ASAP7_75t_L g1227 ( 
.A(n_1054),
.B(n_748),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1035),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1049),
.B(n_1004),
.Y(n_1229)
);

BUFx10_ASAP7_75t_L g1230 ( 
.A(n_1035),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1049),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1052),
.A2(n_824),
.B1(n_1010),
.B2(n_676),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1090),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1054),
.Y(n_1234)
);

NAND2xp33_ASAP7_75t_L g1235 ( 
.A(n_1053),
.B(n_1055),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1035),
.B(n_1038),
.Y(n_1236)
);

NAND2xp33_ASAP7_75t_L g1237 ( 
.A(n_1053),
.B(n_1055),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1099),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1049),
.B(n_1010),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1049),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1070),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1056),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1099),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1085),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1056),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1142),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1142),
.Y(n_1247)
);

INVxp67_ASAP7_75t_SL g1248 ( 
.A(n_1164),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1159),
.B(n_992),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1130),
.Y(n_1250)
);

CKINVDCx16_ASAP7_75t_R g1251 ( 
.A(n_1140),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1143),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1119),
.B(n_852),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1143),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1110),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1110),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1123),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1109),
.B(n_1070),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1133),
.A2(n_1237),
.B(n_1235),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1114),
.Y(n_1260)
);

XOR2xp5_ASAP7_75t_L g1261 ( 
.A(n_1119),
.B(n_852),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1124),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1124),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1115),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1125),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1127),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1127),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1164),
.Y(n_1268)
);

NOR2xp67_ASAP7_75t_L g1269 ( 
.A(n_1138),
.B(n_1010),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1135),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1135),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1115),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1136),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1136),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1155),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1183),
.B(n_1070),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1193),
.B(n_1214),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1168),
.B(n_1070),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1171),
.B(n_853),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1156),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1117),
.B(n_1128),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1169),
.B(n_1035),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1158),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1166),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1239),
.Y(n_1285)
);

CKINVDCx16_ASAP7_75t_R g1286 ( 
.A(n_1175),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1239),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1145),
.Y(n_1288)
);

NAND2xp33_ASAP7_75t_R g1289 ( 
.A(n_1191),
.B(n_853),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1146),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1193),
.B(n_908),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1125),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1165),
.B(n_1057),
.Y(n_1293)
);

NOR2xp67_ASAP7_75t_L g1294 ( 
.A(n_1132),
.B(n_909),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1234),
.A2(n_1091),
.B(n_1085),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1176),
.B(n_1057),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1147),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1229),
.Y(n_1298)
);

XNOR2x2_ASAP7_75t_L g1299 ( 
.A(n_1177),
.B(n_854),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1148),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1113),
.B(n_854),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1113),
.B(n_1126),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1234),
.A2(n_1096),
.B(n_1091),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1217),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1193),
.B(n_911),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1126),
.B(n_889),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1116),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1171),
.B(n_889),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1189),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1154),
.B(n_1059),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1189),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1215),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1215),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1211),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1150),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1150),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1153),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1152),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1121),
.B(n_929),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1152),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1153),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1116),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1203),
.Y(n_1323)
);

XOR2xp5_ASAP7_75t_L g1324 ( 
.A(n_1221),
.B(n_929),
.Y(n_1324)
);

CKINVDCx11_ASAP7_75t_R g1325 ( 
.A(n_1206),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1212),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1182),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1139),
.B(n_1059),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1200),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1144),
.B(n_1035),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1200),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1242),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1180),
.B(n_1061),
.Y(n_1333)
);

XOR2x2_ASAP7_75t_L g1334 ( 
.A(n_1198),
.B(n_820),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1242),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1245),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_1181),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1245),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1122),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1129),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1129),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1120),
.B(n_1061),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1134),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1134),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1137),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1206),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1137),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1244),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1244),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1157),
.Y(n_1350)
);

INVxp33_ASAP7_75t_L g1351 ( 
.A(n_1178),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1206),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1210),
.B(n_912),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1178),
.B(n_1096),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1118),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1206),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1131),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1161),
.B(n_1035),
.Y(n_1358)
);

XNOR2x2_ASAP7_75t_L g1359 ( 
.A(n_1210),
.B(n_630),
.Y(n_1359)
);

XNOR2xp5_ASAP7_75t_L g1360 ( 
.A(n_1194),
.B(n_914),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1167),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1167),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_SL g1363 ( 
.A(n_1186),
.B(n_742),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1197),
.B(n_1098),
.Y(n_1364)
);

INVx1_ASAP7_75t_SL g1365 ( 
.A(n_1196),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1232),
.B(n_917),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1172),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1172),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1179),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1179),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1149),
.B(n_918),
.Y(n_1371)
);

AND2x2_ASAP7_75t_SL g1372 ( 
.A(n_1235),
.B(n_771),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1163),
.B(n_1220),
.Y(n_1373)
);

NAND2x1p5_ASAP7_75t_L g1374 ( 
.A(n_1170),
.B(n_1038),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1185),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1185),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1111),
.B(n_1098),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1187),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1187),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1111),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1111),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1195),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1188),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1195),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1170),
.B(n_919),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1188),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_1186),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1195),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1240),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1240),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1240),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1190),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_1228),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1230),
.Y(n_1394)
);

NAND2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1112),
.B(n_1038),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1190),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1192),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1207),
.B(n_920),
.Y(n_1398)
);

INVxp33_ASAP7_75t_L g1399 ( 
.A(n_1224),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1228),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1192),
.Y(n_1401)
);

INVxp33_ASAP7_75t_L g1402 ( 
.A(n_1243),
.Y(n_1402)
);

INVxp33_ASAP7_75t_SL g1403 ( 
.A(n_1173),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1199),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1218),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1199),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1201),
.Y(n_1407)
);

NOR2xp67_ASAP7_75t_L g1408 ( 
.A(n_1201),
.B(n_923),
.Y(n_1408)
);

XOR2x2_ASAP7_75t_L g1409 ( 
.A(n_1112),
.B(n_747),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1204),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1204),
.Y(n_1411)
);

XNOR2xp5_ASAP7_75t_L g1412 ( 
.A(n_1162),
.B(n_927),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1205),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1205),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1213),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_SL g1416 ( 
.A(n_1162),
.B(n_830),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1213),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1218),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1151),
.B(n_1038),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1219),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_SL g1421 ( 
.A(n_1174),
.B(n_841),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1207),
.B(n_1100),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1219),
.Y(n_1423)
);

OAI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1236),
.A2(n_1102),
.B(n_1101),
.Y(n_1424)
);

XNOR2xp5_ASAP7_75t_L g1425 ( 
.A(n_1174),
.B(n_928),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1231),
.Y(n_1426)
);

XOR2xp5_ASAP7_75t_L g1427 ( 
.A(n_1202),
.B(n_606),
.Y(n_1427)
);

OAI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1241),
.A2(n_1209),
.B(n_1222),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1231),
.B(n_1101),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1222),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1164),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1225),
.Y(n_1432)
);

NAND2xp33_ASAP7_75t_R g1433 ( 
.A(n_1225),
.B(n_1105),
.Y(n_1433)
);

NOR2xp67_ASAP7_75t_L g1434 ( 
.A(n_1233),
.B(n_1238),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1233),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1238),
.Y(n_1436)
);

NAND2x1p5_ASAP7_75t_L g1437 ( 
.A(n_1202),
.B(n_1141),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1151),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1151),
.Y(n_1439)
);

XNOR2xp5_ASAP7_75t_L g1440 ( 
.A(n_1184),
.B(n_930),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1250),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1355),
.B(n_1141),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1281),
.B(n_1323),
.Y(n_1443)
);

NAND2xp33_ASAP7_75t_L g1444 ( 
.A(n_1400),
.B(n_1164),
.Y(n_1444)
);

BUFx6f_ASAP7_75t_L g1445 ( 
.A(n_1325),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_R g1446 ( 
.A(n_1405),
.B(n_1151),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1261),
.B(n_1164),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1264),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1260),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1281),
.B(n_1141),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1403),
.B(n_1160),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1275),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1301),
.B(n_839),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1264),
.Y(n_1454)
);

NAND2xp33_ASAP7_75t_L g1455 ( 
.A(n_1268),
.B(n_1394),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1326),
.B(n_1160),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1298),
.B(n_1160),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1354),
.B(n_1223),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1319),
.B(n_1253),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1265),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1286),
.B(n_1223),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1306),
.B(n_839),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1272),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1393),
.B(n_1223),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1289),
.B(n_1216),
.C(n_838),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1272),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1299),
.A2(n_839),
.B1(n_632),
.B2(n_634),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1354),
.B(n_1230),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1280),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1328),
.B(n_1230),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_1325),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1307),
.Y(n_1472)
);

AND2x6_ASAP7_75t_SL g1473 ( 
.A(n_1308),
.B(n_932),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1328),
.B(n_1237),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1307),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1393),
.B(n_1038),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1302),
.B(n_627),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1249),
.B(n_632),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1322),
.Y(n_1479)
);

AO221x1_ASAP7_75t_L g1480 ( 
.A1(n_1289),
.A2(n_783),
.B1(n_785),
.B2(n_781),
.C(n_771),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1337),
.A2(n_1216),
.B1(n_610),
.B2(n_614),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1283),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1277),
.B(n_1038),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_R g1484 ( 
.A(n_1405),
.B(n_1226),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1277),
.B(n_634),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1431),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1279),
.B(n_933),
.Y(n_1487)
);

AOI221xp5_ASAP7_75t_L g1488 ( 
.A1(n_1329),
.A2(n_936),
.B1(n_937),
.B2(n_935),
.C(n_934),
.Y(n_1488)
);

INVx4_ASAP7_75t_L g1489 ( 
.A(n_1426),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1284),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1337),
.A2(n_616),
.B1(n_621),
.B2(n_607),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1427),
.B(n_635),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1331),
.B(n_635),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1351),
.B(n_636),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1324),
.B(n_938),
.Y(n_1495)
);

NAND2xp33_ASAP7_75t_L g1496 ( 
.A(n_1268),
.B(n_1394),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1322),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1255),
.B(n_1184),
.Y(n_1498)
);

INVxp67_ASAP7_75t_L g1499 ( 
.A(n_1353),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1251),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1288),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1290),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1297),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1327),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1351),
.B(n_636),
.Y(n_1505)
);

O2A1O1Ixp5_ASAP7_75t_L g1506 ( 
.A1(n_1259),
.A2(n_1102),
.B(n_1103),
.C(n_1106),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1341),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1291),
.B(n_639),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1341),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1256),
.B(n_1184),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1291),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1365),
.B(n_639),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1350),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1346),
.B(n_727),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1350),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1257),
.B(n_1208),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1399),
.B(n_727),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1300),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1252),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1254),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1399),
.B(n_825),
.Y(n_1521)
);

BUFx5_ASAP7_75t_L g1522 ( 
.A(n_1431),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1305),
.B(n_939),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1305),
.B(n_825),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1352),
.B(n_826),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1262),
.B(n_1208),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1385),
.B(n_952),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1366),
.A2(n_832),
.B1(n_833),
.B2(n_826),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1294),
.B(n_1372),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1360),
.B(n_832),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1342),
.B(n_833),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1363),
.B(n_836),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1263),
.B(n_1266),
.Y(n_1533)
);

NOR2xp67_ASAP7_75t_L g1534 ( 
.A(n_1292),
.B(n_1103),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1267),
.B(n_868),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1398),
.B(n_840),
.Y(n_1536)
);

INVx8_ASAP7_75t_L g1537 ( 
.A(n_1418),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1310),
.B(n_840),
.Y(n_1538)
);

OAI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1259),
.A2(n_868),
.B(n_1226),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1270),
.B(n_1053),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1379),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_SL g1542 ( 
.A(n_1310),
.B(n_843),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1285),
.B(n_843),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_SL g1544 ( 
.A1(n_1412),
.A2(n_846),
.B1(n_847),
.B2(n_845),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1317),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1314),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1287),
.B(n_1425),
.Y(n_1547)
);

INVx8_ASAP7_75t_L g1548 ( 
.A(n_1418),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1356),
.B(n_845),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1387),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1409),
.A2(n_847),
.B1(n_846),
.B2(n_651),
.Y(n_1551)
);

OR2x6_ASAP7_75t_L g1552 ( 
.A(n_1373),
.B(n_1106),
.Y(n_1552)
);

BUFx8_ASAP7_75t_L g1553 ( 
.A(n_1371),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1374),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1342),
.B(n_1053),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1293),
.B(n_623),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1293),
.B(n_653),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1271),
.B(n_654),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1332),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1373),
.B(n_1053),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1371),
.B(n_655),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1383),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1374),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1383),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_1387),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_SL g1566 ( 
.A1(n_1334),
.A2(n_661),
.B1(n_662),
.B2(n_657),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1273),
.B(n_1055),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1274),
.B(n_665),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1386),
.Y(n_1569)
);

OR2x6_ASAP7_75t_SL g1570 ( 
.A(n_1359),
.B(n_667),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1357),
.B(n_670),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1304),
.B(n_678),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1269),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1386),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1335),
.A2(n_720),
.B1(n_750),
.B2(n_701),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1364),
.A2(n_1421),
.B1(n_1416),
.B2(n_1333),
.Y(n_1576)
);

AND2x2_ASAP7_75t_SL g1577 ( 
.A(n_1364),
.B(n_1268),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1343),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1268),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1440),
.Y(n_1580)
);

O2A1O1Ixp5_ASAP7_75t_L g1581 ( 
.A1(n_1258),
.A2(n_761),
.B(n_750),
.C(n_755),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1246),
.B(n_1055),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1247),
.A2(n_682),
.B1(n_685),
.B2(n_679),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1276),
.B(n_1055),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1348),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1309),
.B(n_1055),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1276),
.B(n_1065),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1311),
.B(n_1065),
.Y(n_1588)
);

O2A1O1Ixp5_ASAP7_75t_L g1589 ( 
.A1(n_1258),
.A2(n_755),
.B(n_758),
.C(n_720),
.Y(n_1589)
);

INVx8_ASAP7_75t_L g1590 ( 
.A(n_1433),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1296),
.B(n_686),
.Y(n_1591)
);

INVxp33_ASAP7_75t_L g1592 ( 
.A(n_1333),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1349),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1312),
.B(n_1065),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1313),
.B(n_1065),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1422),
.B(n_1065),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1336),
.B(n_1065),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1339),
.Y(n_1598)
);

OR2x6_ASAP7_75t_L g1599 ( 
.A(n_1438),
.B(n_758),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1340),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1338),
.B(n_1073),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1344),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1345),
.B(n_1073),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1347),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1296),
.B(n_687),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1248),
.B(n_1105),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1315),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1316),
.B(n_1318),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_SL g1609 ( 
.A(n_1248),
.B(n_704),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1320),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1321),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1408),
.B(n_688),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1278),
.B(n_1073),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1361),
.B(n_1073),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1362),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1422),
.B(n_1073),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1380),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1367),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1429),
.B(n_1074),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1368),
.B(n_1074),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1369),
.B(n_1074),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1381),
.B(n_690),
.Y(n_1622)
);

O2A1O1Ixp5_ASAP7_75t_L g1623 ( 
.A1(n_1295),
.A2(n_817),
.B(n_831),
.C(n_761),
.Y(n_1623)
);

O2A1O1Ixp33_ASAP7_75t_L g1624 ( 
.A1(n_1382),
.A2(n_1388),
.B(n_1389),
.C(n_1384),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1370),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1375),
.B(n_1074),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1376),
.B(n_1074),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1429),
.B(n_1076),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1282),
.B(n_694),
.Y(n_1629)
);

NOR2xp67_ASAP7_75t_L g1630 ( 
.A(n_1390),
.B(n_1062),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1378),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1392),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1396),
.B(n_698),
.Y(n_1633)
);

AND2x4_ASAP7_75t_SL g1634 ( 
.A(n_1391),
.B(n_1076),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1433),
.A2(n_705),
.B1(n_709),
.B2(n_699),
.Y(n_1635)
);

OR2x6_ASAP7_75t_L g1636 ( 
.A(n_1437),
.B(n_817),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1402),
.B(n_710),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1437),
.Y(n_1638)
);

INVx5_ASAP7_75t_L g1639 ( 
.A(n_1395),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1474),
.A2(n_1330),
.B(n_1428),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1504),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1531),
.B(n_1397),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1474),
.A2(n_1470),
.B(n_1458),
.Y(n_1643)
);

INVx2_ASAP7_75t_SL g1644 ( 
.A(n_1537),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1451),
.B(n_1358),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1470),
.A2(n_1303),
.B(n_1377),
.Y(n_1646)
);

AOI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1555),
.A2(n_1434),
.B(n_1419),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1585),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1537),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1523),
.B(n_714),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1458),
.A2(n_1468),
.B(n_1450),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1576),
.B(n_1377),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1468),
.A2(n_1424),
.B(n_1395),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1511),
.Y(n_1654)
);

O2A1O1Ixp33_ASAP7_75t_L g1655 ( 
.A1(n_1538),
.A2(n_715),
.B(n_726),
.C(n_713),
.Y(n_1655)
);

AOI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1530),
.A2(n_1439),
.B1(n_717),
.B2(n_718),
.Y(n_1656)
);

NOR2xp67_ASAP7_75t_L g1657 ( 
.A(n_1489),
.B(n_1401),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1443),
.A2(n_831),
.B1(n_736),
.B2(n_763),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1593),
.Y(n_1659)
);

O2A1O1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1591),
.A2(n_776),
.B(n_777),
.C(n_735),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1592),
.B(n_716),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_SL g1662 ( 
.A(n_1590),
.B(n_1404),
.Y(n_1662)
);

BUFx12f_ASAP7_75t_L g1663 ( 
.A(n_1445),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1492),
.B(n_719),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1443),
.B(n_1407),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1623),
.A2(n_1410),
.B(n_1406),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1449),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1598),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1537),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1450),
.A2(n_1413),
.B(n_1411),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1527),
.B(n_1415),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1613),
.A2(n_1417),
.B(n_1414),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1459),
.B(n_721),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1605),
.B(n_1499),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1544),
.B(n_722),
.Y(n_1675)
);

A2O1A1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1556),
.A2(n_1402),
.B(n_1423),
.C(n_1420),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1441),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1452),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1577),
.B(n_1430),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1590),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1613),
.A2(n_1435),
.B(n_1432),
.Y(n_1681)
);

AO22x1_ASAP7_75t_L g1682 ( 
.A1(n_1553),
.A2(n_1461),
.B1(n_1447),
.B2(n_1517),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1457),
.A2(n_1442),
.B(n_1455),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1547),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1478),
.B(n_1436),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1545),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1548),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1533),
.A2(n_780),
.B1(n_792),
.B2(n_786),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1487),
.B(n_723),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1469),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_1548),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1482),
.Y(n_1692)
);

NOR2x1_ASAP7_75t_L g1693 ( 
.A(n_1489),
.B(n_793),
.Y(n_1693)
);

OAI22x1_ASAP7_75t_L g1694 ( 
.A1(n_1580),
.A2(n_834),
.B1(n_798),
.B2(n_799),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1533),
.A2(n_801),
.B1(n_805),
.B2(n_795),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1600),
.Y(n_1696)
);

BUFx4f_ASAP7_75t_L g1697 ( 
.A(n_1445),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1442),
.A2(n_1086),
.B(n_1076),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1602),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1496),
.A2(n_1086),
.B(n_1076),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1453),
.B(n_1462),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1604),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1609),
.B(n_1076),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1456),
.A2(n_1093),
.B(n_1086),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1566),
.A2(n_725),
.B1(n_731),
.B2(n_730),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1607),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1539),
.A2(n_1093),
.B(n_1086),
.Y(n_1707)
);

INVx1_ASAP7_75t_SL g1708 ( 
.A(n_1484),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1557),
.B(n_732),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_1579),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1521),
.A2(n_733),
.B1(n_738),
.B2(n_737),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1539),
.A2(n_1590),
.B(n_1567),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1446),
.B(n_1093),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1445),
.B(n_1093),
.Y(n_1714)
);

OAI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1581),
.A2(n_1589),
.B(n_1510),
.Y(n_1715)
);

INVx3_ASAP7_75t_L g1716 ( 
.A(n_1639),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1540),
.A2(n_1093),
.B(n_1105),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1498),
.A2(n_1227),
.B(n_1062),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1490),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1540),
.A2(n_1586),
.B(n_1567),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1586),
.A2(n_1105),
.B(n_1062),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1542),
.B(n_741),
.Y(n_1722)
);

BUFx6f_ASAP7_75t_L g1723 ( 
.A(n_1579),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1551),
.A2(n_744),
.B1(n_745),
.B2(n_743),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1588),
.A2(n_1595),
.B(n_1594),
.Y(n_1725)
);

INVx3_ASAP7_75t_L g1726 ( 
.A(n_1639),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_SL g1727 ( 
.A(n_1471),
.B(n_1062),
.Y(n_1727)
);

AOI21x1_ASAP7_75t_L g1728 ( 
.A1(n_1584),
.A2(n_881),
.B(n_873),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1512),
.B(n_749),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1588),
.A2(n_1062),
.B(n_1107),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1579),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_1460),
.Y(n_1732)
);

OAI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1498),
.A2(n_1227),
.B(n_881),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1536),
.B(n_751),
.Y(n_1734)
);

BUFx2_ASAP7_75t_L g1735 ( 
.A(n_1553),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1561),
.B(n_753),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_L g1737 ( 
.A(n_1471),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_1471),
.Y(n_1738)
);

O2A1O1Ixp33_ASAP7_75t_L g1739 ( 
.A1(n_1571),
.A2(n_809),
.B(n_810),
.C(n_808),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1594),
.A2(n_1107),
.B(n_883),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1477),
.B(n_756),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1501),
.Y(n_1742)
);

NOR2xp67_ASAP7_75t_L g1743 ( 
.A(n_1500),
.B(n_515),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1519),
.B(n_757),
.Y(n_1744)
);

A2O1A1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1465),
.A2(n_827),
.B(n_828),
.C(n_815),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1520),
.B(n_1559),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1532),
.B(n_1473),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1491),
.B(n_759),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1595),
.A2(n_1601),
.B(n_1597),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1552),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1548),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1502),
.B(n_760),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1597),
.A2(n_1107),
.B(n_883),
.Y(n_1753)
);

NAND3xp33_ASAP7_75t_L g1754 ( 
.A(n_1635),
.B(n_765),
.C(n_762),
.Y(n_1754)
);

NAND2xp33_ASAP7_75t_L g1755 ( 
.A(n_1522),
.B(n_1227),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1639),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1495),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1503),
.B(n_766),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1637),
.B(n_767),
.Y(n_1759)
);

OAI21xp33_ASAP7_75t_L g1760 ( 
.A1(n_1629),
.A2(n_816),
.B(n_772),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1601),
.A2(n_1616),
.B(n_1596),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1550),
.B(n_768),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1529),
.A2(n_773),
.B1(n_774),
.B2(n_769),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1508),
.B(n_778),
.Y(n_1764)
);

AND2x2_ASAP7_75t_SL g1765 ( 
.A(n_1467),
.B(n_781),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1565),
.B(n_779),
.Y(n_1766)
);

INVx1_ASAP7_75t_SL g1767 ( 
.A(n_1552),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1485),
.B(n_782),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1608),
.B(n_1227),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1524),
.Y(n_1770)
);

AOI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1552),
.A2(n_789),
.B1(n_791),
.B2(n_788),
.Y(n_1771)
);

O2A1O1Ixp33_ASAP7_75t_L g1772 ( 
.A1(n_1543),
.A2(n_835),
.B(n_837),
.C(n_829),
.Y(n_1772)
);

OAI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1510),
.A2(n_1227),
.B(n_884),
.Y(n_1773)
);

INVx2_ASAP7_75t_SL g1774 ( 
.A(n_1636),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1608),
.B(n_1227),
.Y(n_1775)
);

BUFx12f_ASAP7_75t_L g1776 ( 
.A(n_1636),
.Y(n_1776)
);

O2A1O1Ixp33_ASAP7_75t_L g1777 ( 
.A1(n_1493),
.A2(n_842),
.B(n_887),
.C(n_882),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1578),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1518),
.B(n_941),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1546),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1619),
.A2(n_1107),
.B(n_942),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1570),
.B(n_794),
.Y(n_1782)
);

NAND2x1p5_ASAP7_75t_L g1783 ( 
.A(n_1639),
.B(n_946),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1628),
.A2(n_942),
.B(n_940),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1610),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1516),
.A2(n_943),
.B(n_940),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1516),
.A2(n_944),
.B(n_943),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1486),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1528),
.B(n_802),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1494),
.B(n_803),
.Y(n_1790)
);

AND2x2_ASAP7_75t_SL g1791 ( 
.A(n_1444),
.B(n_783),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1505),
.B(n_804),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1464),
.B(n_807),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1573),
.B(n_812),
.Y(n_1794)
);

INVx3_ASAP7_75t_L g1795 ( 
.A(n_1486),
.Y(n_1795)
);

OAI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1535),
.A2(n_781),
.B1(n_783),
.B2(n_771),
.Y(n_1796)
);

INVx11_ASAP7_75t_L g1797 ( 
.A(n_1534),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1488),
.B(n_813),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1514),
.B(n_814),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1575),
.B(n_819),
.Y(n_1800)
);

INVx1_ASAP7_75t_SL g1801 ( 
.A(n_1476),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1575),
.B(n_821),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1526),
.A2(n_949),
.B(n_946),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1525),
.B(n_822),
.Y(n_1804)
);

AOI21xp33_ASAP7_75t_L g1805 ( 
.A1(n_1624),
.A2(n_951),
.B(n_823),
.Y(n_1805)
);

BUFx3_ASAP7_75t_L g1806 ( 
.A(n_1636),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1611),
.B(n_1612),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1448),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1587),
.A2(n_797),
.B(n_781),
.Y(n_1809)
);

O2A1O1Ixp33_ASAP7_75t_L g1810 ( 
.A1(n_1549),
.A2(n_1568),
.B(n_1558),
.C(n_1572),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1615),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_SL g1812 ( 
.A(n_1522),
.B(n_724),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1535),
.A2(n_785),
.B(n_797),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1454),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1481),
.B(n_739),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1522),
.B(n_740),
.Y(n_1816)
);

AOI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1582),
.A2(n_797),
.B(n_785),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1582),
.A2(n_797),
.B(n_785),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1622),
.B(n_797),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_1522),
.Y(n_1820)
);

BUFx2_ASAP7_75t_L g1821 ( 
.A(n_1554),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1618),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_SL g1823 ( 
.A(n_1522),
.B(n_775),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1625),
.B(n_921),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1631),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1603),
.A2(n_1620),
.B(n_1614),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1632),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1674),
.B(n_1617),
.Y(n_1828)
);

AOI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1651),
.A2(n_1614),
.B(n_1603),
.Y(n_1829)
);

AOI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1643),
.A2(n_1621),
.B(n_1620),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1642),
.B(n_1463),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1765),
.A2(n_1480),
.B1(n_1472),
.B2(n_1475),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1791),
.B(n_1638),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1684),
.B(n_1466),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1662),
.B(n_1638),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1757),
.A2(n_1497),
.B1(n_1507),
.B2(n_1479),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1648),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1712),
.A2(n_1626),
.B(n_1621),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1683),
.A2(n_1627),
.B(n_1626),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1748),
.A2(n_1583),
.B1(n_1633),
.B2(n_1599),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1646),
.A2(n_1755),
.B(n_1707),
.Y(n_1841)
);

AOI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1640),
.A2(n_1725),
.B(n_1720),
.Y(n_1842)
);

A2O1A1Ixp33_ASAP7_75t_L g1843 ( 
.A1(n_1660),
.A2(n_1560),
.B(n_1630),
.C(n_1483),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1652),
.A2(n_1599),
.B1(n_1634),
.B2(n_1606),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1685),
.B(n_1509),
.Y(n_1845)
);

AND2x4_ASAP7_75t_L g1846 ( 
.A(n_1767),
.B(n_1554),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1671),
.B(n_1513),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1659),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_SL g1849 ( 
.A(n_1708),
.B(n_1563),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1749),
.A2(n_1627),
.B(n_1606),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1665),
.B(n_1515),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1650),
.B(n_3),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1826),
.A2(n_1506),
.B(n_1599),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1653),
.A2(n_1704),
.B(n_1698),
.Y(n_1854)
);

AOI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1664),
.A2(n_1655),
.B1(n_1772),
.B2(n_1658),
.C(n_1673),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1670),
.A2(n_1645),
.B(n_1662),
.Y(n_1856)
);

AO32x1_ASAP7_75t_L g1857 ( 
.A1(n_1658),
.A2(n_1562),
.A3(n_1569),
.B1(n_1564),
.B2(n_1541),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1701),
.B(n_4),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1708),
.B(n_5),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1747),
.A2(n_1574),
.B1(n_1522),
.B2(n_787),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1718),
.A2(n_784),
.B(n_955),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1746),
.Y(n_1862)
);

AOI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1718),
.A2(n_978),
.B(n_955),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_R g1864 ( 
.A(n_1732),
.B(n_516),
.Y(n_1864)
);

A2O1A1Ixp33_ASAP7_75t_L g1865 ( 
.A1(n_1810),
.A2(n_8),
.B(n_6),
.C(n_7),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1686),
.B(n_1654),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1736),
.A2(n_9),
.B1(n_6),
.B2(n_7),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1675),
.B(n_9),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1667),
.B(n_10),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1700),
.A2(n_979),
.B(n_978),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1717),
.A2(n_979),
.B(n_978),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1820),
.A2(n_979),
.B(n_978),
.Y(n_1872)
);

NOR2x1p5_ASAP7_75t_SL g1873 ( 
.A(n_1728),
.B(n_978),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1688),
.A2(n_991),
.B1(n_999),
.B2(n_979),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1657),
.B(n_979),
.Y(n_1875)
);

O2A1O1Ixp33_ASAP7_75t_L g1876 ( 
.A1(n_1729),
.A2(n_13),
.B(n_11),
.C(n_12),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1770),
.B(n_11),
.Y(n_1877)
);

OA22x2_ASAP7_75t_L g1878 ( 
.A1(n_1694),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1722),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1761),
.A2(n_999),
.B(n_991),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1815),
.A2(n_999),
.B1(n_991),
.B2(n_17),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1641),
.B(n_15),
.Y(n_1882)
);

O2A1O1Ixp33_ASAP7_75t_L g1883 ( 
.A1(n_1739),
.A2(n_19),
.B(n_16),
.C(n_17),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1800),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1703),
.A2(n_999),
.B(n_991),
.Y(n_1885)
);

AOI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1730),
.A2(n_999),
.B(n_991),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1767),
.B(n_21),
.Y(n_1887)
);

AOI21x1_ASAP7_75t_L g1888 ( 
.A1(n_1803),
.A2(n_518),
.B(n_517),
.Y(n_1888)
);

OAI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1661),
.A2(n_22),
.B(n_23),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1672),
.A2(n_22),
.B(n_24),
.Y(n_1890)
);

OAI21xp33_ASAP7_75t_L g1891 ( 
.A1(n_1711),
.A2(n_24),
.B(n_25),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1668),
.Y(n_1892)
);

BUFx6f_ASAP7_75t_L g1893 ( 
.A(n_1649),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1677),
.B(n_25),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1678),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1762),
.B(n_26),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1680),
.B(n_27),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1690),
.Y(n_1898)
);

OAI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1709),
.A2(n_27),
.B(n_28),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1692),
.B(n_28),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1719),
.B(n_29),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1742),
.B(n_30),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1680),
.B(n_30),
.Y(n_1903)
);

NAND2x1_ASAP7_75t_L g1904 ( 
.A(n_1788),
.B(n_519),
.Y(n_1904)
);

BUFx6f_ASAP7_75t_L g1905 ( 
.A(n_1691),
.Y(n_1905)
);

O2A1O1Ixp33_ASAP7_75t_L g1906 ( 
.A1(n_1802),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1681),
.A2(n_32),
.B(n_33),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1801),
.B(n_34),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1780),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_L g1910 ( 
.A(n_1766),
.B(n_34),
.Y(n_1910)
);

OAI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1798),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1785),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1721),
.A2(n_36),
.B(n_37),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1793),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1914)
);

NOR3xp33_ASAP7_75t_L g1915 ( 
.A(n_1688),
.B(n_38),
.C(n_39),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1811),
.Y(n_1916)
);

AOI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1715),
.A2(n_1816),
.B(n_1812),
.Y(n_1917)
);

NOR2x1_ASAP7_75t_L g1918 ( 
.A(n_1693),
.B(n_40),
.Y(n_1918)
);

CKINVDCx10_ASAP7_75t_R g1919 ( 
.A(n_1697),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_SL g1920 ( 
.A(n_1801),
.B(n_41),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1782),
.B(n_42),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_SL g1922 ( 
.A(n_1807),
.B(n_42),
.Y(n_1922)
);

AOI21xp5_ASAP7_75t_L g1923 ( 
.A1(n_1715),
.A2(n_43),
.B(n_45),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1823),
.A2(n_43),
.B(n_45),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1695),
.B(n_46),
.Y(n_1925)
);

INVx3_ASAP7_75t_L g1926 ( 
.A(n_1710),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1644),
.B(n_1669),
.Y(n_1927)
);

AOI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1817),
.A2(n_1818),
.B(n_1713),
.Y(n_1928)
);

INVx3_ASAP7_75t_L g1929 ( 
.A(n_1710),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1769),
.A2(n_46),
.B(n_47),
.Y(n_1930)
);

BUFx12f_ASAP7_75t_L g1931 ( 
.A(n_1663),
.Y(n_1931)
);

A2O1A1Ixp33_ASAP7_75t_L g1932 ( 
.A1(n_1760),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_1932)
);

AOI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1768),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1695),
.B(n_50),
.Y(n_1934)
);

O2A1O1Ixp33_ASAP7_75t_L g1935 ( 
.A1(n_1789),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1822),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1769),
.A2(n_54),
.B(n_55),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_SL g1938 ( 
.A(n_1788),
.B(n_54),
.Y(n_1938)
);

INVx3_ASAP7_75t_L g1939 ( 
.A(n_1710),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1687),
.B(n_1751),
.Y(n_1940)
);

A2O1A1Ixp33_ASAP7_75t_L g1941 ( 
.A1(n_1754),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1735),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1682),
.B(n_57),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1825),
.Y(n_1944)
);

INVx3_ASAP7_75t_L g1945 ( 
.A(n_1723),
.Y(n_1945)
);

AOI22xp33_ASAP7_75t_SL g1946 ( 
.A1(n_1819),
.A2(n_60),
.B1(n_61),
.B2(n_59),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_L g1947 ( 
.A1(n_1775),
.A2(n_58),
.B(n_59),
.Y(n_1947)
);

OAI22x1_ASAP7_75t_L g1948 ( 
.A1(n_1827),
.A2(n_62),
.B1(n_58),
.B2(n_61),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1775),
.A2(n_62),
.B(n_63),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1696),
.Y(n_1950)
);

AOI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1740),
.A2(n_63),
.B(n_64),
.Y(n_1951)
);

AND2x4_ASAP7_75t_L g1952 ( 
.A(n_1806),
.B(n_65),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1699),
.B(n_66),
.Y(n_1953)
);

BUFx2_ASAP7_75t_L g1954 ( 
.A(n_1723),
.Y(n_1954)
);

BUFx6f_ASAP7_75t_L g1955 ( 
.A(n_1697),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1702),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1795),
.B(n_66),
.Y(n_1957)
);

AOI21xp5_ASAP7_75t_L g1958 ( 
.A1(n_1753),
.A2(n_67),
.B(n_68),
.Y(n_1958)
);

INVx5_ASAP7_75t_L g1959 ( 
.A(n_1737),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1706),
.B(n_67),
.Y(n_1960)
);

AOI21x1_ASAP7_75t_L g1961 ( 
.A1(n_1786),
.A2(n_521),
.B(n_520),
.Y(n_1961)
);

OR2x6_ASAP7_75t_L g1962 ( 
.A(n_1679),
.B(n_604),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1774),
.B(n_68),
.Y(n_1963)
);

OAI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1705),
.A2(n_69),
.B(n_70),
.Y(n_1964)
);

NAND3xp33_ASAP7_75t_L g1965 ( 
.A(n_1799),
.B(n_69),
.C(n_70),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1737),
.B(n_71),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1795),
.B(n_71),
.Y(n_1967)
);

OAI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1676),
.A2(n_72),
.B(n_73),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1808),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1814),
.Y(n_1970)
);

OAI21x1_ASAP7_75t_L g1971 ( 
.A1(n_1813),
.A2(n_523),
.B(n_522),
.Y(n_1971)
);

AOI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1804),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1972)
);

AOI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1733),
.A2(n_74),
.B(n_76),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1821),
.B(n_1689),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1778),
.Y(n_1975)
);

HB1xp67_ASAP7_75t_L g1976 ( 
.A(n_1723),
.Y(n_1976)
);

AOI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1794),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_1977)
);

INVx3_ASAP7_75t_SL g1978 ( 
.A(n_1737),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1779),
.Y(n_1979)
);

AOI21x1_ASAP7_75t_L g1980 ( 
.A1(n_1787),
.A2(n_528),
.B(n_524),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1779),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1759),
.B(n_79),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1738),
.B(n_79),
.Y(n_1983)
);

AOI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1733),
.A2(n_80),
.B(n_81),
.Y(n_1984)
);

AOI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1773),
.A2(n_81),
.B(n_82),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1824),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1773),
.A2(n_82),
.B(n_83),
.Y(n_1987)
);

AOI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1776),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1771),
.A2(n_87),
.B1(n_84),
.B2(n_85),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1750),
.B(n_88),
.Y(n_1990)
);

NOR3xp33_ASAP7_75t_L g1991 ( 
.A(n_1734),
.B(n_88),
.C(n_89),
.Y(n_1991)
);

AOI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1656),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_1992)
);

BUFx8_ASAP7_75t_SL g1993 ( 
.A(n_1738),
.Y(n_1993)
);

OAI321xp33_ASAP7_75t_L g1994 ( 
.A1(n_1796),
.A2(n_92),
.A3(n_94),
.B1(n_90),
.B2(n_91),
.C(n_93),
.Y(n_1994)
);

AOI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1764),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1995)
);

OAI21xp33_ASAP7_75t_L g1996 ( 
.A1(n_1724),
.A2(n_96),
.B(n_97),
.Y(n_1996)
);

OAI22xp5_ASAP7_75t_L g1997 ( 
.A1(n_1763),
.A2(n_99),
.B1(n_96),
.B2(n_98),
.Y(n_1997)
);

AOI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1743),
.A2(n_1792),
.B1(n_1790),
.B2(n_1741),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1744),
.B(n_98),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1837),
.Y(n_2000)
);

OAI21xp5_ASAP7_75t_L g2001 ( 
.A1(n_1855),
.A2(n_1805),
.B(n_1809),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1955),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1862),
.B(n_1866),
.Y(n_2003)
);

INVx2_ASAP7_75t_SL g2004 ( 
.A(n_1893),
.Y(n_2004)
);

OA21x2_ASAP7_75t_L g2005 ( 
.A1(n_1842),
.A2(n_1854),
.B(n_1841),
.Y(n_2005)
);

INVx2_ASAP7_75t_SL g2006 ( 
.A(n_1893),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1828),
.B(n_1738),
.Y(n_2007)
);

AOI21xp5_ASAP7_75t_L g2008 ( 
.A1(n_1850),
.A2(n_1796),
.B(n_1714),
.Y(n_2008)
);

A2O1A1Ixp33_ASAP7_75t_L g2009 ( 
.A1(n_1868),
.A2(n_1777),
.B(n_1745),
.C(n_1805),
.Y(n_2009)
);

AOI21xp5_ASAP7_75t_L g2010 ( 
.A1(n_1829),
.A2(n_1666),
.B(n_1727),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1848),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1895),
.B(n_1731),
.Y(n_2012)
);

OAI22x1_ASAP7_75t_L g2013 ( 
.A1(n_1921),
.A2(n_1752),
.B1(n_1758),
.B2(n_1647),
.Y(n_2013)
);

INVxp67_ASAP7_75t_L g2014 ( 
.A(n_1974),
.Y(n_2014)
);

OAI21x1_ASAP7_75t_L g2015 ( 
.A1(n_1853),
.A2(n_1666),
.B(n_1784),
.Y(n_2015)
);

NAND3x1_ASAP7_75t_L g2016 ( 
.A(n_1896),
.B(n_1726),
.C(n_1716),
.Y(n_2016)
);

BUFx12f_ASAP7_75t_L g2017 ( 
.A(n_1931),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1898),
.B(n_1731),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_L g2019 ( 
.A(n_1910),
.B(n_1797),
.Y(n_2019)
);

OR2x6_ASAP7_75t_L g2020 ( 
.A(n_1962),
.B(n_1731),
.Y(n_2020)
);

NOR2x1_ASAP7_75t_SL g2021 ( 
.A(n_1962),
.B(n_1716),
.Y(n_2021)
);

AOI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_1830),
.A2(n_1781),
.B(n_1783),
.Y(n_2022)
);

OAI21x1_ASAP7_75t_L g2023 ( 
.A1(n_1928),
.A2(n_1756),
.B(n_1726),
.Y(n_2023)
);

OAI21xp5_ASAP7_75t_L g2024 ( 
.A1(n_1968),
.A2(n_99),
.B(n_100),
.Y(n_2024)
);

AO21x2_ASAP7_75t_L g2025 ( 
.A1(n_1917),
.A2(n_530),
.B(n_529),
.Y(n_2025)
);

AOI31xp67_ASAP7_75t_L g2026 ( 
.A1(n_1938),
.A2(n_102),
.A3(n_100),
.B(n_101),
.Y(n_2026)
);

AO31x2_ASAP7_75t_L g2027 ( 
.A1(n_1838),
.A2(n_532),
.A3(n_533),
.B(n_531),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1909),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1912),
.B(n_103),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1887),
.B(n_105),
.Y(n_2030)
);

OAI21xp5_ASAP7_75t_L g2031 ( 
.A1(n_1865),
.A2(n_106),
.B(n_107),
.Y(n_2031)
);

NOR2x1_ASAP7_75t_SL g2032 ( 
.A(n_1962),
.B(n_106),
.Y(n_2032)
);

AO32x2_ASAP7_75t_L g2033 ( 
.A1(n_1884),
.A2(n_109),
.A3(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1916),
.B(n_108),
.Y(n_2034)
);

OAI21xp33_ASAP7_75t_L g2035 ( 
.A1(n_1889),
.A2(n_1972),
.B(n_1933),
.Y(n_2035)
);

AO22x2_ASAP7_75t_L g2036 ( 
.A1(n_1950),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1936),
.B(n_111),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1944),
.Y(n_2038)
);

OAI22xp5_ASAP7_75t_L g2039 ( 
.A1(n_1925),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_2039)
);

OAI21x1_ASAP7_75t_L g2040 ( 
.A1(n_1839),
.A2(n_535),
.B(n_534),
.Y(n_2040)
);

NOR2xp67_ASAP7_75t_L g2041 ( 
.A(n_1965),
.B(n_1959),
.Y(n_2041)
);

A2O1A1Ixp33_ASAP7_75t_L g2042 ( 
.A1(n_1998),
.A2(n_116),
.B(n_113),
.C(n_115),
.Y(n_2042)
);

BUFx10_ASAP7_75t_L g2043 ( 
.A(n_1955),
.Y(n_2043)
);

AOI21xp5_ASAP7_75t_L g2044 ( 
.A1(n_1856),
.A2(n_115),
.B(n_116),
.Y(n_2044)
);

BUFx12f_ASAP7_75t_L g2045 ( 
.A(n_1942),
.Y(n_2045)
);

OAI22xp5_ASAP7_75t_L g2046 ( 
.A1(n_1934),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_2046)
);

AOI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_1835),
.A2(n_117),
.B(n_120),
.Y(n_2047)
);

AOI21x1_ASAP7_75t_L g2048 ( 
.A1(n_1923),
.A2(n_121),
.B(n_122),
.Y(n_2048)
);

OAI21x1_ASAP7_75t_L g2049 ( 
.A1(n_1888),
.A2(n_537),
.B(n_536),
.Y(n_2049)
);

OAI21xp5_ASAP7_75t_L g2050 ( 
.A1(n_1973),
.A2(n_121),
.B(n_122),
.Y(n_2050)
);

A2O1A1Ixp33_ASAP7_75t_L g2051 ( 
.A1(n_1891),
.A2(n_126),
.B(n_123),
.C(n_124),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1887),
.B(n_123),
.Y(n_2052)
);

OAI21x1_ASAP7_75t_L g2053 ( 
.A1(n_1961),
.A2(n_539),
.B(n_538),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1831),
.B(n_124),
.Y(n_2054)
);

A2O1A1Ixp33_ASAP7_75t_L g2055 ( 
.A1(n_1996),
.A2(n_128),
.B(n_126),
.C(n_127),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1984),
.A2(n_127),
.B(n_128),
.Y(n_2056)
);

OAI21x1_ASAP7_75t_L g2057 ( 
.A1(n_1980),
.A2(n_541),
.B(n_540),
.Y(n_2057)
);

OAI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_1985),
.A2(n_1987),
.B(n_1964),
.Y(n_2058)
);

AOI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_1915),
.A2(n_132),
.B1(n_129),
.B2(n_130),
.Y(n_2059)
);

INVx2_ASAP7_75t_SL g2060 ( 
.A(n_1893),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1834),
.Y(n_2061)
);

OAI21x1_ASAP7_75t_L g2062 ( 
.A1(n_1863),
.A2(n_543),
.B(n_542),
.Y(n_2062)
);

AO31x2_ASAP7_75t_L g2063 ( 
.A1(n_1979),
.A2(n_546),
.A3(n_547),
.B(n_545),
.Y(n_2063)
);

NAND2x1p5_ASAP7_75t_L g2064 ( 
.A(n_1959),
.B(n_548),
.Y(n_2064)
);

AO32x2_ASAP7_75t_L g2065 ( 
.A1(n_1879),
.A2(n_132),
.A3(n_129),
.B1(n_130),
.B2(n_134),
.Y(n_2065)
);

OAI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_1977),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_2066)
);

OAI21x1_ASAP7_75t_L g2067 ( 
.A1(n_1971),
.A2(n_552),
.B(n_551),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1845),
.B(n_137),
.Y(n_2068)
);

AOI22xp5_ASAP7_75t_L g2069 ( 
.A1(n_1840),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_2069)
);

OR2x6_ASAP7_75t_L g2070 ( 
.A(n_1955),
.B(n_553),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1849),
.B(n_555),
.Y(n_2071)
);

AOI221xp5_ASAP7_75t_L g2072 ( 
.A1(n_1991),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.C(n_144),
.Y(n_2072)
);

OAI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_1899),
.A2(n_141),
.B(n_142),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1986),
.B(n_143),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1981),
.Y(n_2075)
);

BUFx6f_ASAP7_75t_L g2076 ( 
.A(n_1905),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_1976),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1858),
.B(n_144),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1847),
.B(n_145),
.Y(n_2079)
);

AO31x2_ASAP7_75t_L g2080 ( 
.A1(n_1969),
.A2(n_557),
.A3(n_558),
.B(n_556),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1851),
.B(n_145),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1959),
.B(n_559),
.Y(n_2082)
);

AND2x4_ASAP7_75t_L g2083 ( 
.A(n_1846),
.B(n_560),
.Y(n_2083)
);

OAI21x1_ASAP7_75t_L g2084 ( 
.A1(n_1930),
.A2(n_564),
.B(n_562),
.Y(n_2084)
);

NOR3xp33_ASAP7_75t_L g2085 ( 
.A(n_1914),
.B(n_146),
.C(n_147),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1990),
.B(n_147),
.Y(n_2086)
);

OAI21x1_ASAP7_75t_L g2087 ( 
.A1(n_1937),
.A2(n_568),
.B(n_565),
.Y(n_2087)
);

HB1xp67_ASAP7_75t_L g2088 ( 
.A(n_1954),
.Y(n_2088)
);

O2A1O1Ixp5_ASAP7_75t_L g2089 ( 
.A1(n_1911),
.A2(n_151),
.B(n_148),
.C(n_150),
.Y(n_2089)
);

AO31x2_ASAP7_75t_L g2090 ( 
.A1(n_1970),
.A2(n_573),
.A3(n_575),
.B(n_570),
.Y(n_2090)
);

INVx3_ASAP7_75t_SL g2091 ( 
.A(n_1978),
.Y(n_2091)
);

OAI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_1932),
.A2(n_148),
.B(n_150),
.Y(n_2092)
);

INVx3_ASAP7_75t_L g2093 ( 
.A(n_1926),
.Y(n_2093)
);

INVx4_ASAP7_75t_L g2094 ( 
.A(n_1905),
.Y(n_2094)
);

OAI21x1_ASAP7_75t_L g2095 ( 
.A1(n_1947),
.A2(n_580),
.B(n_578),
.Y(n_2095)
);

OAI21x1_ASAP7_75t_L g2096 ( 
.A1(n_1949),
.A2(n_583),
.B(n_581),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1990),
.B(n_151),
.Y(n_2097)
);

OAI21x1_ASAP7_75t_L g2098 ( 
.A1(n_1880),
.A2(n_586),
.B(n_585),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1882),
.B(n_1894),
.Y(n_2099)
);

BUFx3_ASAP7_75t_L g2100 ( 
.A(n_1993),
.Y(n_2100)
);

AOI21xp5_ASAP7_75t_L g2101 ( 
.A1(n_1833),
.A2(n_152),
.B(n_153),
.Y(n_2101)
);

OAI21x1_ASAP7_75t_L g2102 ( 
.A1(n_1871),
.A2(n_592),
.B(n_589),
.Y(n_2102)
);

OAI21x1_ASAP7_75t_L g2103 ( 
.A1(n_1886),
.A2(n_594),
.B(n_593),
.Y(n_2103)
);

OAI21x1_ASAP7_75t_L g2104 ( 
.A1(n_1913),
.A2(n_596),
.B(n_595),
.Y(n_2104)
);

NOR3xp33_ASAP7_75t_L g2105 ( 
.A(n_1876),
.B(n_153),
.C(n_154),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1900),
.B(n_154),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1892),
.Y(n_2107)
);

AND2x4_ASAP7_75t_L g2108 ( 
.A(n_1846),
.B(n_598),
.Y(n_2108)
);

OAI21x1_ASAP7_75t_L g2109 ( 
.A1(n_1890),
.A2(n_600),
.B(n_599),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1956),
.Y(n_2110)
);

AOI21xp5_ASAP7_75t_L g2111 ( 
.A1(n_1844),
.A2(n_1907),
.B(n_1875),
.Y(n_2111)
);

AOI211x1_ASAP7_75t_L g2112 ( 
.A1(n_1867),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_2112)
);

OAI21x1_ASAP7_75t_L g2113 ( 
.A1(n_1870),
.A2(n_602),
.B(n_601),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1901),
.B(n_155),
.Y(n_2114)
);

OAI21xp5_ASAP7_75t_L g2115 ( 
.A1(n_1883),
.A2(n_1935),
.B(n_1906),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2038),
.Y(n_2116)
);

CKINVDCx20_ASAP7_75t_R g2117 ( 
.A(n_2100),
.Y(n_2117)
);

NOR2xp33_ASAP7_75t_L g2118 ( 
.A(n_2019),
.B(n_1905),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_2000),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2038),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2014),
.B(n_1943),
.Y(n_2121)
);

BUFx3_ASAP7_75t_L g2122 ( 
.A(n_2017),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2028),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2075),
.Y(n_2124)
);

A2O1A1Ixp33_ASAP7_75t_L g2125 ( 
.A1(n_2035),
.A2(n_1988),
.B(n_1992),
.C(n_1999),
.Y(n_2125)
);

INVx2_ASAP7_75t_SL g2126 ( 
.A(n_2076),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2003),
.B(n_1902),
.Y(n_2127)
);

INVx2_ASAP7_75t_SL g2128 ( 
.A(n_2076),
.Y(n_2128)
);

OAI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_2024),
.A2(n_1995),
.B1(n_1946),
.B2(n_1881),
.Y(n_2129)
);

NAND3xp33_ASAP7_75t_L g2130 ( 
.A(n_2105),
.B(n_1989),
.C(n_1941),
.Y(n_2130)
);

AOI21xp5_ASAP7_75t_L g2131 ( 
.A1(n_2058),
.A2(n_1994),
.B(n_1958),
.Y(n_2131)
);

BUFx6f_ASAP7_75t_L g2132 ( 
.A(n_2076),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2075),
.Y(n_2133)
);

AO22x1_ASAP7_75t_L g2134 ( 
.A1(n_2073),
.A2(n_1952),
.B1(n_1983),
.B2(n_1966),
.Y(n_2134)
);

AOI21xp5_ASAP7_75t_L g2135 ( 
.A1(n_2008),
.A2(n_1951),
.B(n_1843),
.Y(n_2135)
);

BUFx6f_ASAP7_75t_L g2136 ( 
.A(n_2002),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2088),
.B(n_2077),
.Y(n_2137)
);

BUFx6f_ASAP7_75t_L g2138 ( 
.A(n_2002),
.Y(n_2138)
);

OR2x2_ASAP7_75t_L g2139 ( 
.A(n_2061),
.B(n_2018),
.Y(n_2139)
);

OAI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_2069),
.A2(n_1878),
.B1(n_1997),
.B2(n_1920),
.Y(n_2140)
);

OAI22xp5_ASAP7_75t_L g2141 ( 
.A1(n_2059),
.A2(n_2042),
.B1(n_2036),
.B2(n_2055),
.Y(n_2141)
);

AOI22xp33_ASAP7_75t_L g2142 ( 
.A1(n_2092),
.A2(n_1982),
.B1(n_1852),
.B2(n_1836),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2007),
.B(n_2099),
.Y(n_2143)
);

OAI21x1_ASAP7_75t_L g2144 ( 
.A1(n_2015),
.A2(n_1904),
.B(n_1885),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2012),
.B(n_1869),
.Y(n_2145)
);

AND2x4_ASAP7_75t_L g2146 ( 
.A(n_2021),
.B(n_1952),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_L g2147 ( 
.A(n_2091),
.B(n_1919),
.Y(n_2147)
);

AOI22xp5_ASAP7_75t_L g2148 ( 
.A1(n_2085),
.A2(n_1948),
.B1(n_1918),
.B2(n_1908),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2107),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2054),
.B(n_1877),
.Y(n_2150)
);

INVx3_ASAP7_75t_L g2151 ( 
.A(n_2093),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_2041),
.B(n_1864),
.Y(n_2152)
);

INVxp67_ASAP7_75t_L g2153 ( 
.A(n_2004),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2068),
.B(n_1859),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2110),
.Y(n_2155)
);

NOR2xp33_ASAP7_75t_L g2156 ( 
.A(n_2045),
.B(n_2094),
.Y(n_2156)
);

AOI21x1_ASAP7_75t_L g2157 ( 
.A1(n_2013),
.A2(n_2034),
.B(n_2029),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2011),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2037),
.Y(n_2159)
);

A2O1A1Ixp33_ASAP7_75t_SL g2160 ( 
.A1(n_2050),
.A2(n_1927),
.B(n_1940),
.C(n_1924),
.Y(n_2160)
);

HAxp5_ASAP7_75t_L g2161 ( 
.A(n_2072),
.B(n_156),
.CON(n_2161),
.SN(n_2161)
);

AOI21xp5_ASAP7_75t_L g2162 ( 
.A1(n_2020),
.A2(n_1861),
.B(n_1874),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2036),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2074),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2093),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_2081),
.Y(n_2166)
);

BUFx2_ASAP7_75t_L g2167 ( 
.A(n_2094),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2079),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2021),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2030),
.B(n_1953),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_2063),
.Y(n_2171)
);

AOI22xp33_ASAP7_75t_SL g2172 ( 
.A1(n_2032),
.A2(n_1975),
.B1(n_1960),
.B2(n_1963),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_2063),
.Y(n_2173)
);

AND2x4_ASAP7_75t_L g2174 ( 
.A(n_2020),
.B(n_2006),
.Y(n_2174)
);

OAI22xp5_ASAP7_75t_L g2175 ( 
.A1(n_2051),
.A2(n_1860),
.B1(n_1922),
.B2(n_1874),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2033),
.Y(n_2176)
);

BUFx2_ASAP7_75t_R g2177 ( 
.A(n_2086),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_2097),
.B(n_1926),
.Y(n_2178)
);

AND2x4_ASAP7_75t_L g2179 ( 
.A(n_2060),
.B(n_1929),
.Y(n_2179)
);

NOR2xp33_ASAP7_75t_L g2180 ( 
.A(n_2078),
.B(n_1919),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2033),
.Y(n_2181)
);

O2A1O1Ixp33_ASAP7_75t_L g2182 ( 
.A1(n_2009),
.A2(n_1967),
.B(n_1957),
.C(n_1897),
.Y(n_2182)
);

INVx1_ASAP7_75t_SL g2183 ( 
.A(n_2016),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2033),
.Y(n_2184)
);

AOI21xp5_ASAP7_75t_L g2185 ( 
.A1(n_2005),
.A2(n_1872),
.B(n_1903),
.Y(n_2185)
);

HB1xp67_ASAP7_75t_L g2186 ( 
.A(n_2005),
.Y(n_2186)
);

BUFx12f_ASAP7_75t_L g2187 ( 
.A(n_2043),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2065),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2065),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2065),
.Y(n_2190)
);

AOI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_2066),
.A2(n_1832),
.B1(n_1939),
.B2(n_1929),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2052),
.B(n_2032),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2106),
.B(n_1939),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2143),
.B(n_2010),
.Y(n_2194)
);

BUFx2_ASAP7_75t_L g2195 ( 
.A(n_2167),
.Y(n_2195)
);

CKINVDCx11_ASAP7_75t_R g2196 ( 
.A(n_2117),
.Y(n_2196)
);

BUFx2_ASAP7_75t_L g2197 ( 
.A(n_2137),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2116),
.Y(n_2198)
);

BUFx6f_ASAP7_75t_L g2199 ( 
.A(n_2132),
.Y(n_2199)
);

INVx6_ASAP7_75t_L g2200 ( 
.A(n_2187),
.Y(n_2200)
);

CKINVDCx11_ASAP7_75t_R g2201 ( 
.A(n_2122),
.Y(n_2201)
);

CKINVDCx11_ASAP7_75t_R g2202 ( 
.A(n_2166),
.Y(n_2202)
);

INVx6_ASAP7_75t_L g2203 ( 
.A(n_2146),
.Y(n_2203)
);

OAI21xp5_ASAP7_75t_SL g2204 ( 
.A1(n_2130),
.A2(n_2115),
.B(n_2031),
.Y(n_2204)
);

INVx6_ASAP7_75t_L g2205 ( 
.A(n_2146),
.Y(n_2205)
);

CKINVDCx20_ASAP7_75t_R g2206 ( 
.A(n_2147),
.Y(n_2206)
);

AOI22xp33_ASAP7_75t_L g2207 ( 
.A1(n_2141),
.A2(n_2001),
.B1(n_2046),
.B2(n_2039),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2120),
.Y(n_2208)
);

BUFx12f_ASAP7_75t_L g2209 ( 
.A(n_2132),
.Y(n_2209)
);

INVx6_ASAP7_75t_L g2210 ( 
.A(n_2132),
.Y(n_2210)
);

BUFx10_ASAP7_75t_L g2211 ( 
.A(n_2156),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2124),
.Y(n_2212)
);

OAI22xp5_ASAP7_75t_L g2213 ( 
.A1(n_2141),
.A2(n_2112),
.B1(n_2056),
.B2(n_2044),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2133),
.Y(n_2214)
);

AOI22xp33_ASAP7_75t_L g2215 ( 
.A1(n_2129),
.A2(n_2114),
.B1(n_2101),
.B2(n_2047),
.Y(n_2215)
);

AOI22xp33_ASAP7_75t_L g2216 ( 
.A1(n_2129),
.A2(n_2070),
.B1(n_2025),
.B2(n_2111),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2127),
.B(n_2023),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2119),
.Y(n_2218)
);

NAND2x1p5_ASAP7_75t_L g2219 ( 
.A(n_2152),
.B(n_2083),
.Y(n_2219)
);

AOI22xp33_ASAP7_75t_L g2220 ( 
.A1(n_2140),
.A2(n_2070),
.B1(n_2108),
.B2(n_2083),
.Y(n_2220)
);

OAI22xp5_ASAP7_75t_L g2221 ( 
.A1(n_2148),
.A2(n_2048),
.B1(n_2071),
.B2(n_2108),
.Y(n_2221)
);

INVxp67_ASAP7_75t_SL g2222 ( 
.A(n_2186),
.Y(n_2222)
);

BUFx4f_ASAP7_75t_L g2223 ( 
.A(n_2136),
.Y(n_2223)
);

BUFx2_ASAP7_75t_L g2224 ( 
.A(n_2153),
.Y(n_2224)
);

BUFx4f_ASAP7_75t_SL g2225 ( 
.A(n_2145),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2123),
.Y(n_2226)
);

AOI22xp33_ASAP7_75t_L g2227 ( 
.A1(n_2140),
.A2(n_2109),
.B1(n_2084),
.B2(n_2095),
.Y(n_2227)
);

INVx3_ASAP7_75t_L g2228 ( 
.A(n_2151),
.Y(n_2228)
);

AOI22xp33_ASAP7_75t_L g2229 ( 
.A1(n_2163),
.A2(n_2087),
.B1(n_2096),
.B2(n_2104),
.Y(n_2229)
);

BUFx3_ASAP7_75t_L g2230 ( 
.A(n_2174),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_2158),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2192),
.B(n_2002),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2149),
.Y(n_2233)
);

INVx8_ASAP7_75t_L g2234 ( 
.A(n_2179),
.Y(n_2234)
);

BUFx8_ASAP7_75t_SL g2235 ( 
.A(n_2170),
.Y(n_2235)
);

AOI22xp33_ASAP7_75t_L g2236 ( 
.A1(n_2130),
.A2(n_2082),
.B1(n_2053),
.B2(n_2057),
.Y(n_2236)
);

BUFx3_ASAP7_75t_L g2237 ( 
.A(n_2174),
.Y(n_2237)
);

OAI22xp33_ASAP7_75t_SL g2238 ( 
.A1(n_2176),
.A2(n_2064),
.B1(n_1945),
.B2(n_1857),
.Y(n_2238)
);

CKINVDCx11_ASAP7_75t_R g2239 ( 
.A(n_2136),
.Y(n_2239)
);

AOI22xp33_ASAP7_75t_L g2240 ( 
.A1(n_2181),
.A2(n_2184),
.B1(n_2189),
.B2(n_2188),
.Y(n_2240)
);

AOI22xp33_ASAP7_75t_SL g2241 ( 
.A1(n_2190),
.A2(n_2040),
.B1(n_2049),
.B2(n_2062),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2155),
.Y(n_2242)
);

OAI22xp5_ASAP7_75t_L g2243 ( 
.A1(n_2207),
.A2(n_2125),
.B1(n_2148),
.B2(n_2172),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2218),
.Y(n_2244)
);

HB1xp67_ASAP7_75t_SL g2245 ( 
.A(n_2230),
.Y(n_2245)
);

INVx2_ASAP7_75t_SL g2246 ( 
.A(n_2203),
.Y(n_2246)
);

OAI22xp5_ASAP7_75t_L g2247 ( 
.A1(n_2207),
.A2(n_2131),
.B1(n_2183),
.B2(n_2135),
.Y(n_2247)
);

O2A1O1Ixp5_ASAP7_75t_L g2248 ( 
.A1(n_2194),
.A2(n_2134),
.B(n_2157),
.C(n_2159),
.Y(n_2248)
);

OA21x2_ASAP7_75t_L g2249 ( 
.A1(n_2222),
.A2(n_2185),
.B(n_2173),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2197),
.B(n_2169),
.Y(n_2250)
);

OAI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_2220),
.A2(n_2183),
.B1(n_2142),
.B2(n_2191),
.Y(n_2251)
);

A2O1A1Ixp33_ASAP7_75t_L g2252 ( 
.A1(n_2204),
.A2(n_2182),
.B(n_2150),
.C(n_2089),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2198),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2208),
.Y(n_2254)
);

AOI21xp5_ASAP7_75t_SL g2255 ( 
.A1(n_2221),
.A2(n_2162),
.B(n_2175),
.Y(n_2255)
);

O2A1O1Ixp33_ASAP7_75t_L g2256 ( 
.A1(n_2213),
.A2(n_2161),
.B(n_2160),
.C(n_2175),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2217),
.B(n_2164),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2195),
.B(n_2165),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2224),
.B(n_2151),
.Y(n_2259)
);

OAI22xp5_ASAP7_75t_L g2260 ( 
.A1(n_2220),
.A2(n_2191),
.B1(n_2177),
.B2(n_2178),
.Y(n_2260)
);

AOI21x1_ASAP7_75t_SL g2261 ( 
.A1(n_2232),
.A2(n_2193),
.B(n_2121),
.Y(n_2261)
);

O2A1O1Ixp33_ASAP7_75t_L g2262 ( 
.A1(n_2216),
.A2(n_2168),
.B(n_2154),
.C(n_2180),
.Y(n_2262)
);

OAI22xp5_ASAP7_75t_L g2263 ( 
.A1(n_2216),
.A2(n_2126),
.B1(n_2128),
.B2(n_2179),
.Y(n_2263)
);

AOI21xp5_ASAP7_75t_L g2264 ( 
.A1(n_2227),
.A2(n_2238),
.B(n_2236),
.Y(n_2264)
);

OA21x2_ASAP7_75t_L g2265 ( 
.A1(n_2240),
.A2(n_2171),
.B(n_2144),
.Y(n_2265)
);

O2A1O1Ixp33_ASAP7_75t_L g2266 ( 
.A1(n_2215),
.A2(n_2227),
.B(n_2219),
.C(n_2236),
.Y(n_2266)
);

HB1xp67_ASAP7_75t_L g2267 ( 
.A(n_2226),
.Y(n_2267)
);

NOR2xp67_ASAP7_75t_L g2268 ( 
.A(n_2228),
.B(n_2118),
.Y(n_2268)
);

AO21x2_ASAP7_75t_L g2269 ( 
.A1(n_2264),
.A2(n_2022),
.B(n_2233),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2257),
.B(n_2242),
.Y(n_2270)
);

INVx5_ASAP7_75t_SL g2271 ( 
.A(n_2255),
.Y(n_2271)
);

CKINVDCx5p33_ASAP7_75t_R g2272 ( 
.A(n_2245),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2250),
.B(n_2240),
.Y(n_2273)
);

BUFx2_ASAP7_75t_L g2274 ( 
.A(n_2246),
.Y(n_2274)
);

AOI22xp33_ASAP7_75t_L g2275 ( 
.A1(n_2243),
.A2(n_2215),
.B1(n_2202),
.B2(n_2225),
.Y(n_2275)
);

CKINVDCx5p33_ASAP7_75t_R g2276 ( 
.A(n_2247),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2250),
.B(n_2228),
.Y(n_2277)
);

NOR2xp33_ASAP7_75t_L g2278 ( 
.A(n_2252),
.B(n_2235),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2258),
.B(n_2203),
.Y(n_2279)
);

NOR2xp33_ASAP7_75t_R g2280 ( 
.A(n_2246),
.B(n_2196),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2270),
.Y(n_2281)
);

HB1xp67_ASAP7_75t_L g2282 ( 
.A(n_2269),
.Y(n_2282)
);

BUFx2_ASAP7_75t_L g2283 ( 
.A(n_2280),
.Y(n_2283)
);

INVx3_ASAP7_75t_L g2284 ( 
.A(n_2271),
.Y(n_2284)
);

INVx3_ASAP7_75t_L g2285 ( 
.A(n_2271),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2269),
.B(n_2259),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2270),
.B(n_2267),
.Y(n_2287)
);

OA21x2_ASAP7_75t_L g2288 ( 
.A1(n_2274),
.A2(n_2248),
.B(n_2244),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2283),
.B(n_2274),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2283),
.B(n_2286),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2287),
.Y(n_2291)
);

OAI22xp5_ASAP7_75t_L g2292 ( 
.A1(n_2283),
.A2(n_2271),
.B1(n_2276),
.B2(n_2255),
.Y(n_2292)
);

AND2x4_ASAP7_75t_L g2293 ( 
.A(n_2284),
.B(n_2269),
.Y(n_2293)
);

AOI22xp33_ASAP7_75t_L g2294 ( 
.A1(n_2282),
.A2(n_2269),
.B1(n_2271),
.B2(n_2273),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2287),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_2286),
.B(n_2271),
.Y(n_2296)
);

AND2x4_ASAP7_75t_L g2297 ( 
.A(n_2284),
.B(n_2273),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2282),
.Y(n_2298)
);

INVx3_ASAP7_75t_L g2299 ( 
.A(n_2297),
.Y(n_2299)
);

INVxp67_ASAP7_75t_SL g2300 ( 
.A(n_2289),
.Y(n_2300)
);

OR2x2_ASAP7_75t_L g2301 ( 
.A(n_2291),
.B(n_2281),
.Y(n_2301)
);

OR2x2_ASAP7_75t_L g2302 ( 
.A(n_2291),
.B(n_2281),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2298),
.Y(n_2303)
);

NAND4xp25_ASAP7_75t_L g2304 ( 
.A(n_2290),
.B(n_2289),
.C(n_2256),
.D(n_2296),
.Y(n_2304)
);

INVx3_ASAP7_75t_L g2305 ( 
.A(n_2297),
.Y(n_2305)
);

HB1xp67_ASAP7_75t_L g2306 ( 
.A(n_2297),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2297),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2290),
.B(n_2295),
.Y(n_2308)
);

OAI33xp33_ASAP7_75t_L g2309 ( 
.A1(n_2295),
.A2(n_2262),
.A3(n_2272),
.B1(n_2251),
.B2(n_2266),
.B3(n_2260),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2296),
.B(n_2271),
.Y(n_2310)
);

OR2x2_ASAP7_75t_L g2311 ( 
.A(n_2300),
.B(n_2292),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_2299),
.B(n_2280),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2306),
.Y(n_2313)
);

INVxp67_ASAP7_75t_SL g2314 ( 
.A(n_2299),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2308),
.B(n_2298),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2305),
.B(n_2278),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2305),
.B(n_2273),
.Y(n_2317)
);

NOR2xp33_ASAP7_75t_L g2318 ( 
.A(n_2304),
.B(n_2196),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2307),
.B(n_2294),
.Y(n_2319)
);

INVxp67_ASAP7_75t_L g2320 ( 
.A(n_2318),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_2312),
.B(n_2278),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2314),
.B(n_2304),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2316),
.B(n_2310),
.Y(n_2323)
);

AND2x2_ASAP7_75t_L g2324 ( 
.A(n_2321),
.B(n_2311),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2323),
.B(n_2317),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2320),
.Y(n_2326)
);

AOI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_2322),
.A2(n_2309),
.B(n_2315),
.Y(n_2327)
);

NAND4xp75_ASAP7_75t_SL g2328 ( 
.A(n_2324),
.B(n_2286),
.C(n_2288),
.D(n_2285),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2325),
.B(n_2313),
.Y(n_2329)
);

OAI21xp5_ASAP7_75t_L g2330 ( 
.A1(n_2327),
.A2(n_2315),
.B(n_2319),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2326),
.Y(n_2331)
);

AOI22xp33_ASAP7_75t_L g2332 ( 
.A1(n_2327),
.A2(n_2293),
.B1(n_2303),
.B2(n_2288),
.Y(n_2332)
);

AOI322xp5_ASAP7_75t_L g2333 ( 
.A1(n_2324),
.A2(n_2293),
.A3(n_2275),
.B1(n_2285),
.B2(n_2284),
.C1(n_2288),
.C2(n_2301),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2332),
.B(n_2302),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2331),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2329),
.Y(n_2336)
);

CKINVDCx16_ASAP7_75t_R g2337 ( 
.A(n_2330),
.Y(n_2337)
);

HB1xp67_ASAP7_75t_L g2338 ( 
.A(n_2328),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2333),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2331),
.Y(n_2340)
);

NOR2xp33_ASAP7_75t_L g2341 ( 
.A(n_2329),
.B(n_2201),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2332),
.B(n_2293),
.Y(n_2342)
);

INVx1_ASAP7_75t_SL g2343 ( 
.A(n_2329),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2337),
.B(n_2343),
.Y(n_2344)
);

OAI22xp5_ASAP7_75t_L g2345 ( 
.A1(n_2343),
.A2(n_2293),
.B1(n_2285),
.B2(n_2284),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2336),
.Y(n_2346)
);

OAI21xp5_ASAP7_75t_SL g2347 ( 
.A1(n_2341),
.A2(n_2338),
.B(n_2339),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2335),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2340),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2334),
.B(n_2288),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2342),
.Y(n_2351)
);

OAI21xp33_ASAP7_75t_L g2352 ( 
.A1(n_2341),
.A2(n_2285),
.B(n_2284),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2337),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2337),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2337),
.Y(n_2355)
);

OAI22xp33_ASAP7_75t_L g2356 ( 
.A1(n_2337),
.A2(n_2285),
.B1(n_2288),
.B2(n_2200),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2353),
.B(n_2275),
.Y(n_2357)
);

AOI22xp33_ASAP7_75t_SL g2358 ( 
.A1(n_2350),
.A2(n_2200),
.B1(n_2206),
.B2(n_2211),
.Y(n_2358)
);

OAI211xp5_ASAP7_75t_L g2359 ( 
.A1(n_2347),
.A2(n_2239),
.B(n_2200),
.C(n_2277),
.Y(n_2359)
);

AOI21xp5_ASAP7_75t_L g2360 ( 
.A1(n_2344),
.A2(n_2279),
.B(n_2277),
.Y(n_2360)
);

HB1xp67_ASAP7_75t_L g2361 ( 
.A(n_2354),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2355),
.Y(n_2362)
);

OAI22xp5_ASAP7_75t_L g2363 ( 
.A1(n_2349),
.A2(n_2279),
.B1(n_2277),
.B2(n_2254),
.Y(n_2363)
);

INVxp67_ASAP7_75t_L g2364 ( 
.A(n_2348),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_L g2365 ( 
.A(n_2346),
.B(n_2211),
.Y(n_2365)
);

AOI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2347),
.A2(n_2279),
.B(n_2259),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2352),
.B(n_2258),
.Y(n_2367)
);

OAI22xp33_ASAP7_75t_L g2368 ( 
.A1(n_2351),
.A2(n_2219),
.B1(n_2268),
.B2(n_2263),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2345),
.B(n_2253),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_2356),
.B(n_2253),
.Y(n_2370)
);

OAI211xp5_ASAP7_75t_SL g2371 ( 
.A1(n_2347),
.A2(n_2239),
.B(n_159),
.C(n_157),
.Y(n_2371)
);

OR2x2_ASAP7_75t_L g2372 ( 
.A(n_2361),
.B(n_2254),
.Y(n_2372)
);

OAI22xp5_ASAP7_75t_L g2373 ( 
.A1(n_2362),
.A2(n_2229),
.B1(n_2241),
.B2(n_2210),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2364),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_2358),
.B(n_2199),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2366),
.B(n_2249),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2371),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2357),
.Y(n_2378)
);

NOR2xp33_ASAP7_75t_L g2379 ( 
.A(n_2359),
.B(n_158),
.Y(n_2379)
);

NOR2x1p5_ASAP7_75t_L g2380 ( 
.A(n_2369),
.B(n_2209),
.Y(n_2380)
);

INVx1_ASAP7_75t_SL g2381 ( 
.A(n_2365),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2367),
.B(n_2203),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2360),
.B(n_2249),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2370),
.B(n_2249),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2363),
.Y(n_2385)
);

NOR3xp33_ASAP7_75t_L g2386 ( 
.A(n_2374),
.B(n_2368),
.C(n_2067),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_L g2387 ( 
.A(n_2377),
.B(n_2378),
.Y(n_2387)
);

NOR3xp33_ASAP7_75t_L g2388 ( 
.A(n_2381),
.B(n_159),
.C(n_160),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2372),
.B(n_2249),
.Y(n_2389)
);

XOR2xp5_ASAP7_75t_L g2390 ( 
.A(n_2385),
.B(n_160),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_SL g2391 ( 
.A(n_2379),
.B(n_2043),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2383),
.Y(n_2392)
);

NAND3xp33_ASAP7_75t_SL g2393 ( 
.A(n_2375),
.B(n_2229),
.C(n_161),
.Y(n_2393)
);

NAND3xp33_ASAP7_75t_SL g2394 ( 
.A(n_2376),
.B(n_2384),
.C(n_2382),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2380),
.B(n_2205),
.Y(n_2395)
);

NAND2x1_ASAP7_75t_L g2396 ( 
.A(n_2373),
.B(n_2205),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_SL g2397 ( 
.A(n_2377),
.B(n_2199),
.Y(n_2397)
);

A2O1A1Ixp33_ASAP7_75t_SL g2398 ( 
.A1(n_2374),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_2398)
);

NAND4xp25_ASAP7_75t_L g2399 ( 
.A(n_2377),
.B(n_164),
.C(n_162),
.D(n_163),
.Y(n_2399)
);

AOI322xp5_ASAP7_75t_L g2400 ( 
.A1(n_2377),
.A2(n_2244),
.A3(n_2026),
.B1(n_2261),
.B2(n_2214),
.C1(n_2212),
.C2(n_2265),
.Y(n_2400)
);

OAI22xp5_ASAP7_75t_L g2401 ( 
.A1(n_2372),
.A2(n_2210),
.B1(n_2205),
.B2(n_2223),
.Y(n_2401)
);

BUFx3_ASAP7_75t_L g2402 ( 
.A(n_2374),
.Y(n_2402)
);

AOI221xp5_ASAP7_75t_L g2403 ( 
.A1(n_2374),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.C(n_167),
.Y(n_2403)
);

AOI22xp5_ASAP7_75t_L g2404 ( 
.A1(n_2377),
.A2(n_2209),
.B1(n_2265),
.B2(n_2210),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_2382),
.B(n_2230),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2378),
.B(n_2265),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2378),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2402),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2390),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_L g2410 ( 
.A(n_2407),
.B(n_2399),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2387),
.Y(n_2411)
);

AOI21xp33_ASAP7_75t_L g2412 ( 
.A1(n_2392),
.A2(n_168),
.B(n_169),
.Y(n_2412)
);

NOR2x1_ASAP7_75t_L g2413 ( 
.A(n_2394),
.B(n_168),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2406),
.Y(n_2414)
);

NOR2xp33_ASAP7_75t_L g2415 ( 
.A(n_2393),
.B(n_2397),
.Y(n_2415)
);

INVxp67_ASAP7_75t_L g2416 ( 
.A(n_2388),
.Y(n_2416)
);

NAND3xp33_ASAP7_75t_L g2417 ( 
.A(n_2398),
.B(n_169),
.C(n_170),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2405),
.B(n_170),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2403),
.B(n_171),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2391),
.B(n_172),
.Y(n_2420)
);

NAND4xp25_ASAP7_75t_L g2421 ( 
.A(n_2395),
.B(n_174),
.C(n_172),
.D(n_173),
.Y(n_2421)
);

OR2x2_ASAP7_75t_L g2422 ( 
.A(n_2389),
.B(n_173),
.Y(n_2422)
);

NAND3xp33_ASAP7_75t_L g2423 ( 
.A(n_2386),
.B(n_174),
.C(n_175),
.Y(n_2423)
);

INVx2_ASAP7_75t_SL g2424 ( 
.A(n_2396),
.Y(n_2424)
);

OAI22xp5_ASAP7_75t_L g2425 ( 
.A1(n_2404),
.A2(n_2223),
.B1(n_2199),
.B2(n_2136),
.Y(n_2425)
);

NOR3x1_ASAP7_75t_L g2426 ( 
.A(n_2401),
.B(n_175),
.C(n_176),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2400),
.B(n_176),
.Y(n_2427)
);

AND3x1_ASAP7_75t_L g2428 ( 
.A(n_2388),
.B(n_177),
.C(n_178),
.Y(n_2428)
);

OAI21xp33_ASAP7_75t_L g2429 ( 
.A1(n_2402),
.A2(n_2237),
.B(n_2199),
.Y(n_2429)
);

INVx1_ASAP7_75t_SL g2430 ( 
.A(n_2402),
.Y(n_2430)
);

NAND3xp33_ASAP7_75t_SL g2431 ( 
.A(n_2407),
.B(n_178),
.C(n_179),
.Y(n_2431)
);

AND2x2_ASAP7_75t_L g2432 ( 
.A(n_2402),
.B(n_2237),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2398),
.B(n_179),
.Y(n_2433)
);

O2A1O1Ixp33_ASAP7_75t_L g2434 ( 
.A1(n_2407),
.A2(n_182),
.B(n_180),
.C(n_181),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2402),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2398),
.B(n_180),
.Y(n_2436)
);

OAI211xp5_ASAP7_75t_L g2437 ( 
.A1(n_2402),
.A2(n_184),
.B(n_182),
.C(n_183),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2402),
.Y(n_2438)
);

AND2x2_ASAP7_75t_L g2439 ( 
.A(n_2402),
.B(n_2234),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2402),
.Y(n_2440)
);

NAND4xp25_ASAP7_75t_L g2441 ( 
.A(n_2387),
.B(n_185),
.C(n_183),
.D(n_184),
.Y(n_2441)
);

AND3x1_ASAP7_75t_L g2442 ( 
.A(n_2407),
.B(n_185),
.C(n_186),
.Y(n_2442)
);

AOI311xp33_ASAP7_75t_L g2443 ( 
.A1(n_2407),
.A2(n_189),
.A3(n_186),
.B(n_187),
.C(n_190),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2398),
.B(n_187),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2442),
.Y(n_2445)
);

NAND2x1_ASAP7_75t_SL g2446 ( 
.A(n_2408),
.B(n_189),
.Y(n_2446)
);

NAND3xp33_ASAP7_75t_SL g2447 ( 
.A(n_2430),
.B(n_191),
.C(n_192),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2442),
.Y(n_2448)
);

OAI211xp5_ASAP7_75t_L g2449 ( 
.A1(n_2435),
.A2(n_194),
.B(n_191),
.C(n_193),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2413),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2424),
.B(n_2027),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2438),
.B(n_2027),
.Y(n_2452)
);

NOR3xp33_ASAP7_75t_SL g2453 ( 
.A(n_2410),
.B(n_193),
.C(n_194),
.Y(n_2453)
);

NOR4xp25_ASAP7_75t_L g2454 ( 
.A(n_2440),
.B(n_2414),
.C(n_2409),
.D(n_2411),
.Y(n_2454)
);

AOI211xp5_ASAP7_75t_L g2455 ( 
.A1(n_2415),
.A2(n_197),
.B(n_195),
.C(n_196),
.Y(n_2455)
);

NAND2x1p5_ASAP7_75t_L g2456 ( 
.A(n_2426),
.B(n_2138),
.Y(n_2456)
);

NOR3xp33_ASAP7_75t_L g2457 ( 
.A(n_2412),
.B(n_195),
.C(n_196),
.Y(n_2457)
);

AOI221xp5_ASAP7_75t_L g2458 ( 
.A1(n_2423),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.C(n_200),
.Y(n_2458)
);

OAI321xp33_ASAP7_75t_L g2459 ( 
.A1(n_2427),
.A2(n_2139),
.A3(n_2138),
.B1(n_200),
.B2(n_202),
.C(n_198),
.Y(n_2459)
);

NAND3xp33_ASAP7_75t_L g2460 ( 
.A(n_2433),
.B(n_199),
.C(n_201),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2436),
.B(n_2027),
.Y(n_2461)
);

NAND3xp33_ASAP7_75t_L g2462 ( 
.A(n_2444),
.B(n_201),
.C(n_202),
.Y(n_2462)
);

AOI221x1_ASAP7_75t_L g2463 ( 
.A1(n_2420),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.C(n_206),
.Y(n_2463)
);

AOI211xp5_ASAP7_75t_L g2464 ( 
.A1(n_2431),
.A2(n_207),
.B(n_204),
.C(n_206),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2428),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2432),
.B(n_2234),
.Y(n_2466)
);

AOI22xp5_ASAP7_75t_L g2467 ( 
.A1(n_2416),
.A2(n_2417),
.B1(n_2418),
.B2(n_2439),
.Y(n_2467)
);

AOI211xp5_ASAP7_75t_L g2468 ( 
.A1(n_2437),
.A2(n_2434),
.B(n_2421),
.C(n_2422),
.Y(n_2468)
);

AOI22xp5_ASAP7_75t_L g2469 ( 
.A1(n_2419),
.A2(n_2138),
.B1(n_2234),
.B2(n_1945),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2429),
.B(n_2441),
.Y(n_2470)
);

OAI322xp33_ASAP7_75t_L g2471 ( 
.A1(n_2425),
.A2(n_207),
.A3(n_208),
.B1(n_209),
.B2(n_210),
.C1(n_211),
.C2(n_212),
.Y(n_2471)
);

NAND5xp2_ASAP7_75t_L g2472 ( 
.A(n_2443),
.B(n_210),
.C(n_208),
.D(n_209),
.E(n_213),
.Y(n_2472)
);

NAND4xp25_ASAP7_75t_L g2473 ( 
.A(n_2430),
.B(n_215),
.C(n_213),
.D(n_214),
.Y(n_2473)
);

INVx2_ASAP7_75t_SL g2474 ( 
.A(n_2432),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2442),
.Y(n_2475)
);

NAND4xp25_ASAP7_75t_L g2476 ( 
.A(n_2430),
.B(n_216),
.C(n_214),
.D(n_215),
.Y(n_2476)
);

OAI21xp33_ASAP7_75t_L g2477 ( 
.A1(n_2430),
.A2(n_1873),
.B(n_2102),
.Y(n_2477)
);

AOI21x1_ASAP7_75t_L g2478 ( 
.A1(n_2408),
.A2(n_216),
.B(n_217),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_SL g2479 ( 
.A(n_2430),
.B(n_217),
.Y(n_2479)
);

AOI211xp5_ASAP7_75t_L g2480 ( 
.A1(n_2430),
.A2(n_220),
.B(n_218),
.C(n_219),
.Y(n_2480)
);

AND4x1_ASAP7_75t_L g2481 ( 
.A(n_2408),
.B(n_221),
.C(n_219),
.D(n_220),
.Y(n_2481)
);

NAND4xp25_ASAP7_75t_SL g2482 ( 
.A(n_2464),
.B(n_2470),
.C(n_2458),
.D(n_2468),
.Y(n_2482)
);

NAND4xp25_ASAP7_75t_L g2483 ( 
.A(n_2472),
.B(n_223),
.C(n_221),
.D(n_222),
.Y(n_2483)
);

AOI211x1_ASAP7_75t_L g2484 ( 
.A1(n_2460),
.A2(n_225),
.B(n_223),
.C(n_224),
.Y(n_2484)
);

OAI211xp5_ASAP7_75t_L g2485 ( 
.A1(n_2454),
.A2(n_227),
.B(n_225),
.C(n_226),
.Y(n_2485)
);

NAND3xp33_ASAP7_75t_SL g2486 ( 
.A(n_2450),
.B(n_226),
.C(n_227),
.Y(n_2486)
);

XNOR2xp5_ASAP7_75t_L g2487 ( 
.A(n_2481),
.B(n_228),
.Y(n_2487)
);

NOR4xp25_ASAP7_75t_L g2488 ( 
.A(n_2445),
.B(n_231),
.C(n_229),
.D(n_230),
.Y(n_2488)
);

NOR2x1_ASAP7_75t_L g2489 ( 
.A(n_2473),
.B(n_229),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2466),
.B(n_232),
.Y(n_2490)
);

NOR2x1_ASAP7_75t_L g2491 ( 
.A(n_2476),
.B(n_232),
.Y(n_2491)
);

NAND4xp75_ASAP7_75t_L g2492 ( 
.A(n_2448),
.B(n_2475),
.C(n_2474),
.D(n_2467),
.Y(n_2492)
);

AOI221xp5_ASAP7_75t_L g2493 ( 
.A1(n_2459),
.A2(n_237),
.B1(n_234),
.B2(n_236),
.C(n_238),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2446),
.Y(n_2494)
);

NAND3xp33_ASAP7_75t_SL g2495 ( 
.A(n_2465),
.B(n_236),
.C(n_238),
.Y(n_2495)
);

AOI211xp5_ASAP7_75t_L g2496 ( 
.A1(n_2462),
.A2(n_241),
.B(n_239),
.C(n_240),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2478),
.Y(n_2497)
);

NOR2xp67_ASAP7_75t_L g2498 ( 
.A(n_2449),
.B(n_239),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2481),
.Y(n_2499)
);

NAND3xp33_ASAP7_75t_SL g2500 ( 
.A(n_2457),
.B(n_240),
.C(n_241),
.Y(n_2500)
);

NOR4xp25_ASAP7_75t_L g2501 ( 
.A(n_2447),
.B(n_244),
.C(n_242),
.D(n_243),
.Y(n_2501)
);

NAND4xp25_ASAP7_75t_SL g2502 ( 
.A(n_2469),
.B(n_245),
.C(n_243),
.D(n_244),
.Y(n_2502)
);

NOR3xp33_ASAP7_75t_SL g2503 ( 
.A(n_2479),
.B(n_245),
.C(n_246),
.Y(n_2503)
);

NAND4xp25_ASAP7_75t_L g2504 ( 
.A(n_2463),
.B(n_2455),
.C(n_2480),
.D(n_2461),
.Y(n_2504)
);

NAND4xp25_ASAP7_75t_L g2505 ( 
.A(n_2452),
.B(n_248),
.C(n_246),
.D(n_247),
.Y(n_2505)
);

NOR4xp25_ASAP7_75t_L g2506 ( 
.A(n_2471),
.B(n_249),
.C(n_247),
.D(n_248),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2456),
.B(n_250),
.Y(n_2507)
);

NAND4xp25_ASAP7_75t_L g2508 ( 
.A(n_2451),
.B(n_252),
.C(n_250),
.D(n_251),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_L g2509 ( 
.A(n_2453),
.B(n_251),
.Y(n_2509)
);

AOI221x1_ASAP7_75t_L g2510 ( 
.A1(n_2477),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.C(n_255),
.Y(n_2510)
);

NOR2x1_ASAP7_75t_L g2511 ( 
.A(n_2473),
.B(n_253),
.Y(n_2511)
);

NOR2xp67_ASAP7_75t_SL g2512 ( 
.A(n_2445),
.B(n_254),
.Y(n_2512)
);

NOR3xp33_ASAP7_75t_L g2513 ( 
.A(n_2474),
.B(n_255),
.C(n_256),
.Y(n_2513)
);

NOR2xp67_ASAP7_75t_L g2514 ( 
.A(n_2473),
.B(n_257),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2446),
.B(n_257),
.Y(n_2515)
);

OAI211xp5_ASAP7_75t_L g2516 ( 
.A1(n_2454),
.A2(n_260),
.B(n_258),
.C(n_259),
.Y(n_2516)
);

NAND4xp25_ASAP7_75t_SL g2517 ( 
.A(n_2464),
.B(n_261),
.C(n_258),
.D(n_259),
.Y(n_2517)
);

NOR3x1_ASAP7_75t_L g2518 ( 
.A(n_2449),
.B(n_261),
.C(n_262),
.Y(n_2518)
);

NOR3xp33_ASAP7_75t_L g2519 ( 
.A(n_2474),
.B(n_262),
.C(n_263),
.Y(n_2519)
);

BUFx2_ASAP7_75t_L g2520 ( 
.A(n_2446),
.Y(n_2520)
);

NOR2x1_ASAP7_75t_L g2521 ( 
.A(n_2473),
.B(n_264),
.Y(n_2521)
);

NOR2x1_ASAP7_75t_L g2522 ( 
.A(n_2473),
.B(n_265),
.Y(n_2522)
);

OAI221xp5_ASAP7_75t_L g2523 ( 
.A1(n_2454),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.C(n_268),
.Y(n_2523)
);

NOR3xp33_ASAP7_75t_L g2524 ( 
.A(n_2474),
.B(n_267),
.C(n_268),
.Y(n_2524)
);

NAND3xp33_ASAP7_75t_SL g2525 ( 
.A(n_2454),
.B(n_269),
.C(n_271),
.Y(n_2525)
);

AOI222xp33_ASAP7_75t_L g2526 ( 
.A1(n_2445),
.A2(n_269),
.B1(n_272),
.B2(n_273),
.C1(n_274),
.C2(n_275),
.Y(n_2526)
);

NAND4xp25_ASAP7_75t_L g2527 ( 
.A(n_2472),
.B(n_277),
.C(n_274),
.D(n_276),
.Y(n_2527)
);

OAI321xp33_ASAP7_75t_L g2528 ( 
.A1(n_2450),
.A2(n_277),
.A3(n_278),
.B1(n_279),
.B2(n_280),
.C(n_281),
.Y(n_2528)
);

AOI221xp5_ASAP7_75t_L g2529 ( 
.A1(n_2454),
.A2(n_283),
.B1(n_278),
.B2(n_279),
.C(n_284),
.Y(n_2529)
);

OAI211xp5_ASAP7_75t_L g2530 ( 
.A1(n_2454),
.A2(n_286),
.B(n_284),
.C(n_285),
.Y(n_2530)
);

XOR2xp5_ASAP7_75t_L g2531 ( 
.A(n_2467),
.B(n_285),
.Y(n_2531)
);

NOR2x1_ASAP7_75t_L g2532 ( 
.A(n_2473),
.B(n_287),
.Y(n_2532)
);

NAND3xp33_ASAP7_75t_SL g2533 ( 
.A(n_2454),
.B(n_287),
.C(n_289),
.Y(n_2533)
);

NOR2x1_ASAP7_75t_L g2534 ( 
.A(n_2473),
.B(n_289),
.Y(n_2534)
);

AOI211xp5_ASAP7_75t_L g2535 ( 
.A1(n_2454),
.A2(n_293),
.B(n_290),
.C(n_291),
.Y(n_2535)
);

NAND4xp75_ASAP7_75t_L g2536 ( 
.A(n_2450),
.B(n_295),
.C(n_291),
.D(n_293),
.Y(n_2536)
);

NAND3xp33_ASAP7_75t_L g2537 ( 
.A(n_2445),
.B(n_295),
.C(n_296),
.Y(n_2537)
);

OA211x2_ASAP7_75t_L g2538 ( 
.A1(n_2479),
.A2(n_298),
.B(n_296),
.C(n_297),
.Y(n_2538)
);

NOR2x1_ASAP7_75t_L g2539 ( 
.A(n_2473),
.B(n_298),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2499),
.B(n_299),
.Y(n_2540)
);

AOI22xp5_ASAP7_75t_L g2541 ( 
.A1(n_2492),
.A2(n_2514),
.B1(n_2494),
.B2(n_2483),
.Y(n_2541)
);

NOR2xp33_ASAP7_75t_R g2542 ( 
.A(n_2525),
.B(n_299),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2520),
.B(n_300),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_SL g2544 ( 
.A(n_2488),
.B(n_301),
.Y(n_2544)
);

NAND2xp33_ASAP7_75t_R g2545 ( 
.A(n_2503),
.B(n_301),
.Y(n_2545)
);

CKINVDCx16_ASAP7_75t_R g2546 ( 
.A(n_2533),
.Y(n_2546)
);

AOI222xp33_ASAP7_75t_L g2547 ( 
.A1(n_2497),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.C1(n_306),
.C2(n_307),
.Y(n_2547)
);

BUFx2_ASAP7_75t_L g2548 ( 
.A(n_2515),
.Y(n_2548)
);

XNOR2xp5_ASAP7_75t_L g2549 ( 
.A(n_2487),
.B(n_302),
.Y(n_2549)
);

AOI322xp5_ASAP7_75t_L g2550 ( 
.A1(n_2489),
.A2(n_2090),
.A3(n_2080),
.B1(n_308),
.B2(n_309),
.C1(n_310),
.C2(n_311),
.Y(n_2550)
);

OAI322xp33_ASAP7_75t_L g2551 ( 
.A1(n_2507),
.A2(n_303),
.A3(n_307),
.B1(n_308),
.B2(n_309),
.C1(n_311),
.C2(n_312),
.Y(n_2551)
);

XOR2xp5_ASAP7_75t_L g2552 ( 
.A(n_2531),
.B(n_313),
.Y(n_2552)
);

OAI22xp33_ASAP7_75t_L g2553 ( 
.A1(n_2527),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_2553)
);

INVx2_ASAP7_75t_SL g2554 ( 
.A(n_2490),
.Y(n_2554)
);

AOI221x1_ASAP7_75t_L g2555 ( 
.A1(n_2513),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.C(n_318),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2491),
.Y(n_2556)
);

AOI22xp5_ASAP7_75t_L g2557 ( 
.A1(n_2511),
.A2(n_2113),
.B1(n_2103),
.B2(n_2098),
.Y(n_2557)
);

AOI21x1_ASAP7_75t_L g2558 ( 
.A1(n_2512),
.A2(n_316),
.B(n_319),
.Y(n_2558)
);

AOI22xp5_ASAP7_75t_L g2559 ( 
.A1(n_2521),
.A2(n_2231),
.B1(n_2218),
.B2(n_321),
.Y(n_2559)
);

HB1xp67_ASAP7_75t_L g2560 ( 
.A(n_2498),
.Y(n_2560)
);

NAND4xp75_ASAP7_75t_L g2561 ( 
.A(n_2518),
.B(n_2484),
.C(n_2538),
.D(n_2532),
.Y(n_2561)
);

AOI211xp5_ASAP7_75t_L g2562 ( 
.A1(n_2523),
.A2(n_323),
.B(n_319),
.C(n_320),
.Y(n_2562)
);

AOI22xp33_ASAP7_75t_L g2563 ( 
.A1(n_2522),
.A2(n_2539),
.B1(n_2534),
.B2(n_2500),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2509),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2501),
.B(n_323),
.Y(n_2565)
);

INVxp33_ASAP7_75t_L g2566 ( 
.A(n_2519),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2535),
.B(n_324),
.Y(n_2567)
);

NAND3xp33_ASAP7_75t_L g2568 ( 
.A(n_2529),
.B(n_324),
.C(n_325),
.Y(n_2568)
);

OAI21xp33_ASAP7_75t_L g2569 ( 
.A1(n_2504),
.A2(n_325),
.B(n_326),
.Y(n_2569)
);

HB1xp67_ASAP7_75t_L g2570 ( 
.A(n_2536),
.Y(n_2570)
);

NOR4xp25_ASAP7_75t_L g2571 ( 
.A(n_2482),
.B(n_328),
.C(n_326),
.D(n_327),
.Y(n_2571)
);

O2A1O1Ixp33_ASAP7_75t_L g2572 ( 
.A1(n_2486),
.A2(n_2516),
.B(n_2530),
.C(n_2485),
.Y(n_2572)
);

INVx1_ASAP7_75t_SL g2573 ( 
.A(n_2537),
.Y(n_2573)
);

AND2x4_ASAP7_75t_L g2574 ( 
.A(n_2524),
.B(n_327),
.Y(n_2574)
);

NOR2xp33_ASAP7_75t_L g2575 ( 
.A(n_2495),
.B(n_328),
.Y(n_2575)
);

BUFx3_ASAP7_75t_L g2576 ( 
.A(n_2496),
.Y(n_2576)
);

NOR2x1_ASAP7_75t_L g2577 ( 
.A(n_2517),
.B(n_329),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2506),
.B(n_329),
.Y(n_2578)
);

OAI22xp5_ASAP7_75t_L g2579 ( 
.A1(n_2496),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.Y(n_2579)
);

HB1xp67_ASAP7_75t_L g2580 ( 
.A(n_2502),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_R g2581 ( 
.A(n_2528),
.B(n_330),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2508),
.Y(n_2582)
);

NOR2xp33_ASAP7_75t_R g2583 ( 
.A(n_2526),
.B(n_333),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2505),
.Y(n_2584)
);

OAI22xp33_ASAP7_75t_L g2585 ( 
.A1(n_2510),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_2585)
);

INVx1_ASAP7_75t_SL g2586 ( 
.A(n_2493),
.Y(n_2586)
);

AND2x2_ASAP7_75t_L g2587 ( 
.A(n_2499),
.B(n_335),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2520),
.B(n_336),
.Y(n_2588)
);

AOI22xp5_ASAP7_75t_L g2589 ( 
.A1(n_2499),
.A2(n_2231),
.B1(n_339),
.B2(n_337),
.Y(n_2589)
);

AOI21xp5_ASAP7_75t_L g2590 ( 
.A1(n_2507),
.A2(n_337),
.B(n_338),
.Y(n_2590)
);

AOI21xp33_ASAP7_75t_SL g2591 ( 
.A1(n_2487),
.A2(n_340),
.B(n_341),
.Y(n_2591)
);

OAI21xp5_ASAP7_75t_SL g2592 ( 
.A1(n_2487),
.A2(n_340),
.B(n_341),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2499),
.B(n_342),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_L g2594 ( 
.A(n_2520),
.B(n_342),
.Y(n_2594)
);

NOR2xp33_ASAP7_75t_R g2595 ( 
.A(n_2525),
.B(n_343),
.Y(n_2595)
);

HB1xp67_ASAP7_75t_L g2596 ( 
.A(n_2520),
.Y(n_2596)
);

NOR2x1_ASAP7_75t_L g2597 ( 
.A(n_2543),
.B(n_343),
.Y(n_2597)
);

NAND2x1p5_ASAP7_75t_L g2598 ( 
.A(n_2554),
.B(n_2576),
.Y(n_2598)
);

NOR2xp67_ASAP7_75t_L g2599 ( 
.A(n_2596),
.B(n_2579),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2558),
.Y(n_2600)
);

OR2x2_ASAP7_75t_L g2601 ( 
.A(n_2571),
.B(n_344),
.Y(n_2601)
);

NOR2x1_ASAP7_75t_L g2602 ( 
.A(n_2588),
.B(n_2592),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2560),
.Y(n_2603)
);

INVx3_ASAP7_75t_L g2604 ( 
.A(n_2561),
.Y(n_2604)
);

NAND4xp75_ASAP7_75t_L g2605 ( 
.A(n_2541),
.B(n_346),
.C(n_344),
.D(n_345),
.Y(n_2605)
);

OR2x6_ASAP7_75t_L g2606 ( 
.A(n_2548),
.B(n_345),
.Y(n_2606)
);

HB1xp67_ASAP7_75t_L g2607 ( 
.A(n_2549),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2546),
.B(n_346),
.Y(n_2608)
);

NOR2x1p5_ASAP7_75t_L g2609 ( 
.A(n_2565),
.B(n_347),
.Y(n_2609)
);

NOR2xp67_ASAP7_75t_L g2610 ( 
.A(n_2568),
.B(n_348),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2578),
.Y(n_2611)
);

NAND2x1p5_ASAP7_75t_L g2612 ( 
.A(n_2573),
.B(n_348),
.Y(n_2612)
);

NAND5xp2_ASAP7_75t_L g2613 ( 
.A(n_2563),
.B(n_349),
.C(n_350),
.D(n_351),
.E(n_352),
.Y(n_2613)
);

NAND4xp75_ASAP7_75t_L g2614 ( 
.A(n_2556),
.B(n_349),
.C(n_350),
.D(n_353),
.Y(n_2614)
);

INVxp67_ASAP7_75t_SL g2615 ( 
.A(n_2594),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2540),
.Y(n_2616)
);

AOI22xp5_ASAP7_75t_L g2617 ( 
.A1(n_2545),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2577),
.Y(n_2618)
);

NOR2xp33_ASAP7_75t_L g2619 ( 
.A(n_2591),
.B(n_354),
.Y(n_2619)
);

AND2x2_ASAP7_75t_L g2620 ( 
.A(n_2574),
.B(n_2570),
.Y(n_2620)
);

OAI22xp5_ASAP7_75t_L g2621 ( 
.A1(n_2566),
.A2(n_2580),
.B1(n_2586),
.B2(n_2567),
.Y(n_2621)
);

AO22x1_ASAP7_75t_L g2622 ( 
.A1(n_2587),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2593),
.Y(n_2623)
);

NAND4xp75_ASAP7_75t_L g2624 ( 
.A(n_2564),
.B(n_356),
.C(n_357),
.D(n_358),
.Y(n_2624)
);

INVx1_ASAP7_75t_SL g2625 ( 
.A(n_2581),
.Y(n_2625)
);

AND2x4_ASAP7_75t_L g2626 ( 
.A(n_2582),
.B(n_2584),
.Y(n_2626)
);

NOR2x1_ASAP7_75t_L g2627 ( 
.A(n_2551),
.B(n_358),
.Y(n_2627)
);

NOR2x1_ASAP7_75t_L g2628 ( 
.A(n_2552),
.B(n_359),
.Y(n_2628)
);

NOR2xp33_ASAP7_75t_L g2629 ( 
.A(n_2544),
.B(n_360),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2572),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2574),
.B(n_360),
.Y(n_2631)
);

NOR2x1_ASAP7_75t_L g2632 ( 
.A(n_2553),
.B(n_361),
.Y(n_2632)
);

NAND4xp75_ASAP7_75t_L g2633 ( 
.A(n_2555),
.B(n_361),
.C(n_362),
.D(n_363),
.Y(n_2633)
);

AND2x4_ASAP7_75t_L g2634 ( 
.A(n_2590),
.B(n_364),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2575),
.Y(n_2635)
);

XNOR2x1_ASAP7_75t_L g2636 ( 
.A(n_2585),
.B(n_2559),
.Y(n_2636)
);

OAI221xp5_ASAP7_75t_L g2637 ( 
.A1(n_2569),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.C(n_369),
.Y(n_2637)
);

AND2x4_ASAP7_75t_L g2638 ( 
.A(n_2589),
.B(n_367),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2542),
.Y(n_2639)
);

INVx3_ASAP7_75t_L g2640 ( 
.A(n_2595),
.Y(n_2640)
);

NOR2x1_ASAP7_75t_L g2641 ( 
.A(n_2547),
.B(n_368),
.Y(n_2641)
);

XOR2x2_ASAP7_75t_L g2642 ( 
.A(n_2562),
.B(n_369),
.Y(n_2642)
);

NAND4xp75_ASAP7_75t_L g2643 ( 
.A(n_2583),
.B(n_370),
.C(n_371),
.D(n_372),
.Y(n_2643)
);

NOR2xp67_ASAP7_75t_L g2644 ( 
.A(n_2557),
.B(n_370),
.Y(n_2644)
);

OA211x2_ASAP7_75t_L g2645 ( 
.A1(n_2629),
.A2(n_2550),
.B(n_372),
.C(n_373),
.Y(n_2645)
);

NAND4xp75_ASAP7_75t_L g2646 ( 
.A(n_2599),
.B(n_371),
.C(n_373),
.D(n_374),
.Y(n_2646)
);

NOR3xp33_ASAP7_75t_L g2647 ( 
.A(n_2603),
.B(n_375),
.C(n_376),
.Y(n_2647)
);

OR2x2_ASAP7_75t_L g2648 ( 
.A(n_2598),
.B(n_2612),
.Y(n_2648)
);

NOR3xp33_ASAP7_75t_SL g2649 ( 
.A(n_2621),
.B(n_375),
.C(n_376),
.Y(n_2649)
);

OAI21xp33_ASAP7_75t_L g2650 ( 
.A1(n_2613),
.A2(n_377),
.B(n_378),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2600),
.B(n_378),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2609),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2604),
.B(n_379),
.Y(n_2653)
);

AND3x2_ASAP7_75t_L g2654 ( 
.A(n_2618),
.B(n_379),
.C(n_380),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2628),
.Y(n_2655)
);

NOR2x1_ASAP7_75t_L g2656 ( 
.A(n_2630),
.B(n_380),
.Y(n_2656)
);

NAND3xp33_ASAP7_75t_SL g2657 ( 
.A(n_2625),
.B(n_381),
.C(n_382),
.Y(n_2657)
);

NAND5xp2_ASAP7_75t_L g2658 ( 
.A(n_2620),
.B(n_381),
.C(n_383),
.D(n_384),
.E(n_385),
.Y(n_2658)
);

NOR3xp33_ASAP7_75t_SL g2659 ( 
.A(n_2615),
.B(n_383),
.C(n_384),
.Y(n_2659)
);

NAND5xp2_ASAP7_75t_L g2660 ( 
.A(n_2616),
.B(n_385),
.C(n_386),
.D(n_387),
.E(n_388),
.Y(n_2660)
);

NAND4xp25_ASAP7_75t_L g2661 ( 
.A(n_2617),
.B(n_386),
.C(n_387),
.D(n_388),
.Y(n_2661)
);

OR3x2_ASAP7_75t_L g2662 ( 
.A(n_2611),
.B(n_389),
.C(n_391),
.Y(n_2662)
);

NAND4xp25_ASAP7_75t_SL g2663 ( 
.A(n_2637),
.B(n_389),
.C(n_391),
.D(n_392),
.Y(n_2663)
);

AND5x1_ASAP7_75t_L g2664 ( 
.A(n_2619),
.B(n_392),
.C(n_393),
.D(n_394),
.E(n_395),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2597),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2640),
.B(n_2623),
.Y(n_2666)
);

NOR4xp25_ASAP7_75t_L g2667 ( 
.A(n_2639),
.B(n_393),
.C(n_394),
.D(n_395),
.Y(n_2667)
);

NAND5xp2_ASAP7_75t_L g2668 ( 
.A(n_2635),
.B(n_396),
.C(n_397),
.D(n_398),
.E(n_399),
.Y(n_2668)
);

AND4x1_ASAP7_75t_L g2669 ( 
.A(n_2602),
.B(n_396),
.C(n_397),
.D(n_398),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2601),
.Y(n_2670)
);

NOR5xp2_ASAP7_75t_L g2671 ( 
.A(n_2607),
.B(n_399),
.C(n_400),
.D(n_401),
.E(n_402),
.Y(n_2671)
);

NAND3xp33_ASAP7_75t_L g2672 ( 
.A(n_2608),
.B(n_2606),
.C(n_2626),
.Y(n_2672)
);

NAND4xp25_ASAP7_75t_L g2673 ( 
.A(n_2610),
.B(n_400),
.C(n_401),
.D(n_402),
.Y(n_2673)
);

NOR5xp2_ASAP7_75t_L g2674 ( 
.A(n_2643),
.B(n_403),
.C(n_404),
.D(n_405),
.E(n_406),
.Y(n_2674)
);

NOR2x1_ASAP7_75t_L g2675 ( 
.A(n_2606),
.B(n_403),
.Y(n_2675)
);

AOI211xp5_ASAP7_75t_L g2676 ( 
.A1(n_2622),
.A2(n_405),
.B(n_406),
.C(n_407),
.Y(n_2676)
);

NOR5xp2_ASAP7_75t_L g2677 ( 
.A(n_2636),
.B(n_407),
.C(n_408),
.D(n_409),
.E(n_410),
.Y(n_2677)
);

INVxp67_ASAP7_75t_SL g2678 ( 
.A(n_2631),
.Y(n_2678)
);

OAI211xp5_ASAP7_75t_SL g2679 ( 
.A1(n_2627),
.A2(n_408),
.B(n_409),
.C(n_410),
.Y(n_2679)
);

NAND5xp2_ASAP7_75t_L g2680 ( 
.A(n_2642),
.B(n_411),
.C(n_412),
.D(n_413),
.E(n_415),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2633),
.Y(n_2681)
);

NAND4xp75_ASAP7_75t_L g2682 ( 
.A(n_2641),
.B(n_2632),
.C(n_2644),
.D(n_2624),
.Y(n_2682)
);

NOR2x1_ASAP7_75t_L g2683 ( 
.A(n_2605),
.B(n_412),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2648),
.Y(n_2684)
);

CKINVDCx5p33_ASAP7_75t_R g2685 ( 
.A(n_2678),
.Y(n_2685)
);

BUFx2_ASAP7_75t_L g2686 ( 
.A(n_2675),
.Y(n_2686)
);

OAI221xp5_ASAP7_75t_L g2687 ( 
.A1(n_2667),
.A2(n_2605),
.B1(n_2614),
.B2(n_2634),
.C(n_2638),
.Y(n_2687)
);

NAND3xp33_ASAP7_75t_L g2688 ( 
.A(n_2672),
.B(n_413),
.C(n_415),
.Y(n_2688)
);

CKINVDCx20_ASAP7_75t_R g2689 ( 
.A(n_2666),
.Y(n_2689)
);

NOR2xp33_ASAP7_75t_R g2690 ( 
.A(n_2681),
.B(n_416),
.Y(n_2690)
);

CKINVDCx5p33_ASAP7_75t_R g2691 ( 
.A(n_2652),
.Y(n_2691)
);

CKINVDCx5p33_ASAP7_75t_R g2692 ( 
.A(n_2670),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2659),
.B(n_417),
.Y(n_2693)
);

INVx6_ASAP7_75t_L g2694 ( 
.A(n_2655),
.Y(n_2694)
);

OR2x2_ASAP7_75t_L g2695 ( 
.A(n_2665),
.B(n_418),
.Y(n_2695)
);

CKINVDCx5p33_ASAP7_75t_R g2696 ( 
.A(n_2649),
.Y(n_2696)
);

CKINVDCx20_ASAP7_75t_R g2697 ( 
.A(n_2664),
.Y(n_2697)
);

XOR2xp5_ASAP7_75t_L g2698 ( 
.A(n_2662),
.B(n_2682),
.Y(n_2698)
);

NOR2xp33_ASAP7_75t_L g2699 ( 
.A(n_2680),
.B(n_418),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2654),
.Y(n_2700)
);

CKINVDCx16_ASAP7_75t_R g2701 ( 
.A(n_2656),
.Y(n_2701)
);

BUFx6f_ASAP7_75t_L g2702 ( 
.A(n_2651),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2653),
.Y(n_2703)
);

BUFx2_ASAP7_75t_L g2704 ( 
.A(n_2683),
.Y(n_2704)
);

INVx1_ASAP7_75t_SL g2705 ( 
.A(n_2646),
.Y(n_2705)
);

BUFx2_ASAP7_75t_L g2706 ( 
.A(n_2673),
.Y(n_2706)
);

CKINVDCx5p33_ASAP7_75t_R g2707 ( 
.A(n_2650),
.Y(n_2707)
);

INVxp33_ASAP7_75t_L g2708 ( 
.A(n_2647),
.Y(n_2708)
);

AOI22x1_ASAP7_75t_L g2709 ( 
.A1(n_2684),
.A2(n_2671),
.B1(n_2677),
.B2(n_2674),
.Y(n_2709)
);

AOI22xp33_ASAP7_75t_L g2710 ( 
.A1(n_2694),
.A2(n_2679),
.B1(n_2645),
.B2(n_2657),
.Y(n_2710)
);

NAND3xp33_ASAP7_75t_SL g2711 ( 
.A(n_2689),
.B(n_2676),
.C(n_2669),
.Y(n_2711)
);

AOI322xp5_ASAP7_75t_L g2712 ( 
.A1(n_2697),
.A2(n_2663),
.A3(n_2661),
.B1(n_2658),
.B2(n_2660),
.C1(n_2668),
.C2(n_425),
.Y(n_2712)
);

AOI322xp5_ASAP7_75t_L g2713 ( 
.A1(n_2699),
.A2(n_419),
.A3(n_420),
.B1(n_421),
.B2(n_422),
.C1(n_423),
.C2(n_426),
.Y(n_2713)
);

AND2x4_ASAP7_75t_L g2714 ( 
.A(n_2686),
.B(n_419),
.Y(n_2714)
);

NAND3xp33_ASAP7_75t_SL g2715 ( 
.A(n_2685),
.B(n_420),
.C(n_421),
.Y(n_2715)
);

INVx2_ASAP7_75t_SL g2716 ( 
.A(n_2694),
.Y(n_2716)
);

OR3x1_ASAP7_75t_L g2717 ( 
.A(n_2703),
.B(n_422),
.C(n_423),
.Y(n_2717)
);

AOI22xp33_ASAP7_75t_SL g2718 ( 
.A1(n_2701),
.A2(n_426),
.B1(n_427),
.B2(n_428),
.Y(n_2718)
);

AOI22x1_ASAP7_75t_L g2719 ( 
.A1(n_2698),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.Y(n_2719)
);

AOI322xp5_ASAP7_75t_L g2720 ( 
.A1(n_2704),
.A2(n_429),
.A3(n_430),
.B1(n_432),
.B2(n_433),
.C1(n_434),
.C2(n_435),
.Y(n_2720)
);

AOI32xp33_ASAP7_75t_L g2721 ( 
.A1(n_2693),
.A2(n_2692),
.A3(n_2708),
.B1(n_2691),
.B2(n_2705),
.Y(n_2721)
);

AOI322xp5_ASAP7_75t_L g2722 ( 
.A1(n_2700),
.A2(n_430),
.A3(n_432),
.B1(n_433),
.B2(n_434),
.C1(n_437),
.C2(n_438),
.Y(n_2722)
);

INVx1_ASAP7_75t_SL g2723 ( 
.A(n_2690),
.Y(n_2723)
);

AOI22xp33_ASAP7_75t_L g2724 ( 
.A1(n_2702),
.A2(n_438),
.B1(n_439),
.B2(n_440),
.Y(n_2724)
);

OAI322xp33_ASAP7_75t_L g2725 ( 
.A1(n_2687),
.A2(n_440),
.A3(n_441),
.B1(n_442),
.B2(n_443),
.C1(n_444),
.C2(n_446),
.Y(n_2725)
);

AOI322xp5_ASAP7_75t_L g2726 ( 
.A1(n_2696),
.A2(n_443),
.A3(n_444),
.B1(n_446),
.B2(n_447),
.C1(n_448),
.C2(n_449),
.Y(n_2726)
);

OAI211xp5_ASAP7_75t_SL g2727 ( 
.A1(n_2702),
.A2(n_448),
.B(n_450),
.C(n_451),
.Y(n_2727)
);

O2A1O1Ixp33_ASAP7_75t_L g2728 ( 
.A1(n_2706),
.A2(n_451),
.B(n_452),
.C(n_453),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2716),
.Y(n_2729)
);

OAI22x1_ASAP7_75t_L g2730 ( 
.A1(n_2709),
.A2(n_2707),
.B1(n_2688),
.B2(n_2695),
.Y(n_2730)
);

OAI22x1_ASAP7_75t_L g2731 ( 
.A1(n_2719),
.A2(n_2702),
.B1(n_453),
.B2(n_454),
.Y(n_2731)
);

AOI22xp5_ASAP7_75t_L g2732 ( 
.A1(n_2711),
.A2(n_452),
.B1(n_454),
.B2(n_455),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2717),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2714),
.Y(n_2734)
);

OAI22x1_ASAP7_75t_L g2735 ( 
.A1(n_2723),
.A2(n_455),
.B1(n_456),
.B2(n_457),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2710),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2715),
.Y(n_2737)
);

OAI22x1_ASAP7_75t_L g2738 ( 
.A1(n_2714),
.A2(n_456),
.B1(n_457),
.B2(n_458),
.Y(n_2738)
);

OAI22x1_ASAP7_75t_L g2739 ( 
.A1(n_2721),
.A2(n_459),
.B1(n_460),
.B2(n_461),
.Y(n_2739)
);

CKINVDCx20_ASAP7_75t_R g2740 ( 
.A(n_2712),
.Y(n_2740)
);

NAND3xp33_ASAP7_75t_L g2741 ( 
.A(n_2729),
.B(n_2713),
.C(n_2718),
.Y(n_2741)
);

AOI221xp5_ASAP7_75t_L g2742 ( 
.A1(n_2733),
.A2(n_2736),
.B1(n_2730),
.B2(n_2731),
.C(n_2737),
.Y(n_2742)
);

NOR4xp25_ASAP7_75t_L g2743 ( 
.A(n_2734),
.B(n_2727),
.C(n_2728),
.D(n_2725),
.Y(n_2743)
);

NOR2x1p5_ASAP7_75t_L g2744 ( 
.A(n_2740),
.B(n_2724),
.Y(n_2744)
);

NOR4xp25_ASAP7_75t_L g2745 ( 
.A(n_2739),
.B(n_2722),
.C(n_2726),
.D(n_2720),
.Y(n_2745)
);

XNOR2xp5_ASAP7_75t_L g2746 ( 
.A(n_2738),
.B(n_459),
.Y(n_2746)
);

AOI22xp5_ASAP7_75t_L g2747 ( 
.A1(n_2735),
.A2(n_462),
.B1(n_463),
.B2(n_464),
.Y(n_2747)
);

HB1xp67_ASAP7_75t_L g2748 ( 
.A(n_2744),
.Y(n_2748)
);

AO21x2_ASAP7_75t_L g2749 ( 
.A1(n_2741),
.A2(n_2732),
.B(n_463),
.Y(n_2749)
);

NOR2xp33_ASAP7_75t_R g2750 ( 
.A(n_2746),
.B(n_462),
.Y(n_2750)
);

NAND2x1p5_ASAP7_75t_L g2751 ( 
.A(n_2742),
.B(n_465),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2747),
.Y(n_2752)
);

NAND2xp33_ASAP7_75t_SL g2753 ( 
.A(n_2743),
.B(n_465),
.Y(n_2753)
);

XNOR2x1_ASAP7_75t_L g2754 ( 
.A(n_2748),
.B(n_2745),
.Y(n_2754)
);

AOI22xp5_ASAP7_75t_L g2755 ( 
.A1(n_2753),
.A2(n_466),
.B1(n_467),
.B2(n_468),
.Y(n_2755)
);

NOR2xp33_ASAP7_75t_L g2756 ( 
.A(n_2751),
.B(n_466),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2752),
.B(n_467),
.Y(n_2757)
);

AOI22xp33_ASAP7_75t_L g2758 ( 
.A1(n_2754),
.A2(n_2750),
.B1(n_2749),
.B2(n_470),
.Y(n_2758)
);

OAI22xp5_ASAP7_75t_L g2759 ( 
.A1(n_2755),
.A2(n_468),
.B1(n_469),
.B2(n_471),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2756),
.B(n_469),
.Y(n_2760)
);

AOI22xp5_ASAP7_75t_SL g2761 ( 
.A1(n_2757),
.A2(n_471),
.B1(n_472),
.B2(n_473),
.Y(n_2761)
);

OAI21x1_ASAP7_75t_SL g2762 ( 
.A1(n_2754),
.A2(n_473),
.B(n_474),
.Y(n_2762)
);

AOI22xp5_ASAP7_75t_L g2763 ( 
.A1(n_2758),
.A2(n_2760),
.B1(n_2759),
.B2(n_2761),
.Y(n_2763)
);

OAI21x1_ASAP7_75t_L g2764 ( 
.A1(n_2762),
.A2(n_474),
.B(n_475),
.Y(n_2764)
);

AO21x1_ASAP7_75t_L g2765 ( 
.A1(n_2760),
.A2(n_475),
.B(n_476),
.Y(n_2765)
);

OAI21xp5_ASAP7_75t_L g2766 ( 
.A1(n_2758),
.A2(n_476),
.B(n_477),
.Y(n_2766)
);

AOI22xp5_ASAP7_75t_L g2767 ( 
.A1(n_2765),
.A2(n_478),
.B1(n_479),
.B2(n_480),
.Y(n_2767)
);

AOI22xp5_ASAP7_75t_L g2768 ( 
.A1(n_2763),
.A2(n_481),
.B1(n_482),
.B2(n_483),
.Y(n_2768)
);

AO22x2_ASAP7_75t_L g2769 ( 
.A1(n_2766),
.A2(n_481),
.B1(n_483),
.B2(n_484),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2767),
.B(n_2764),
.Y(n_2770)
);

OAI21xp5_ASAP7_75t_L g2771 ( 
.A1(n_2768),
.A2(n_485),
.B(n_486),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2770),
.Y(n_2772)
);

AOI221x1_ASAP7_75t_L g2773 ( 
.A1(n_2772),
.A2(n_2769),
.B1(n_2771),
.B2(n_487),
.C(n_488),
.Y(n_2773)
);

AOI21xp5_ASAP7_75t_L g2774 ( 
.A1(n_2773),
.A2(n_485),
.B(n_486),
.Y(n_2774)
);

AOI211xp5_ASAP7_75t_L g2775 ( 
.A1(n_2774),
.A2(n_489),
.B(n_490),
.C(n_491),
.Y(n_2775)
);


endmodule