module fake_jpeg_30603_n_495 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_495);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_495;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g51 ( 
.A(n_22),
.B(n_13),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_51),
.B(n_54),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

NAND2xp33_ASAP7_75t_SL g54 ( 
.A(n_22),
.B(n_13),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

HAxp5_ASAP7_75t_SL g57 ( 
.A(n_22),
.B(n_0),
.CON(n_57),
.SN(n_57)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_57),
.B(n_72),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_26),
.B(n_13),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_26),
.B(n_10),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_73),
.Y(n_104)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_SL g72 ( 
.A(n_22),
.B(n_45),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_75),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_80),
.Y(n_118)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_45),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_91),
.Y(n_130)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVxp67_ASAP7_75t_SL g131 ( 
.A(n_90),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_27),
.B(n_10),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_38),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_94),
.Y(n_146)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_93),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_42),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_43),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

BUFx24_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVxp67_ASAP7_75t_SL g173 ( 
.A(n_107),
.Y(n_173)
);

INVx6_ASAP7_75t_SL g112 ( 
.A(n_85),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_112),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_70),
.B(n_27),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_123),
.B(n_143),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_124),
.Y(n_188)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_93),
.A2(n_40),
.B1(n_21),
.B2(n_44),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_46),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_87),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_142),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_59),
.A2(n_44),
.B1(n_28),
.B2(n_48),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_134),
.A2(n_140),
.B1(n_52),
.B2(n_55),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_84),
.A2(n_40),
.B1(n_31),
.B2(n_41),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_67),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_62),
.B(n_19),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_63),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_90),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_97),
.B(n_19),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_158),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_99),
.B(n_24),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_159),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_161),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_162),
.B(n_178),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_43),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_163),
.B(n_167),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_107),
.A2(n_58),
.B1(n_81),
.B2(n_50),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_164),
.A2(n_172),
.B1(n_193),
.B2(n_197),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_165),
.B(n_212),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_166),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_49),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_170),
.Y(n_249)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_171),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_134),
.A2(n_78),
.B1(n_77),
.B2(n_48),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_174),
.A2(n_179),
.B1(n_182),
.B2(n_213),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_153),
.A2(n_76),
.B1(n_61),
.B2(n_53),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_175),
.A2(n_116),
.B1(n_129),
.B2(n_4),
.Y(n_258)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_177),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_108),
.A2(n_66),
.B1(n_63),
.B2(n_49),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_145),
.A2(n_66),
.B1(n_49),
.B2(n_90),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_118),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_194),
.Y(n_228)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_185),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_100),
.Y(n_186)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_186),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_102),
.Y(n_189)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_189),
.Y(n_246)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_138),
.Y(n_190)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_190),
.Y(n_252)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_118),
.Y(n_192)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_192),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_117),
.A2(n_46),
.B1(n_41),
.B2(n_39),
.Y(n_193)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_103),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_200),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_113),
.A2(n_46),
.B1(n_41),
.B2(n_39),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_198),
.A2(n_204),
.B1(n_215),
.B2(n_115),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_151),
.A2(n_47),
.B1(n_49),
.B2(n_24),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_199),
.A2(n_202),
.B1(n_214),
.B2(n_181),
.Y(n_242)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_120),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_151),
.A2(n_47),
.B1(n_8),
.B2(n_2),
.Y(n_202)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_208),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_101),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_104),
.B(n_8),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_205),
.B(n_206),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_104),
.B(n_8),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_130),
.B(n_0),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_207),
.B(n_211),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_130),
.B(n_0),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_105),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_209),
.B(n_210),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_101),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_149),
.B(n_1),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_113),
.B(n_1),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_137),
.A2(n_114),
.B1(n_141),
.B2(n_103),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_153),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_152),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_128),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_216),
.B(n_218),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_202),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_173),
.B(n_132),
.C(n_154),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_222),
.B(n_225),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_1),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_232),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_136),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g232 ( 
.A(n_160),
.Y(n_232)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_173),
.B(n_124),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_236),
.B(n_240),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_165),
.B(n_136),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_164),
.B(n_131),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_254),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_242),
.A2(n_250),
.B1(n_213),
.B2(n_159),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g244 ( 
.A1(n_174),
.A2(n_141),
.B1(n_148),
.B2(n_128),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_244),
.A2(n_258),
.B1(n_170),
.B2(n_204),
.Y(n_272)
);

AOI21xp33_ASAP7_75t_L g245 ( 
.A1(n_182),
.A2(n_2),
.B(n_3),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_245),
.B(n_3),
.Y(n_296)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_247),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_175),
.A2(n_115),
.B1(n_135),
.B2(n_133),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_248),
.A2(n_260),
.B1(n_161),
.B2(n_198),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_176),
.A2(n_106),
.B1(n_148),
.B2(n_116),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_169),
.B(n_135),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_195),
.B(n_133),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_257),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_179),
.B(n_106),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_200),
.A2(n_129),
.B1(n_3),
.B2(n_5),
.Y(n_260)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_219),
.B(n_256),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_264),
.B(n_270),
.Y(n_325)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_254),
.Y(n_265)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_268),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_261),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_177),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_271),
.B(n_280),
.Y(n_331)
);

OA22x2_ASAP7_75t_L g317 ( 
.A1(n_272),
.A2(n_227),
.B1(n_243),
.B2(n_249),
.Y(n_317)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_203),
.B1(n_184),
.B2(n_194),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_235),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_228),
.B(n_188),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_220),
.Y(n_281)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_226),
.Y(n_282)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_234),
.B(n_178),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_283),
.B(n_287),
.Y(n_336)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_226),
.Y(n_284)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_284),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_233),
.A2(n_166),
.B1(n_187),
.B2(n_186),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_285),
.A2(n_289),
.B1(n_244),
.B2(n_258),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_216),
.B(n_218),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_288),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_231),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_225),
.B(n_185),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_233),
.A2(n_210),
.B1(n_178),
.B2(n_191),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_230),
.B(n_185),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_290),
.B(n_295),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_239),
.B(n_210),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_297),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_217),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_293),
.Y(n_320)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_246),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_294),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_222),
.B(n_2),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_296),
.A2(n_221),
.B(n_236),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_229),
.B(n_5),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_259),
.B(n_5),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_298),
.B(n_300),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_240),
.A2(n_5),
.B(n_7),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_299),
.A2(n_223),
.B(n_252),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_243),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_242),
.B(n_7),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_301),
.B(n_223),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_240),
.B(n_257),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_302),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_303),
.A2(n_314),
.B1(n_317),
.B2(n_330),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_266),
.A2(n_224),
.B1(n_241),
.B2(n_221),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_307),
.A2(n_326),
.B1(n_333),
.B2(n_329),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_322),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_273),
.B(n_221),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_316),
.B(n_324),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_268),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_323),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_273),
.B(n_236),
.C(n_246),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_266),
.A2(n_227),
.B1(n_249),
.B2(n_235),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_285),
.A2(n_289),
.B1(n_301),
.B2(n_274),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_332),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_329),
.A2(n_278),
.B(n_302),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_272),
.A2(n_252),
.B1(n_237),
.B2(n_238),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_278),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_237),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_269),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_290),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_337),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_293),
.B(n_238),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_288),
.B(n_279),
.Y(n_338)
);

XNOR2x1_ASAP7_75t_L g370 ( 
.A(n_338),
.B(n_295),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_263),
.B(n_270),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_339),
.B(n_287),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_341),
.B(n_305),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_343),
.Y(n_392)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_344),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_370),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_286),
.Y(n_346)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_346),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_308),
.B(n_265),
.Y(n_348)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_348),
.Y(n_384)
);

INVx13_ASAP7_75t_L g349 ( 
.A(n_309),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_349),
.Y(n_387)
);

BUFx5_ASAP7_75t_L g350 ( 
.A(n_320),
.Y(n_350)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_350),
.Y(n_386)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_319),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_351),
.Y(n_385)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_334),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_357),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_304),
.A2(n_296),
.B(n_278),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_360),
.Y(n_374)
);

OAI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_312),
.A2(n_308),
.B1(n_310),
.B2(n_303),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_355),
.A2(n_367),
.B1(n_307),
.B2(n_277),
.Y(n_381)
);

INVx13_ASAP7_75t_L g356 ( 
.A(n_311),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_356),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_334),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_304),
.A2(n_269),
.B(n_279),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_358),
.A2(n_371),
.B(n_299),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_325),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_359),
.Y(n_395)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_312),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_362),
.Y(n_397)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_326),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_318),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_368),
.Y(n_376)
);

INVx13_ASAP7_75t_L g364 ( 
.A(n_311),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_364),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_320),
.B(n_284),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_366),
.Y(n_399)
);

OAI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_317),
.A2(n_327),
.B1(n_336),
.B2(n_332),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_318),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_315),
.A2(n_321),
.B(n_324),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_375),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_359),
.A2(n_339),
.B1(n_331),
.B2(n_328),
.Y(n_377)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_377),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_R g380 ( 
.A(n_354),
.B(n_323),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_380),
.B(n_398),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_381),
.A2(n_282),
.B1(n_294),
.B2(n_300),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_342),
.B(n_317),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_382),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_341),
.B(n_321),
.Y(n_383)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_383),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_316),
.C(n_338),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_388),
.B(n_371),
.C(n_370),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_365),
.A2(n_315),
.B1(n_317),
.B2(n_292),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_389),
.A2(n_344),
.B1(n_368),
.B2(n_363),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_350),
.B(n_313),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_390),
.B(n_353),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_369),
.A2(n_292),
.B1(n_322),
.B2(n_306),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_393),
.A2(n_340),
.B1(n_357),
.B2(n_342),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_394),
.B(n_343),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_366),
.Y(n_398)
);

XNOR2x1_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_340),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_401),
.B(n_406),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_347),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_372),
.C(n_374),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_404),
.A2(n_412),
.B1(n_411),
.B2(n_402),
.Y(n_441)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_379),
.Y(n_405)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_405),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_398),
.B(n_353),
.Y(n_407)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_407),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_408),
.B(n_372),
.Y(n_425)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_409),
.Y(n_436)
);

FAx1_ASAP7_75t_SL g410 ( 
.A(n_394),
.B(n_346),
.CI(n_358),
.CON(n_410),
.SN(n_410)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_411),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_382),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_382),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_418),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_392),
.A2(n_360),
.B(n_362),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_413),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_SL g414 ( 
.A1(n_395),
.A2(n_262),
.B1(n_352),
.B2(n_351),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_414),
.A2(n_386),
.B(n_379),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_375),
.B(n_348),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_392),
.A2(n_361),
.B(n_345),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_419),
.B(n_420),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_395),
.B(n_306),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_421),
.B(n_399),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_422),
.A2(n_384),
.B1(n_389),
.B2(n_399),
.Y(n_429)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_423),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_425),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_440),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_429),
.A2(n_441),
.B1(n_420),
.B2(n_413),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_408),
.B(n_384),
.C(n_397),
.Y(n_434)
);

MAJx2_ASAP7_75t_L g446 ( 
.A(n_434),
.B(n_437),
.C(n_438),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_417),
.A2(n_386),
.B(n_376),
.Y(n_435)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_435),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_403),
.B(n_397),
.C(n_393),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_406),
.B(n_381),
.C(n_378),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_401),
.B(n_378),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_436),
.Y(n_442)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_442),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_445),
.A2(n_453),
.B1(n_448),
.B2(n_456),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_432),
.B(n_416),
.Y(n_447)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_447),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_SL g448 ( 
.A(n_428),
.B(n_407),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_448),
.A2(n_453),
.B(n_439),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_433),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_451),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_SL g450 ( 
.A1(n_431),
.A2(n_405),
.B1(n_415),
.B2(n_400),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_450),
.A2(n_430),
.B1(n_402),
.B2(n_438),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_396),
.Y(n_451)
);

OA21x2_ASAP7_75t_SL g452 ( 
.A1(n_424),
.A2(n_417),
.B(n_410),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_452),
.A2(n_447),
.B(n_444),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_441),
.A2(n_419),
.B(n_430),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_434),
.B(n_410),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_454),
.B(n_437),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_459),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_455),
.A2(n_433),
.B1(n_404),
.B2(n_440),
.Y(n_458)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_458),
.Y(n_472)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_460),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_442),
.B(n_385),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_466),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_425),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_443),
.C(n_446),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_465),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_451),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_468),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_463),
.A2(n_439),
.B(n_396),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_473),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_468),
.A2(n_446),
.B(n_373),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_474),
.B(n_475),
.Y(n_482)
);

OA21x2_ASAP7_75t_SL g478 ( 
.A1(n_470),
.A2(n_467),
.B(n_459),
.Y(n_478)
);

A2O1A1Ixp33_ASAP7_75t_L g484 ( 
.A1(n_478),
.A2(n_474),
.B(n_477),
.C(n_473),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_476),
.A2(n_458),
.B1(n_465),
.B2(n_461),
.Y(n_480)
);

AOI322xp5_ASAP7_75t_L g486 ( 
.A1(n_480),
.A2(n_469),
.A3(n_391),
.B1(n_364),
.B2(n_356),
.C1(n_475),
.C2(n_349),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_471),
.B(n_387),
.Y(n_481)
);

AOI21xp33_ASAP7_75t_L g485 ( 
.A1(n_481),
.A2(n_373),
.B(n_391),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_387),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_483),
.B(n_469),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_484),
.A2(n_485),
.B(n_481),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_486),
.B(n_487),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_488),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_490),
.B(n_489),
.Y(n_491)
);

AOI322xp5_ASAP7_75t_L g492 ( 
.A1(n_491),
.A2(n_479),
.A3(n_482),
.B1(n_364),
.B2(n_356),
.C1(n_349),
.C2(n_300),
.Y(n_492)
);

BUFx24_ASAP7_75t_SL g493 ( 
.A(n_492),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_493),
.A2(n_443),
.B1(n_464),
.B2(n_267),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_494),
.A2(n_281),
.B(n_267),
.Y(n_495)
);


endmodule