module real_aes_164_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_755;
wire n_656;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_0), .B(n_121), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_1), .A2(n_130), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_2), .B(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_3), .B(n_137), .Y(n_200) );
INVx1_ASAP7_75t_L g128 ( .A(n_4), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_5), .B(n_137), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_6), .B(n_141), .Y(n_470) );
INVx1_ASAP7_75t_L g504 ( .A(n_7), .Y(n_504) );
OAI22xp5_ASAP7_75t_SL g804 ( .A1(n_8), .A2(n_805), .B1(n_808), .B2(n_809), .Y(n_804) );
INVx1_ASAP7_75t_L g808 ( .A(n_8), .Y(n_808) );
CKINVDCx16_ASAP7_75t_R g821 ( .A(n_9), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_10), .Y(n_542) );
NAND2xp33_ASAP7_75t_L g138 ( .A(n_11), .B(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g118 ( .A(n_12), .Y(n_118) );
AOI221x1_ASAP7_75t_L g216 ( .A1(n_13), .A2(n_25), .B1(n_121), .B2(n_130), .C(n_217), .Y(n_216) );
CKINVDCx16_ASAP7_75t_R g435 ( .A(n_14), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g120 ( .A(n_15), .B(n_121), .Y(n_120) );
AO21x2_ASAP7_75t_L g115 ( .A1(n_16), .A2(n_116), .B(n_119), .Y(n_115) );
INVx1_ASAP7_75t_L g479 ( .A(n_17), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_18), .B(n_155), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_19), .B(n_137), .Y(n_164) );
AO21x1_ASAP7_75t_L g195 ( .A1(n_20), .A2(n_121), .B(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g438 ( .A(n_21), .Y(n_438) );
INVx1_ASAP7_75t_L g477 ( .A(n_22), .Y(n_477) );
INVx1_ASAP7_75t_SL g487 ( .A(n_23), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_24), .B(n_122), .Y(n_570) );
NAND2x1_ASAP7_75t_L g186 ( .A(n_26), .B(n_137), .Y(n_186) );
AOI33xp33_ASAP7_75t_L g516 ( .A1(n_27), .A2(n_54), .A3(n_454), .B1(n_459), .B2(n_517), .B3(n_518), .Y(n_516) );
NAND2x1_ASAP7_75t_L g174 ( .A(n_28), .B(n_139), .Y(n_174) );
INVx1_ASAP7_75t_L g536 ( .A(n_29), .Y(n_536) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_30), .A2(n_89), .B(n_118), .Y(n_117) );
OR2x2_ASAP7_75t_L g142 ( .A(n_30), .B(n_89), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_31), .B(n_462), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_32), .B(n_139), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_33), .B(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_34), .B(n_139), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_35), .A2(n_130), .B(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g127 ( .A(n_36), .B(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g131 ( .A(n_36), .B(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g453 ( .A(n_36), .Y(n_453) );
OR2x6_ASAP7_75t_L g436 ( .A(n_37), .B(n_437), .Y(n_436) );
NOR3xp33_ASAP7_75t_L g819 ( .A(n_37), .B(n_435), .C(n_820), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_38), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_39), .B(n_121), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_40), .B(n_462), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_41), .A2(n_141), .B1(n_148), .B2(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_42), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_43), .B(n_122), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_44), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_45), .B(n_139), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_46), .A2(n_777), .B1(n_778), .B2(n_779), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_46), .Y(n_777) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_47), .B(n_116), .Y(n_506) );
XNOR2xp5_ASAP7_75t_SL g800 ( .A(n_47), .B(n_801), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_48), .B(n_122), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_49), .A2(n_130), .B(n_173), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_50), .Y(n_567) );
XOR2xp5_ASAP7_75t_L g779 ( .A(n_51), .B(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_52), .B(n_139), .Y(n_187) );
AOI22xp33_ASAP7_75t_SL g783 ( .A1(n_53), .A2(n_776), .B1(n_784), .B2(n_786), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_55), .B(n_122), .Y(n_528) );
INVx1_ASAP7_75t_L g124 ( .A(n_56), .Y(n_124) );
INVx1_ASAP7_75t_L g134 ( .A(n_56), .Y(n_134) );
AND2x2_ASAP7_75t_L g529 ( .A(n_57), .B(n_155), .Y(n_529) );
AOI221xp5_ASAP7_75t_L g502 ( .A1(n_58), .A2(n_75), .B1(n_451), .B2(n_462), .C(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_59), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_60), .B(n_137), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_61), .B(n_148), .Y(n_544) );
AOI21xp5_ASAP7_75t_SL g450 ( .A1(n_62), .A2(n_451), .B(n_456), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_63), .A2(n_130), .B(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g473 ( .A(n_64), .Y(n_473) );
AO21x1_ASAP7_75t_L g197 ( .A1(n_65), .A2(n_130), .B(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_66), .B(n_121), .Y(n_150) );
INVx1_ASAP7_75t_L g527 ( .A(n_67), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_68), .B(n_121), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_69), .A2(n_451), .B(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g210 ( .A(n_70), .B(n_156), .Y(n_210) );
INVx1_ASAP7_75t_L g126 ( .A(n_71), .Y(n_126) );
INVx1_ASAP7_75t_L g132 ( .A(n_71), .Y(n_132) );
AND2x2_ASAP7_75t_L g178 ( .A(n_72), .B(n_147), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_73), .B(n_462), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_74), .B(n_796), .Y(n_795) );
OAI22xp5_ASAP7_75t_SL g805 ( .A1(n_76), .A2(n_87), .B1(n_806), .B2(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_76), .Y(n_806) );
AND2x2_ASAP7_75t_L g489 ( .A(n_77), .B(n_147), .Y(n_489) );
INVx1_ASAP7_75t_L g474 ( .A(n_78), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_79), .A2(n_451), .B(n_486), .Y(n_485) );
INVxp33_ASAP7_75t_L g823 ( .A(n_80), .Y(n_823) );
A2O1A1Ixp33_ASAP7_75t_L g568 ( .A1(n_81), .A2(n_451), .B(n_511), .C(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g439 ( .A(n_82), .Y(n_439) );
AND2x2_ASAP7_75t_L g146 ( .A(n_83), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_84), .B(n_121), .Y(n_166) );
AND2x2_ASAP7_75t_SL g448 ( .A(n_85), .B(n_147), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_86), .A2(n_451), .B1(n_514), .B2(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g807 ( .A(n_87), .Y(n_807) );
AND2x2_ASAP7_75t_L g196 ( .A(n_88), .B(n_141), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_90), .B(n_139), .Y(n_165) );
AND2x2_ASAP7_75t_L g190 ( .A(n_91), .B(n_147), .Y(n_190) );
INVx1_ASAP7_75t_L g457 ( .A(n_92), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_93), .B(n_137), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_94), .A2(n_130), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_95), .B(n_139), .Y(n_218) );
AND2x2_ASAP7_75t_L g520 ( .A(n_96), .B(n_147), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_97), .A2(n_98), .B1(n_781), .B2(n_782), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_97), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_98), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_99), .B(n_137), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_100), .A2(n_534), .B(n_535), .C(n_537), .Y(n_533) );
BUFx2_ASAP7_75t_L g794 ( .A(n_101), .Y(n_794) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_102), .A2(n_130), .B(n_135), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_103), .B(n_122), .Y(n_460) );
AOI21xp33_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_813), .B(n_822), .Y(n_104) );
OA22x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_790), .B1(n_794), .B2(n_799), .Y(n_105) );
OAI21xp5_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_776), .B(n_783), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OAI22xp5_ASAP7_75t_SL g108 ( .A1(n_109), .A2(n_431), .B1(n_440), .B2(n_774), .Y(n_108) );
INVx2_ASAP7_75t_L g785 ( .A(n_109), .Y(n_785) );
OAI22x1_ASAP7_75t_SL g801 ( .A1(n_109), .A2(n_802), .B1(n_803), .B2(n_804), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_109), .Y(n_802) );
AND2x4_ASAP7_75t_L g109 ( .A(n_110), .B(n_352), .Y(n_109) );
NOR3xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_264), .C(n_304), .Y(n_110) );
OAI221xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_179), .B1(n_228), .B2(n_243), .C(n_246), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_143), .Y(n_113) );
INVx2_ASAP7_75t_L g261 ( .A(n_114), .Y(n_261) );
AND2x2_ASAP7_75t_L g291 ( .A(n_114), .B(n_292), .Y(n_291) );
BUFx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g229 ( .A(n_115), .B(n_230), .Y(n_229) );
OR2x2_ASAP7_75t_L g236 ( .A(n_115), .B(n_169), .Y(n_236) );
INVx2_ASAP7_75t_L g242 ( .A(n_115), .Y(n_242) );
AND2x2_ASAP7_75t_L g251 ( .A(n_115), .B(n_145), .Y(n_251) );
INVx1_ASAP7_75t_L g267 ( .A(n_115), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_115), .B(n_313), .Y(n_312) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_116), .A2(n_502), .B(n_506), .Y(n_501) );
INVx2_ASAP7_75t_SL g511 ( .A(n_116), .Y(n_511) );
BUFx4f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx3_ASAP7_75t_L g148 ( .A(n_117), .Y(n_148) );
AND2x4_ASAP7_75t_L g141 ( .A(n_118), .B(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_SL g156 ( .A(n_118), .B(n_142), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_129), .B(n_141), .Y(n_119) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_127), .Y(n_121) );
INVx1_ASAP7_75t_L g475 ( .A(n_122), .Y(n_475) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_125), .Y(n_122) );
AND2x6_ASAP7_75t_L g139 ( .A(n_123), .B(n_132), .Y(n_139) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x4_ASAP7_75t_L g137 ( .A(n_125), .B(n_134), .Y(n_137) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx5_ASAP7_75t_L g140 ( .A(n_127), .Y(n_140) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_127), .Y(n_537) );
AND2x2_ASAP7_75t_L g133 ( .A(n_128), .B(n_134), .Y(n_133) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_128), .Y(n_464) );
AND2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
BUFx3_ASAP7_75t_L g465 ( .A(n_131), .Y(n_465) );
INVx2_ASAP7_75t_L g455 ( .A(n_132), .Y(n_455) );
AND2x4_ASAP7_75t_L g451 ( .A(n_133), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g459 ( .A(n_134), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_138), .B(n_140), .Y(n_135) );
INVxp67_ASAP7_75t_L g480 ( .A(n_137), .Y(n_480) );
INVxp67_ASAP7_75t_L g478 ( .A(n_139), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_140), .A2(n_153), .B(n_154), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_140), .A2(n_164), .B(n_165), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_140), .A2(n_174), .B(n_175), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_140), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_140), .A2(n_199), .B(n_200), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_140), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_140), .A2(n_218), .B(n_219), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g456 ( .A1(n_140), .A2(n_457), .B(n_458), .C(n_460), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_140), .B(n_141), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_SL g486 ( .A1(n_140), .A2(n_458), .B(n_487), .C(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_SL g503 ( .A1(n_140), .A2(n_458), .B(n_504), .C(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g514 ( .A(n_140), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_140), .A2(n_458), .B(n_527), .C(n_528), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_140), .A2(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_SL g160 ( .A(n_141), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_141), .B(n_202), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_141), .A2(n_450), .B(n_461), .Y(n_449) );
AND2x2_ASAP7_75t_SL g143 ( .A(n_144), .B(n_157), .Y(n_143) );
INVx4_ASAP7_75t_L g232 ( .A(n_144), .Y(n_232) );
AND2x2_ASAP7_75t_L g263 ( .A(n_144), .B(n_170), .Y(n_263) );
AND2x2_ASAP7_75t_L g339 ( .A(n_144), .B(n_313), .Y(n_339) );
NAND2x1p5_ASAP7_75t_L g381 ( .A(n_144), .B(n_169), .Y(n_381) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_145), .B(n_169), .Y(n_268) );
AND2x2_ASAP7_75t_L g292 ( .A(n_145), .B(n_170), .Y(n_292) );
BUFx2_ASAP7_75t_L g308 ( .A(n_145), .Y(n_308) );
NOR2x1_ASAP7_75t_SL g411 ( .A(n_145), .B(n_313), .Y(n_411) );
OR2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_149), .Y(n_145) );
INVx3_ASAP7_75t_L g189 ( .A(n_147), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_147), .A2(n_189), .B1(n_533), .B2(n_538), .Y(n_532) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_148), .B(n_541), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_155), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_155), .Y(n_177) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_155), .A2(n_216), .B(n_220), .Y(n_215) );
OA21x2_ASAP7_75t_L g278 ( .A1(n_155), .A2(n_216), .B(n_220), .Y(n_278) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g288 ( .A(n_157), .Y(n_288) );
AOI221xp5_ASAP7_75t_L g354 ( .A1(n_157), .A2(n_355), .B1(n_357), .B2(n_359), .C(n_364), .Y(n_354) );
AND2x2_ASAP7_75t_L g374 ( .A(n_157), .B(n_267), .Y(n_374) );
AND2x4_ASAP7_75t_L g157 ( .A(n_158), .B(n_169), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g230 ( .A(n_159), .Y(n_230) );
INVx1_ASAP7_75t_L g283 ( .A(n_159), .Y(n_283) );
AO21x2_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_167), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_160), .B(n_168), .Y(n_167) );
AO21x2_ASAP7_75t_L g313 ( .A1(n_160), .A2(n_161), .B(n_167), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_166), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_169), .B(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g252 ( .A(n_169), .B(n_240), .Y(n_252) );
INVx2_ASAP7_75t_L g294 ( .A(n_169), .Y(n_294) );
AND2x2_ASAP7_75t_L g427 ( .A(n_169), .B(n_242), .Y(n_427) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_170), .Y(n_284) );
AO21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_177), .B(n_178), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_176), .Y(n_171) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_177), .A2(n_483), .B(n_489), .Y(n_482) );
NOR3xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_211), .C(n_226), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_191), .Y(n_180) );
INVx2_ASAP7_75t_L g341 ( .A(n_181), .Y(n_341) );
AND2x2_ASAP7_75t_L g386 ( .A(n_181), .B(n_263), .Y(n_386) );
BUFx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g331 ( .A(n_182), .Y(n_331) );
AND2x4_ASAP7_75t_SL g346 ( .A(n_182), .B(n_258), .Y(n_346) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_189), .B(n_190), .Y(n_182) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_183), .A2(n_189), .B(n_190), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_188), .Y(n_183) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_189), .A2(n_204), .B(n_210), .Y(n_203) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_189), .A2(n_204), .B(n_210), .Y(n_223) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_189), .A2(n_523), .B(n_529), .Y(n_522) );
AO21x2_ASAP7_75t_L g552 ( .A1(n_189), .A2(n_523), .B(n_529), .Y(n_552) );
INVx2_ASAP7_75t_L g300 ( .A(n_191), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_191), .B(n_330), .Y(n_356) );
AND2x4_ASAP7_75t_L g389 ( .A(n_191), .B(n_336), .Y(n_389) );
AND2x4_ASAP7_75t_L g191 ( .A(n_192), .B(n_203), .Y(n_191) );
AND2x2_ASAP7_75t_L g227 ( .A(n_192), .B(n_222), .Y(n_227) );
OR2x2_ASAP7_75t_L g257 ( .A(n_192), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_SL g326 ( .A(n_192), .B(n_278), .Y(n_326) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
BUFx2_ASAP7_75t_L g271 ( .A(n_193), .Y(n_271) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g245 ( .A(n_194), .Y(n_245) );
OAI21x1_ASAP7_75t_SL g194 ( .A1(n_195), .A2(n_197), .B(n_201), .Y(n_194) );
INVx1_ASAP7_75t_L g202 ( .A(n_196), .Y(n_202) );
INVx2_ASAP7_75t_L g258 ( .A(n_203), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_205), .B(n_209), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_211), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_221), .Y(n_212) );
AND2x2_ASAP7_75t_L g226 ( .A(n_213), .B(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g299 ( .A(n_213), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g384 ( .A(n_213), .Y(n_384) );
BUFx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x4_ASAP7_75t_L g244 ( .A(n_214), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g363 ( .A(n_214), .B(n_223), .Y(n_363) );
AND2x2_ASAP7_75t_L g367 ( .A(n_214), .B(n_233), .Y(n_367) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g336 ( .A(n_215), .Y(n_336) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_215), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_221), .B(n_244), .Y(n_320) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_224), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_222), .B(n_245), .Y(n_430) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g234 ( .A(n_223), .B(n_225), .Y(n_234) );
AND2x2_ASAP7_75t_L g316 ( .A(n_223), .B(n_278), .Y(n_316) );
AND2x2_ASAP7_75t_L g335 ( .A(n_223), .B(n_224), .Y(n_335) );
BUFx2_ASAP7_75t_L g256 ( .A(n_224), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_224), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
BUFx3_ASAP7_75t_L g233 ( .A(n_225), .Y(n_233) );
INVxp67_ASAP7_75t_L g276 ( .A(n_225), .Y(n_276) );
INVx1_ASAP7_75t_L g249 ( .A(n_227), .Y(n_249) );
AND2x2_ASAP7_75t_L g285 ( .A(n_227), .B(n_256), .Y(n_285) );
NAND2xp33_ASAP7_75t_L g366 ( .A(n_227), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g403 ( .A(n_227), .B(n_404), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_231), .B1(n_234), .B2(n_235), .C(n_237), .Y(n_228) );
AND2x2_ASAP7_75t_L g332 ( .A(n_229), .B(n_232), .Y(n_332) );
AND2x2_ASAP7_75t_SL g351 ( .A(n_229), .B(n_292), .Y(n_351) );
AND2x2_ASAP7_75t_L g369 ( .A(n_229), .B(n_294), .Y(n_369) );
AND2x2_ASAP7_75t_L g424 ( .A(n_229), .B(n_263), .Y(n_424) );
INVx1_ASAP7_75t_L g240 ( .A(n_230), .Y(n_240) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_230), .Y(n_296) );
CKINVDCx16_ASAP7_75t_R g376 ( .A(n_231), .Y(n_376) );
AND2x4_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_232), .B(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_232), .B(n_283), .Y(n_358) );
AND2x2_ASAP7_75t_L g325 ( .A(n_233), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g361 ( .A(n_233), .Y(n_361) );
AND2x2_ASAP7_75t_L g270 ( .A(n_234), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_234), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g412 ( .A(n_234), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_234), .B(n_336), .Y(n_422) );
AND2x4_ASAP7_75t_L g338 ( .A(n_235), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g409 ( .A(n_236), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_241), .Y(n_238) );
OR2x2_ASAP7_75t_L g280 ( .A(n_241), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g287 ( .A(n_242), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g318 ( .A(n_242), .B(n_292), .Y(n_318) );
AND2x2_ASAP7_75t_L g392 ( .A(n_242), .B(n_313), .Y(n_392) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g340 ( .A(n_244), .B(n_341), .Y(n_340) );
OAI32xp33_ASAP7_75t_L g405 ( .A1(n_244), .A2(n_406), .A3(n_408), .B1(n_409), .B2(n_412), .Y(n_405) );
AND2x4_ASAP7_75t_L g277 ( .A(n_245), .B(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g375 ( .A(n_245), .B(n_278), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_250), .B1(n_253), .B2(n_259), .Y(n_246) );
INVxp67_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_SL g364 ( .A1(n_248), .A2(n_262), .B(n_365), .C(n_366), .Y(n_364) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g348 ( .A(n_249), .B(n_276), .Y(n_348) );
INVx1_ASAP7_75t_SL g419 ( .A(n_250), .Y(n_419) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AND2x4_ASAP7_75t_L g322 ( .A(n_252), .B(n_261), .Y(n_322) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_252), .A2(n_401), .B1(n_402), .B2(n_403), .C(n_405), .Y(n_400) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_257), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OAI22xp33_ASAP7_75t_L g342 ( .A1(n_260), .A2(n_290), .B1(n_343), .B2(n_344), .Y(n_342) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
OAI211xp5_ASAP7_75t_SL g378 ( .A1(n_261), .A2(n_379), .B(n_387), .C(n_400), .Y(n_378) );
INVx2_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g298 ( .A(n_263), .B(n_267), .Y(n_298) );
OAI211xp5_ASAP7_75t_SL g264 ( .A1(n_265), .A2(n_269), .B(n_272), .C(n_301), .Y(n_264) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g295 ( .A(n_267), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g415 ( .A(n_267), .B(n_411), .Y(n_415) );
OAI32xp33_ASAP7_75t_L g372 ( .A1(n_268), .A2(n_373), .A3(n_375), .B1(n_376), .B2(n_377), .Y(n_372) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_SL g362 ( .A(n_271), .B(n_363), .Y(n_362) );
AOI221xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_279), .B1(n_285), .B2(n_286), .C(n_289), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g429 ( .A(n_276), .B(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_277), .B(n_341), .Y(n_343) );
A2O1A1O1Ixp25_ASAP7_75t_L g414 ( .A1(n_277), .A2(n_346), .B(n_362), .C(n_408), .D(n_415), .Y(n_414) );
AOI31xp33_ASAP7_75t_L g416 ( .A1(n_277), .A2(n_298), .A3(n_408), .B(n_415), .Y(n_416) );
AND2x2_ASAP7_75t_L g330 ( .A(n_278), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_280), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx2_ASAP7_75t_L g407 ( .A(n_282), .Y(n_407) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g402 ( .A(n_283), .B(n_294), .Y(n_402) );
INVx1_ASAP7_75t_L g317 ( .A(n_285), .Y(n_317) );
AND2x2_ASAP7_75t_L g302 ( .A(n_286), .B(n_303), .Y(n_302) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
AOI31xp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_293), .A3(n_297), .B(n_299), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_292), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g425 ( .A(n_292), .B(n_371), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x2_ASAP7_75t_L g370 ( .A(n_294), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g396 ( .A(n_294), .Y(n_396) );
INVxp67_ASAP7_75t_L g365 ( .A(n_295), .Y(n_365) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g303 ( .A(n_299), .Y(n_303) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND3xp33_ASAP7_75t_SL g304 ( .A(n_305), .B(n_321), .C(n_337), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_314), .B1(n_318), .B2(n_319), .Y(n_305) );
INVxp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx2_ASAP7_75t_L g391 ( .A(n_308), .Y(n_391) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_312), .Y(n_371) );
INVxp67_ASAP7_75t_SL g397 ( .A(n_312), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_312), .B(n_381), .Y(n_398) );
NAND2xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx1_ASAP7_75t_L g349 ( .A(n_316), .Y(n_349) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_323), .B1(n_332), .B2(n_333), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_324), .B(n_327), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_330), .A2(n_335), .B1(n_369), .B2(n_370), .C(n_372), .Y(n_368) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2x1_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g408 ( .A(n_335), .Y(n_408) );
AND2x2_ASAP7_75t_L g345 ( .A(n_336), .B(n_346), .Y(n_345) );
O2A1O1Ixp33_ASAP7_75t_SL g393 ( .A1(n_336), .A2(n_394), .B(n_398), .C(n_399), .Y(n_393) );
AOI211xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .B(n_342), .C(n_347), .Y(n_337) );
AND2x2_ASAP7_75t_L g388 ( .A(n_341), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g399 ( .A(n_346), .Y(n_399) );
AOI21xp33_ASAP7_75t_SL g347 ( .A1(n_348), .A2(n_349), .B(n_350), .Y(n_347) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
NOR3xp33_ASAP7_75t_L g352 ( .A(n_353), .B(n_378), .C(n_413), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_354), .B(n_368), .Y(n_353) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_L g377 ( .A(n_362), .Y(n_377) );
INVxp67_ASAP7_75t_L g401 ( .A(n_366), .Y(n_401) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g385 ( .A(n_375), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_382), .B1(n_385), .B2(n_386), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .B(n_393), .Y(n_387) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g426 ( .A(n_411), .B(n_427), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .B1(n_417), .B2(n_420), .C(n_423), .Y(n_413) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI31xp33_ASAP7_75t_SL g423 ( .A1(n_424), .A2(n_425), .A3(n_426), .B(n_428), .Y(n_423) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx4_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVx3_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g784 ( .A1(n_433), .A2(n_441), .B1(n_774), .B2(n_785), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_434), .Y(n_433) );
AND2x6_ASAP7_75t_SL g434 ( .A(n_435), .B(n_436), .Y(n_434) );
OR2x6_ASAP7_75t_SL g774 ( .A(n_435), .B(n_775), .Y(n_774) );
OR2x2_ASAP7_75t_L g789 ( .A(n_435), .B(n_436), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_435), .B(n_775), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g775 ( .A(n_436), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_438), .B(n_439), .Y(n_818) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND3x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_661), .C(n_738), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_613), .Y(n_442) );
NOR2xp67_ASAP7_75t_L g443 ( .A(n_444), .B(n_553), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_490), .B1(n_497), .B2(n_546), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_466), .Y(n_445) );
NOR2xp67_ASAP7_75t_SL g596 ( .A(n_446), .B(n_597), .Y(n_596) );
AND2x4_ASAP7_75t_L g611 ( .A(n_446), .B(n_612), .Y(n_611) );
NOR2x1_ASAP7_75t_L g628 ( .A(n_446), .B(n_629), .Y(n_628) );
AND2x4_ASAP7_75t_SL g668 ( .A(n_446), .B(n_669), .Y(n_668) );
INVx4_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_447), .B(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_447), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g603 ( .A(n_447), .Y(n_603) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_447), .Y(n_608) );
AND2x2_ASAP7_75t_L g637 ( .A(n_447), .B(n_577), .Y(n_637) );
OR2x2_ASAP7_75t_L g641 ( .A(n_447), .B(n_482), .Y(n_641) );
AND2x4_ASAP7_75t_L g654 ( .A(n_447), .B(n_612), .Y(n_654) );
NOR2x1_ASAP7_75t_SL g656 ( .A(n_447), .B(n_469), .Y(n_656) );
AND2x2_ASAP7_75t_L g684 ( .A(n_447), .B(n_562), .Y(n_684) );
OR2x6_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
INVxp67_ASAP7_75t_L g543 ( .A(n_451), .Y(n_543) );
NOR2x1p5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVx1_ASAP7_75t_L g518 ( .A(n_454), .Y(n_518) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x6_ASAP7_75t_L g458 ( .A(n_455), .B(n_459), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_458), .A2(n_473), .B1(n_474), .B2(n_475), .Y(n_472) );
INVxp67_ASAP7_75t_L g534 ( .A(n_458), .Y(n_534) );
INVx2_ASAP7_75t_L g572 ( .A(n_458), .Y(n_572) );
AND2x2_ASAP7_75t_L g463 ( .A(n_459), .B(n_464), .Y(n_463) );
INVxp33_ASAP7_75t_L g517 ( .A(n_459), .Y(n_517) );
INVx1_ASAP7_75t_L g545 ( .A(n_462), .Y(n_545) );
AND2x4_ASAP7_75t_L g462 ( .A(n_463), .B(n_465), .Y(n_462) );
INVx1_ASAP7_75t_L g565 ( .A(n_463), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_465), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_466), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_467), .A2(n_742), .B1(n_744), .B2(n_747), .Y(n_741) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_482), .Y(n_467) );
INVx1_ASAP7_75t_L g496 ( .A(n_468), .Y(n_496) );
AND2x2_ASAP7_75t_L g599 ( .A(n_468), .B(n_600), .Y(n_599) );
AND2x4_ASAP7_75t_L g604 ( .A(n_468), .B(n_562), .Y(n_604) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g561 ( .A(n_469), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g577 ( .A(n_469), .Y(n_577) );
AND2x2_ASAP7_75t_L g610 ( .A(n_469), .B(n_482), .Y(n_610) );
AND2x4_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_476), .B(n_481), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_475), .B(n_536), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B1(n_479), .B2(n_480), .Y(n_476) );
INVx2_ASAP7_75t_L g494 ( .A(n_482), .Y(n_494) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_482), .Y(n_579) );
INVx1_ASAP7_75t_L g598 ( .A(n_482), .Y(n_598) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_482), .Y(n_667) );
INVx1_ASAP7_75t_L g679 ( .A(n_482), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OAI31xp33_ASAP7_75t_SL g733 ( .A1(n_491), .A2(n_734), .A3(n_735), .B(n_736), .Y(n_733) );
NOR2x1_ASAP7_75t_L g491 ( .A(n_492), .B(n_495), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g658 ( .A(n_493), .B(n_560), .Y(n_658) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g574 ( .A(n_494), .Y(n_574) );
AND2x4_ASAP7_75t_SL g694 ( .A(n_496), .B(n_598), .Y(n_694) );
OAI21xp5_ASAP7_75t_L g614 ( .A1(n_497), .A2(n_615), .B(n_618), .Y(n_614) );
OR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_507), .Y(n_497) );
INVx2_ASAP7_75t_L g587 ( .A(n_498), .Y(n_587) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2x1p5_ASAP7_75t_L g714 ( .A(n_499), .B(n_622), .Y(n_714) );
BUFx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g624 ( .A(n_500), .B(n_530), .Y(n_624) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVxp67_ASAP7_75t_L g549 ( .A(n_501), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_501), .B(n_510), .Y(n_584) );
AND2x4_ASAP7_75t_L g594 ( .A(n_501), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g639 ( .A(n_501), .B(n_531), .Y(n_639) );
INVx2_ASAP7_75t_L g647 ( .A(n_501), .Y(n_647) );
INVx1_ASAP7_75t_L g746 ( .A(n_501), .Y(n_746) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_501), .Y(n_755) );
INVx1_ASAP7_75t_L g692 ( .A(n_507), .Y(n_692) );
NAND2x1p5_ASAP7_75t_L g507 ( .A(n_508), .B(n_521), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g548 ( .A(n_509), .B(n_549), .Y(n_548) );
AND2x4_ASAP7_75t_L g687 ( .A(n_509), .B(n_622), .Y(n_687) );
AND2x2_ASAP7_75t_L g704 ( .A(n_509), .B(n_522), .Y(n_704) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_510), .B(n_552), .Y(n_727) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_520), .Y(n_510) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_511), .A2(n_512), .B(n_520), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_513), .B(n_519), .Y(n_512) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g650 ( .A(n_521), .B(n_548), .Y(n_650) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_530), .Y(n_521) );
INVx2_ASAP7_75t_L g556 ( .A(n_522), .Y(n_556) );
NOR2xp67_ASAP7_75t_L g737 ( .A(n_522), .B(n_530), .Y(n_737) );
NOR2x1_ASAP7_75t_L g745 ( .A(n_522), .B(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
AND2x2_ASAP7_75t_L g653 ( .A(n_530), .B(n_557), .Y(n_653) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_531), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g582 ( .A(n_531), .Y(n_582) );
AND2x4_ASAP7_75t_L g646 ( .A(n_531), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g676 ( .A(n_531), .Y(n_676) );
OR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_539), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_539) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_547), .A2(n_560), .B1(n_698), .B2(n_699), .C(n_700), .Y(n_697) );
NAND2x1p5_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
AND2x2_ASAP7_75t_L g674 ( .A(n_548), .B(n_675), .Y(n_674) );
BUFx2_ASAP7_75t_L g717 ( .A(n_548), .Y(n_717) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g660 ( .A(n_551), .B(n_584), .Y(n_660) );
INVx3_ASAP7_75t_L g622 ( .A(n_552), .Y(n_622) );
AND2x2_ASAP7_75t_L g754 ( .A(n_552), .B(n_755), .Y(n_754) );
NAND3xp33_ASAP7_75t_SL g553 ( .A(n_554), .B(n_585), .C(n_601), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_558), .B1(n_575), .B2(n_580), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_555), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g685 ( .A(n_555), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g696 ( .A(n_555), .B(n_591), .Y(n_696) );
AND2x2_ASAP7_75t_L g766 ( .A(n_555), .B(n_639), .Y(n_766) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
INVx2_ASAP7_75t_L g595 ( .A(n_557), .Y(n_595) );
INVx1_ASAP7_75t_L g644 ( .A(n_557), .Y(n_644) );
INVxp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OAI222xp33_ASAP7_75t_L g711 ( .A1(n_559), .A2(n_712), .B1(n_713), .B2(n_715), .C1(n_716), .C2(n_718), .Y(n_711) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_573), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_560), .B(n_587), .Y(n_586) );
NOR2x1_ASAP7_75t_L g719 ( .A(n_560), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g678 ( .A(n_561), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g734 ( .A(n_561), .B(n_608), .Y(n_734) );
INVx2_ASAP7_75t_L g600 ( .A(n_562), .Y(n_600) );
INVx1_ASAP7_75t_L g612 ( .A(n_562), .Y(n_612) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_562), .Y(n_669) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_568), .Y(n_562) );
NOR3xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .C(n_567), .Y(n_564) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_574), .Y(n_617) );
INVx3_ASAP7_75t_L g636 ( .A(n_574), .Y(n_636) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g702 ( .A(n_576), .Y(n_702) );
NAND2x1_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_L g689 ( .A(n_578), .Y(n_689) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
INVx1_ASAP7_75t_L g690 ( .A(n_581), .Y(n_690) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g591 ( .A(n_582), .Y(n_591) );
AND2x2_ASAP7_75t_L g709 ( .A(n_582), .B(n_594), .Y(n_709) );
AND2x2_ASAP7_75t_L g772 ( .A(n_582), .B(n_704), .Y(n_772) );
AND2x2_ASAP7_75t_L g701 ( .A(n_583), .B(n_621), .Y(n_701) );
INVx1_ASAP7_75t_L g712 ( .A(n_583), .Y(n_712) );
AND2x2_ASAP7_75t_L g729 ( .A(n_583), .B(n_676), .Y(n_729) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_588), .B1(n_592), .B2(n_596), .Y(n_585) );
OAI21xp5_ASAP7_75t_L g601 ( .A1(n_588), .A2(n_602), .B(n_605), .Y(n_601) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g633 ( .A(n_591), .B(n_594), .Y(n_633) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x4_ASAP7_75t_L g736 ( .A(n_594), .B(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_L g699 ( .A(n_597), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_598), .Y(n_627) );
AND2x2_ASAP7_75t_SL g607 ( .A(n_599), .B(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g672 ( .A(n_599), .Y(n_672) );
AND2x2_ASAP7_75t_L g770 ( .A(n_599), .B(n_667), .Y(n_770) );
INVx1_ASAP7_75t_L g725 ( .A(n_600), .Y(n_725) );
INVx1_ASAP7_75t_L g631 ( .A(n_602), .Y(n_631) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g720 ( .A(n_603), .Y(n_720) );
INVx4_ASAP7_75t_L g629 ( .A(n_604), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AOI32xp33_ASAP7_75t_L g700 ( .A1(n_607), .A2(n_701), .A3(n_702), .B1(n_703), .B2(n_704), .Y(n_700) );
AND2x2_ASAP7_75t_L g695 ( .A(n_608), .B(n_610), .Y(n_695) );
O2A1O1Ixp33_ASAP7_75t_SL g758 ( .A1(n_608), .A2(n_759), .B(n_760), .C(n_762), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
AND2x2_ASAP7_75t_SL g723 ( .A(n_610), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g762 ( .A(n_610), .Y(n_762) );
AND2x2_ASAP7_75t_L g616 ( .A(n_611), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g743 ( .A(n_611), .Y(n_743) );
AND2x2_ASAP7_75t_L g749 ( .A(n_611), .B(n_636), .Y(n_749) );
NOR3x1_ASAP7_75t_L g613 ( .A(n_614), .B(n_630), .C(n_648), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_625), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
AND2x2_ASAP7_75t_L g638 ( .A(n_621), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g681 ( .A(n_621), .B(n_646), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_621), .B(n_667), .Y(n_708) );
INVx3_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_629), .B(n_636), .Y(n_735) );
INVx2_ASAP7_75t_L g757 ( .A(n_629), .Y(n_757) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B(n_634), .Y(n_630) );
OAI221xp5_ASAP7_75t_L g721 ( .A1(n_631), .A2(n_722), .B1(n_726), .B2(n_728), .C(n_733), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_632), .A2(n_752), .B1(n_753), .B2(n_756), .Y(n_751) );
INVx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_638), .B1(n_640), .B2(n_642), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
AND2x2_ASAP7_75t_L g680 ( .A(n_636), .B(n_656), .Y(n_680) );
INVx1_ASAP7_75t_L g686 ( .A(n_636), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_636), .B(n_654), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_639), .B(n_707), .Y(n_773) );
NAND2x1_ASAP7_75t_L g756 ( .A(n_640), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
NOR2x1_ASAP7_75t_L g671 ( .A(n_641), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
NAND2x1_ASAP7_75t_SL g759 ( .A(n_644), .B(n_646), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_644), .B(n_744), .Y(n_765) );
OR2x2_ASAP7_75t_L g726 ( .A(n_645), .B(n_727), .Y(n_726) );
INVx3_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g761 ( .A(n_646), .B(n_687), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_649), .B(n_655), .Y(n_648) );
OAI21xp33_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_651), .B(n_654), .Y(n_649) );
OR2x2_ASAP7_75t_L g713 ( .A(n_652), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g747 ( .A(n_653), .B(n_745), .Y(n_747) );
AND2x2_ASAP7_75t_SL g693 ( .A(n_654), .B(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g703 ( .A(n_654), .Y(n_703) );
OAI21xp33_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B(n_659), .Y(n_655) );
AND2x2_ASAP7_75t_L g688 ( .A(n_656), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_705), .Y(n_662) );
NOR3xp33_ASAP7_75t_SL g663 ( .A(n_664), .B(n_682), .C(n_697), .Y(n_663) );
A2O1A1Ixp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_670), .B(n_673), .C(n_677), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
BUFx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
BUFx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g731 ( .A(n_676), .Y(n_731) );
AND2x2_ASAP7_75t_L g744 ( .A(n_676), .B(n_745), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .B(n_681), .Y(n_677) );
INVx1_ASAP7_75t_L g752 ( .A(n_678), .Y(n_752) );
OAI21xp5_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_690), .B(n_691), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_685), .B1(n_687), .B2(n_688), .Y(n_683) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_684), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B1(n_695), .B2(n_696), .Y(n_691) );
INVx1_ASAP7_75t_SL g698 ( .A(n_696), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_702), .B(n_743), .Y(n_742) );
OAI22xp33_ASAP7_75t_SL g768 ( .A1(n_703), .A2(n_769), .B1(n_771), .B2(n_773), .Y(n_768) );
AOI211x1_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_710), .B(n_711), .C(n_721), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
OAI21xp5_ASAP7_75t_L g763 ( .A1(n_723), .A2(n_764), .B(n_766), .Y(n_763) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g732 ( .A(n_727), .Y(n_732) );
NOR2xp67_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_730), .B(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NAND4xp25_ASAP7_75t_L g739 ( .A(n_740), .B(n_750), .C(n_763), .D(n_767), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_748), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_758), .Y(n_750) );
INVxp67_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_SL g787 ( .A(n_788), .Y(n_787) );
INVx3_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_795), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
HB1xp67_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
OAI21xp5_ASAP7_75t_L g799 ( .A1(n_795), .A2(n_800), .B(n_810), .Y(n_799) );
INVx1_ASAP7_75t_SL g796 ( .A(n_797), .Y(n_796) );
BUFx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
BUFx2_ASAP7_75t_L g812 ( .A(n_798), .Y(n_812) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g809 ( .A(n_805), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_SL g815 ( .A(n_816), .Y(n_815) );
INVx3_ASAP7_75t_SL g816 ( .A(n_817), .Y(n_816) );
BUFx2_ASAP7_75t_L g824 ( .A(n_817), .Y(n_824) );
AND2x2_ASAP7_75t_SL g817 ( .A(n_818), .B(n_819), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
endmodule