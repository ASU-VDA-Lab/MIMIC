module fake_netlist_6_1017_n_1674 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1674);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1674;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_87),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_92),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_0),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_67),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_21),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_32),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_25),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_76),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_44),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_102),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_6),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_34),
.Y(n_170)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_42),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_104),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_115),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_79),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_29),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_60),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_83),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_64),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_25),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_80),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_133),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_114),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_109),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_113),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_98),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_82),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_23),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_40),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_62),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_58),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_122),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_34),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_112),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_88),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_26),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_42),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_140),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_132),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_61),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_12),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_27),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_33),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_81),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_68),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_55),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_0),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_107),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_50),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_56),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_108),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_48),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_74),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_124),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_116),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_50),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_39),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_21),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_99),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_44),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_145),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_93),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_69),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_106),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_100),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_71),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_46),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_22),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_95),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_131),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_118),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_36),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_77),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_10),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_134),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_4),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_142),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_52),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_121),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_41),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_40),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_49),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_78),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_45),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_137),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_10),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_36),
.Y(n_251)
);

BUFx8_ASAP7_75t_SL g252 ( 
.A(n_52),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_59),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_29),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_17),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_154),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_54),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_33),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_46),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_12),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_48),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_26),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_126),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_11),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_136),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_20),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_54),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_111),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_49),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_19),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_89),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_15),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_63),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_73),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_96),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_147),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_28),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_97),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_8),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_119),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_1),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_139),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_15),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_75),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_51),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_150),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_117),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_23),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_31),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_65),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_53),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_28),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_1),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_31),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_3),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_110),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_146),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_141),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_105),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_135),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_2),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_72),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_123),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_128),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_138),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_195),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_252),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_297),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_2),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_221),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_221),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_225),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_221),
.Y(n_314)
);

NOR2xp67_ASAP7_75t_L g315 ( 
.A(n_166),
.B(n_3),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_221),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_269),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_237),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_155),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_221),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_221),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_156),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_224),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_246),
.B(n_4),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_162),
.B(n_5),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_263),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_224),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_246),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_186),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_L g330 ( 
.A(n_166),
.B(n_5),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_224),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_264),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_292),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_292),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_157),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_161),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_165),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_224),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_168),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_224),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_224),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_281),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_281),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_166),
.B(n_7),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_172),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_160),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_281),
.Y(n_347)
);

BUFx6f_ASAP7_75t_SL g348 ( 
.A(n_160),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_173),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_175),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_176),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_281),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_180),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_264),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_281),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_302),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_184),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_281),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_163),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_163),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_185),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_201),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_196),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_170),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_201),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_170),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_188),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_193),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_158),
.B(n_7),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_198),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_242),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_242),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_199),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_264),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_267),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_267),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_208),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_177),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_177),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_215),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_311),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_356),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_356),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_315),
.B(n_166),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_311),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_356),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_312),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_340),
.B(n_218),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_312),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_314),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_314),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_356),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_316),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_320),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_196),
.Y(n_396)
);

INVx6_ASAP7_75t_L g397 ( 
.A(n_346),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_341),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_320),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_341),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_321),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_321),
.B(n_323),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_323),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_327),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_327),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_331),
.B(n_219),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_331),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_309),
.B(n_212),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_338),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_338),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_342),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_342),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_343),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_317),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_329),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_376),
.B(n_262),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_347),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_325),
.B(n_308),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_347),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_352),
.Y(n_421)
);

NOR2x1_ASAP7_75t_L g422 ( 
.A(n_315),
.B(n_183),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_344),
.B(n_183),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_352),
.Y(n_424)
);

NAND2xp33_ASAP7_75t_SL g425 ( 
.A(n_324),
.B(n_200),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

AND2x6_ASAP7_75t_L g427 ( 
.A(n_355),
.B(n_302),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_358),
.Y(n_428)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_358),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_359),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_359),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_363),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_363),
.B(n_262),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_360),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_360),
.B(n_272),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_344),
.B(n_229),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_378),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_378),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_362),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_362),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_310),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_330),
.B(n_230),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_379),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_334),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_379),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_365),
.B(n_272),
.Y(n_446)
);

AND2x6_ASAP7_75t_L g447 ( 
.A(n_369),
.B(n_302),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_365),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_371),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_388),
.B(n_319),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_388),
.B(n_322),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_386),
.Y(n_452)
);

BUFx10_ASAP7_75t_L g453 ( 
.A(n_419),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_396),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_335),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_419),
.A2(n_380),
.B1(n_361),
.B2(n_367),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_436),
.B(n_336),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_396),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_403),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_337),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_406),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_386),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_417),
.B(n_371),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_403),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_408),
.B(n_345),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_415),
.B(n_351),
.Y(n_466)
);

INVxp33_ASAP7_75t_L g467 ( 
.A(n_441),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_386),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_417),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_408),
.A2(n_333),
.B1(n_301),
.B2(n_200),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_442),
.B(n_353),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_403),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_417),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_386),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_415),
.B(n_357),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_437),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_386),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_406),
.B(n_368),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_387),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_423),
.B(n_370),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_435),
.B(n_446),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_387),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_389),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_389),
.Y(n_484)
);

INVx5_ASAP7_75t_L g485 ( 
.A(n_427),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_435),
.B(n_158),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_423),
.B(n_373),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_386),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_391),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_391),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_423),
.B(n_377),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_425),
.B(n_332),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_386),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_403),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_437),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_386),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_393),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_397),
.B(n_339),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_405),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_405),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_405),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_405),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_438),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_397),
.B(n_349),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_425),
.B(n_332),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_393),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_397),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_423),
.B(n_346),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_438),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_393),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_443),
.Y(n_511)
);

AND2x2_ASAP7_75t_SL g512 ( 
.A(n_423),
.B(n_209),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_397),
.B(n_350),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_416),
.Y(n_514)
);

OAI22xp33_ASAP7_75t_L g515 ( 
.A1(n_432),
.A2(n_328),
.B1(n_374),
.B2(n_354),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_423),
.B(n_217),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_410),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_410),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_410),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_410),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_447),
.B(n_397),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_435),
.B(n_372),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_447),
.B(n_226),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_443),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_445),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_416),
.B(n_307),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_432),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_447),
.A2(n_289),
.B1(n_191),
.B2(n_291),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_445),
.Y(n_529)
);

NAND2xp33_ASAP7_75t_L g530 ( 
.A(n_447),
.B(n_302),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_432),
.B(n_354),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_427),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_433),
.B(n_374),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_433),
.B(n_328),
.Y(n_534)
);

AND3x2_ASAP7_75t_L g535 ( 
.A(n_441),
.B(n_303),
.C(n_241),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_393),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_393),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_433),
.B(n_364),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_392),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_447),
.A2(n_222),
.B1(n_191),
.B2(n_213),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_384),
.B(n_160),
.Y(n_541)
);

AO22x2_ASAP7_75t_L g542 ( 
.A1(n_384),
.A2(n_222),
.B1(n_213),
.B2(n_220),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_393),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_393),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_394),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_384),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_393),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_447),
.A2(n_348),
.B1(n_318),
.B2(n_326),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_444),
.B(n_366),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_418),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_447),
.B(n_227),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_394),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_447),
.B(n_273),
.Y(n_553)
);

AND2x2_ASAP7_75t_SL g554 ( 
.A(n_384),
.B(n_209),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_444),
.Y(n_555)
);

BUFx4f_ASAP7_75t_L g556 ( 
.A(n_447),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_384),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_384),
.B(n_302),
.Y(n_558)
);

BUFx10_ASAP7_75t_L g559 ( 
.A(n_447),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_395),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_399),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_404),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_404),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_399),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_418),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_411),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_418),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_404),
.Y(n_568)
);

NOR2x1p5_ASAP7_75t_L g569 ( 
.A(n_446),
.B(n_171),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_404),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_411),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_446),
.B(n_174),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_422),
.B(n_234),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_422),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_431),
.B(n_306),
.Y(n_575)
);

INVx5_ASAP7_75t_L g576 ( 
.A(n_427),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_418),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_429),
.B(n_348),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_431),
.B(n_220),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_448),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_404),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_429),
.B(n_348),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_429),
.B(n_235),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_448),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_404),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_429),
.B(n_239),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_429),
.B(n_243),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_404),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_412),
.B(n_249),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_414),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_420),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_463),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_461),
.B(n_421),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_463),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_554),
.B(n_302),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_465),
.B(n_453),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_557),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_512),
.B(n_421),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_557),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_459),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_549),
.B(n_159),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_481),
.B(n_313),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_454),
.Y(n_603)
);

NOR2x1p5_ASAP7_75t_L g604 ( 
.A(n_549),
.B(n_164),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_531),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_512),
.B(n_265),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_453),
.B(n_271),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_556),
.B(n_241),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_534),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_556),
.B(n_298),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_507),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_450),
.B(n_448),
.Y(n_612)
);

NOR2xp67_ASAP7_75t_SL g613 ( 
.A(n_485),
.B(n_174),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_542),
.A2(n_244),
.B1(n_245),
.B2(n_236),
.Y(n_614)
);

AND2x6_ASAP7_75t_SL g615 ( 
.A(n_538),
.B(n_232),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_459),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_453),
.B(n_167),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_451),
.B(n_448),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_574),
.B(n_169),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_507),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_514),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_538),
.B(n_182),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_464),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_546),
.Y(n_624)
);

NOR2xp67_ASAP7_75t_L g625 ( 
.A(n_456),
.B(n_274),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_574),
.B(n_192),
.Y(n_626)
);

AO22x2_ASAP7_75t_L g627 ( 
.A1(n_492),
.A2(n_296),
.B1(n_247),
.B2(n_253),
.Y(n_627)
);

AO221x1_ASAP7_75t_L g628 ( 
.A1(n_542),
.A2(n_232),
.B1(n_236),
.B2(n_244),
.C(n_245),
.Y(n_628)
);

O2A1O1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_458),
.A2(n_473),
.B(n_469),
.C(n_481),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_522),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_478),
.B(n_381),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_546),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_522),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_556),
.B(n_298),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_498),
.B(n_278),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_521),
.A2(n_402),
.B(n_383),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_476),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_538),
.B(n_250),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_504),
.B(n_513),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_467),
.B(n_538),
.Y(n_640)
);

AOI221xp5_ASAP7_75t_L g641 ( 
.A1(n_470),
.A2(n_285),
.B1(n_240),
.B2(n_250),
.C(n_254),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_559),
.B(n_305),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_580),
.B(n_381),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_580),
.B(n_381),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_467),
.B(n_264),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_455),
.B(n_205),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_542),
.A2(n_254),
.B1(n_260),
.B2(n_277),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_457),
.B(n_385),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_514),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_559),
.B(n_305),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_460),
.B(n_206),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_471),
.B(n_207),
.Y(n_652)
);

OAI22xp33_ASAP7_75t_L g653 ( 
.A1(n_579),
.A2(n_260),
.B1(n_277),
.B2(n_279),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_508),
.B(n_385),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_584),
.A2(n_280),
.B1(n_282),
.B2(n_284),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_516),
.B(n_385),
.Y(n_656)
);

NOR2xp67_ASAP7_75t_L g657 ( 
.A(n_548),
.B(n_286),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_495),
.B(n_390),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_486),
.B(n_572),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_472),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_503),
.B(n_509),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_511),
.B(n_390),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_569),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_542),
.A2(n_279),
.B1(n_291),
.B2(n_294),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_472),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_524),
.B(n_390),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_480),
.B(n_210),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_494),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_487),
.B(n_211),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_491),
.B(n_290),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_533),
.B(n_216),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_579),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_452),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_466),
.B(n_231),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_559),
.B(n_299),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_525),
.Y(n_676)
);

OAI22xp33_ASAP7_75t_L g677 ( 
.A1(n_579),
.A2(n_294),
.B1(n_178),
.B2(n_253),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_475),
.B(n_527),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_583),
.A2(n_402),
.B(n_382),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_529),
.B(n_401),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_479),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_523),
.B(n_551),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_584),
.B(n_160),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_505),
.B(n_238),
.Y(n_684)
);

INVx8_ASAP7_75t_L g685 ( 
.A(n_486),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_479),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_575),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_553),
.B(n_486),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_494),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_572),
.B(n_204),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_539),
.B(n_401),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_589),
.B(n_248),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_527),
.B(n_251),
.Y(n_693)
);

O2A1O1Ixp5_ASAP7_75t_L g694 ( 
.A1(n_541),
.A2(n_407),
.B(n_428),
.C(n_268),
.Y(n_694)
);

INVx4_ASAP7_75t_L g695 ( 
.A(n_452),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_575),
.B(n_375),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_499),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_482),
.Y(n_698)
);

BUFx6f_ASAP7_75t_SL g699 ( 
.A(n_579),
.Y(n_699)
);

BUFx2_ASAP7_75t_L g700 ( 
.A(n_555),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_482),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_499),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_545),
.B(n_552),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_564),
.B(n_407),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_566),
.B(n_407),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_571),
.B(n_255),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_483),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_586),
.A2(n_194),
.B1(n_179),
.B2(n_181),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_555),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_483),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_526),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_484),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_500),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_515),
.B(n_204),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_484),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_452),
.B(n_430),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_489),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_590),
.B(n_428),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_489),
.B(n_430),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_490),
.B(n_430),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_587),
.A2(n_194),
.B1(n_187),
.B2(n_304),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_490),
.B(n_257),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_578),
.B(n_375),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_573),
.A2(n_190),
.B1(n_187),
.B2(n_304),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_582),
.B(n_258),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_452),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_497),
.B(n_430),
.Y(n_727)
);

AND2x2_ASAP7_75t_SL g728 ( 
.A(n_530),
.B(n_189),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_497),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_497),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_560),
.B(n_259),
.Y(n_731)
);

BUFx4f_ASAP7_75t_L g732 ( 
.A(n_558),
.Y(n_732)
);

OAI221xp5_ASAP7_75t_L g733 ( 
.A1(n_540),
.A2(n_528),
.B1(n_561),
.B2(n_560),
.C(n_202),
.Y(n_733)
);

OAI221xp5_ASAP7_75t_L g734 ( 
.A1(n_561),
.A2(n_197),
.B1(n_203),
.B2(n_214),
.C(n_223),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_497),
.B(n_430),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_462),
.B(n_430),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_500),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_501),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_558),
.A2(n_197),
.B1(n_203),
.B2(n_287),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_L g740 ( 
.A(n_558),
.B(n_214),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_462),
.B(n_434),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_501),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_502),
.Y(n_743)
);

AND2x6_ASAP7_75t_SL g744 ( 
.A(n_535),
.B(n_223),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_468),
.B(n_261),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_468),
.B(n_266),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_468),
.B(n_434),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_474),
.B(n_434),
.Y(n_748)
);

OR2x6_ASAP7_75t_L g749 ( 
.A(n_497),
.B(n_228),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_681),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_686),
.Y(n_751)
);

OAI21xp5_ASAP7_75t_L g752 ( 
.A1(n_682),
.A2(n_530),
.B(n_474),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_673),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_601),
.B(n_693),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_614),
.A2(n_558),
.B1(n_233),
.B2(n_247),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_624),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_600),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_631),
.B(n_493),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_648),
.B(n_493),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_609),
.B(n_493),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_621),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_646),
.B(n_651),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_685),
.Y(n_763)
);

OR2x6_ASAP7_75t_L g764 ( 
.A(n_685),
.B(n_256),
.Y(n_764)
);

OAI321xp33_ASAP7_75t_L g765 ( 
.A1(n_641),
.A2(n_268),
.A3(n_275),
.B1(n_287),
.B2(n_276),
.C(n_449),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_646),
.B(n_543),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_602),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_688),
.A2(n_496),
.B(n_488),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_645),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_652),
.B(n_543),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_682),
.A2(n_544),
.B(n_547),
.Y(n_771)
);

NOR2x1p5_ASAP7_75t_SL g772 ( 
.A(n_616),
.B(n_502),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_652),
.B(n_544),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_624),
.Y(n_774)
);

OA21x2_ASAP7_75t_L g775 ( 
.A1(n_595),
.A2(n_591),
.B(n_577),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_596),
.A2(n_275),
.B(n_276),
.C(n_270),
.Y(n_776)
);

AOI21x1_ASAP7_75t_L g777 ( 
.A1(n_716),
.A2(n_565),
.B(n_520),
.Y(n_777)
);

AOI21x1_ASAP7_75t_L g778 ( 
.A1(n_727),
.A2(n_565),
.B(n_520),
.Y(n_778)
);

O2A1O1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_629),
.A2(n_518),
.B(n_517),
.C(n_577),
.Y(n_779)
);

BUFx12f_ASAP7_75t_L g780 ( 
.A(n_744),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_593),
.B(n_544),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_688),
.A2(n_496),
.B(n_477),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_698),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_612),
.A2(n_496),
.B(n_477),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_618),
.A2(n_488),
.B(n_570),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_703),
.B(n_547),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_703),
.B(n_563),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_692),
.B(n_563),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_595),
.A2(n_598),
.B(n_636),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_701),
.Y(n_790)
);

AOI21x1_ASAP7_75t_L g791 ( 
.A1(n_727),
.A2(n_519),
.B(n_518),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_685),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_596),
.A2(n_568),
.B1(n_563),
.B2(n_581),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_605),
.B(n_283),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_692),
.B(n_568),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_623),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_649),
.B(n_288),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_695),
.A2(n_485),
.B(n_532),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_679),
.A2(n_550),
.B(n_517),
.Y(n_799)
);

INVxp67_ASAP7_75t_SL g800 ( 
.A(n_624),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_707),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_630),
.Y(n_802)
);

NOR3xp33_ASAP7_75t_L g803 ( 
.A(n_617),
.B(n_683),
.C(n_678),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_614),
.A2(n_293),
.B(n_295),
.C(n_567),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_647),
.A2(n_550),
.B(n_567),
.C(n_449),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_639),
.A2(n_568),
.B1(n_581),
.B2(n_510),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_723),
.B(n_581),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_624),
.B(n_506),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_710),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_712),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_715),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_717),
.B(n_506),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_660),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_665),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_654),
.A2(n_485),
.B(n_532),
.Y(n_815)
);

OAI21x1_ASAP7_75t_L g816 ( 
.A1(n_736),
.A2(n_382),
.B(n_383),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_632),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_667),
.B(n_506),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_632),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_668),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_608),
.A2(n_485),
.B(n_532),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_689),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_667),
.B(n_506),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_669),
.B(n_506),
.Y(n_824)
);

AOI21x1_ASAP7_75t_L g825 ( 
.A1(n_735),
.A2(n_382),
.B(n_383),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_642),
.A2(n_650),
.B(n_675),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_617),
.B(n_537),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_632),
.B(n_537),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_632),
.B(n_537),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_669),
.B(n_537),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_700),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_673),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_650),
.A2(n_576),
.B(n_537),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_656),
.A2(n_576),
.B(n_536),
.Y(n_834)
);

AO21x1_ASAP7_75t_L g835 ( 
.A1(n_608),
.A2(n_420),
.B(n_426),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_619),
.B(n_536),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_643),
.B(n_510),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_637),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_659),
.B(n_536),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_697),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_676),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_606),
.A2(n_420),
.B(n_426),
.C(n_424),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_659),
.A2(n_536),
.B1(n_510),
.B2(n_588),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_603),
.Y(n_844)
);

AOI21xp33_ASAP7_75t_L g845 ( 
.A1(n_674),
.A2(n_8),
.B(n_9),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_619),
.B(n_510),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_599),
.B(n_510),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_644),
.B(n_588),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_661),
.B(n_588),
.Y(n_849)
);

AOI21x1_ASAP7_75t_L g850 ( 
.A1(n_735),
.A2(n_382),
.B(n_383),
.Y(n_850)
);

NOR3xp33_ASAP7_75t_L g851 ( 
.A(n_696),
.B(n_439),
.C(n_449),
.Y(n_851)
);

AO21x1_ASAP7_75t_L g852 ( 
.A1(n_610),
.A2(n_424),
.B(n_426),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_626),
.B(n_204),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_626),
.B(n_588),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_599),
.B(n_576),
.Y(n_855)
);

OAI21x1_ASAP7_75t_L g856 ( 
.A1(n_741),
.A2(n_398),
.B(n_424),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_633),
.B(n_204),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_711),
.B(n_585),
.Y(n_858)
);

NAND2x1p5_ASAP7_75t_L g859 ( 
.A(n_732),
.B(n_585),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_610),
.A2(n_398),
.B(n_427),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_611),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_634),
.A2(n_562),
.B(n_585),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_597),
.A2(n_562),
.B1(n_449),
.B2(n_439),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_634),
.A2(n_562),
.B(n_398),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_702),
.Y(n_865)
);

OAI21xp33_ASAP7_75t_L g866 ( 
.A1(n_674),
.A2(n_440),
.B(n_434),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_732),
.A2(n_562),
.B(n_413),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_747),
.A2(n_413),
.B(n_409),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_647),
.B(n_440),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_592),
.B(n_440),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_719),
.A2(n_427),
.B(n_400),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_594),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_709),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_720),
.A2(n_427),
.B(n_400),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_748),
.A2(n_413),
.B(n_409),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_664),
.B(n_440),
.Y(n_876)
);

O2A1O1Ixp5_ASAP7_75t_L g877 ( 
.A1(n_694),
.A2(n_400),
.B(n_427),
.C(n_434),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_722),
.B(n_440),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_640),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_726),
.A2(n_729),
.B(n_730),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_663),
.B(n_9),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_722),
.B(n_440),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_725),
.B(n_440),
.Y(n_883)
);

NOR2x1_ASAP7_75t_L g884 ( 
.A(n_607),
.B(n_400),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_677),
.A2(n_400),
.B(n_13),
.C(n_14),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_677),
.A2(n_11),
.B(n_13),
.C(n_14),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_738),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_611),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_664),
.B(n_440),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_687),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_728),
.B(n_434),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_742),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_728),
.B(n_434),
.Y(n_893)
);

CKINVDCx8_ASAP7_75t_R g894 ( 
.A(n_615),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_684),
.A2(n_746),
.B1(n_745),
.B2(n_657),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_671),
.B(n_16),
.Y(n_896)
);

AOI21xp33_ASAP7_75t_L g897 ( 
.A1(n_684),
.A2(n_16),
.B(n_17),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_726),
.A2(n_413),
.B(n_409),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_611),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_671),
.B(n_18),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_713),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_737),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_672),
.B(n_66),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_731),
.B(n_18),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_745),
.A2(n_427),
.B1(n_413),
.B2(n_409),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_611),
.B(n_404),
.Y(n_906)
);

BUFx12f_ASAP7_75t_L g907 ( 
.A(n_604),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_729),
.A2(n_413),
.B(n_409),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_746),
.B(n_413),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_706),
.B(n_409),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_730),
.A2(n_409),
.B(n_427),
.Y(n_911)
);

BUFx12f_ASAP7_75t_L g912 ( 
.A(n_622),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_690),
.B(n_706),
.Y(n_913)
);

OAI21xp33_ASAP7_75t_L g914 ( 
.A1(n_655),
.A2(n_19),
.B(n_20),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_638),
.B(n_24),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_743),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_658),
.Y(n_917)
);

AO21x1_ASAP7_75t_L g918 ( 
.A1(n_635),
.A2(n_27),
.B(n_30),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_620),
.B(n_84),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_620),
.A2(n_427),
.B(n_85),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_733),
.A2(n_70),
.B1(n_151),
.B2(n_148),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_620),
.B(n_57),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_662),
.B(n_427),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_666),
.B(n_30),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_762),
.B(n_917),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_913),
.B(n_625),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_818),
.A2(n_670),
.B(n_740),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_750),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_900),
.A2(n_714),
.B(n_653),
.C(n_734),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_913),
.B(n_627),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_831),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_836),
.B(n_627),
.Y(n_932)
);

NOR2xp67_ASAP7_75t_SL g933 ( 
.A(n_763),
.B(n_691),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_900),
.A2(n_708),
.B(n_721),
.C(n_724),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_755),
.A2(n_895),
.B1(n_896),
.B2(n_804),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_813),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_761),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_754),
.B(n_638),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_873),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_769),
.B(n_638),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_836),
.B(n_627),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_824),
.A2(n_705),
.B(n_680),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_794),
.B(n_628),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_769),
.B(n_699),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_767),
.B(n_749),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_763),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_830),
.A2(n_749),
.B(n_718),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_883),
.A2(n_704),
.B(n_739),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_R g949 ( 
.A(n_890),
.B(n_699),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_813),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_907),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_767),
.B(n_35),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_R g953 ( 
.A(n_761),
.B(n_86),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_853),
.B(n_35),
.Y(n_954)
);

NOR2x1p5_ASAP7_75t_L g955 ( 
.A(n_912),
.B(n_613),
.Y(n_955)
);

INVx6_ASAP7_75t_L g956 ( 
.A(n_780),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_888),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_797),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_766),
.A2(n_130),
.B(n_125),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_846),
.B(n_37),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_903),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_SL g962 ( 
.A(n_914),
.B(n_120),
.Y(n_962)
);

NOR2x1_ASAP7_75t_L g963 ( 
.A(n_792),
.B(n_103),
.Y(n_963)
);

NOR3xp33_ASAP7_75t_SL g964 ( 
.A(n_915),
.B(n_38),
.C(n_41),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_879),
.B(n_101),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_846),
.B(n_38),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_894),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_753),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_857),
.B(n_43),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_792),
.B(n_94),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_888),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_770),
.A2(n_43),
.B(n_45),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_753),
.Y(n_973)
);

CKINVDCx11_ASAP7_75t_R g974 ( 
.A(n_764),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_802),
.B(n_854),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_804),
.A2(n_47),
.B1(n_55),
.B2(n_802),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_800),
.A2(n_750),
.B1(n_801),
.B2(n_872),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_753),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_753),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_832),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_773),
.A2(n_795),
.B(n_788),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_854),
.B(n_801),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_803),
.B(n_844),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_800),
.A2(n_751),
.B1(n_783),
.B2(n_790),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_807),
.A2(n_826),
.B(n_784),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_903),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_809),
.A2(n_811),
.B1(n_810),
.B2(n_869),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_897),
.A2(n_845),
.B(n_803),
.C(n_765),
.Y(n_988)
);

BUFx5_ASAP7_75t_L g989 ( 
.A(n_887),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_827),
.B(n_858),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_832),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_904),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_838),
.B(n_841),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_827),
.B(n_858),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_789),
.A2(n_851),
.B(n_760),
.C(n_924),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_851),
.B(n_760),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_758),
.B(n_759),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_869),
.A2(n_889),
.B1(n_876),
.B2(n_786),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_787),
.B(n_837),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_764),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_916),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_886),
.A2(n_881),
.B(n_885),
.C(n_918),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_757),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_796),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_817),
.B(n_888),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_805),
.A2(n_843),
.B1(n_891),
.B2(n_893),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_785),
.A2(n_909),
.B(n_768),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_782),
.A2(n_849),
.B(n_781),
.Y(n_1008)
);

NAND2xp33_ASAP7_75t_L g1009 ( 
.A(n_888),
.B(n_899),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_899),
.Y(n_1010)
);

INVx4_ASAP7_75t_L g1011 ( 
.A(n_899),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_839),
.A2(n_881),
.B1(n_764),
.B2(n_915),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_921),
.A2(n_848),
.B(n_922),
.C(n_919),
.Y(n_1013)
);

OA21x2_ASAP7_75t_L g1014 ( 
.A1(n_856),
.A2(n_816),
.B(n_752),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_899),
.B(n_832),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_805),
.A2(n_756),
.B1(n_819),
.B2(n_774),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_892),
.B(n_756),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_774),
.B(n_819),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_832),
.Y(n_1019)
);

INVxp67_ASAP7_75t_L g1020 ( 
.A(n_814),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_878),
.A2(n_882),
.B(n_866),
.C(n_910),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_820),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_861),
.B(n_822),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_840),
.B(n_902),
.Y(n_1024)
);

CKINVDCx11_ASAP7_75t_R g1025 ( 
.A(n_865),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_861),
.B(n_901),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_859),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_859),
.Y(n_1028)
);

XOR2x2_ASAP7_75t_SL g1029 ( 
.A(n_870),
.B(n_793),
.Y(n_1029)
);

AOI222xp33_ASAP7_75t_L g1030 ( 
.A1(n_847),
.A2(n_812),
.B1(n_771),
.B2(n_828),
.C1(n_829),
.C2(n_808),
.Y(n_1030)
);

AO21x1_ASAP7_75t_L g1031 ( 
.A1(n_808),
.A2(n_829),
.B(n_847),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_806),
.B(n_834),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_884),
.B(n_775),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_775),
.B(n_923),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_906),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_855),
.B(n_906),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_779),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_880),
.B(n_905),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_SL g1039 ( 
.A(n_821),
.B(n_920),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_863),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_799),
.A2(n_798),
.B(n_862),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_842),
.A2(n_772),
.B(n_877),
.C(n_864),
.Y(n_1042)
);

NOR3xp33_ASAP7_75t_SL g1043 ( 
.A(n_860),
.B(n_911),
.C(n_871),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_815),
.A2(n_867),
.B(n_833),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_777),
.A2(n_778),
.B(n_791),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_825),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_850),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_775),
.B(n_835),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_868),
.A2(n_875),
.B(n_898),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_852),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_908),
.Y(n_1051)
);

OR2x6_ASAP7_75t_L g1052 ( 
.A(n_874),
.B(n_685),
.Y(n_1052)
);

NAND2xp33_ASAP7_75t_SL g1053 ( 
.A(n_762),
.B(n_896),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_831),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_818),
.A2(n_556),
.B(n_823),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_762),
.A2(n_755),
.B1(n_900),
.B2(n_895),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_762),
.B(n_917),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_762),
.B(n_913),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_762),
.B(n_596),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_750),
.Y(n_1060)
);

AOI21x1_ASAP7_75t_L g1061 ( 
.A1(n_983),
.A2(n_1055),
.B(n_982),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_992),
.B(n_958),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_1054),
.Y(n_1063)
);

O2A1O1Ixp5_ASAP7_75t_L g1064 ( 
.A1(n_1059),
.A2(n_1056),
.B(n_1053),
.C(n_926),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_928),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_981),
.A2(n_1007),
.B(n_1021),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_961),
.B(n_986),
.Y(n_1067)
);

AO31x2_ASAP7_75t_L g1068 ( 
.A1(n_995),
.A2(n_1031),
.A3(n_1048),
.B(n_1056),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1060),
.Y(n_1069)
);

NAND2x1p5_ASAP7_75t_L g1070 ( 
.A(n_946),
.B(n_931),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_937),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_1057),
.B(n_925),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_1008),
.A2(n_994),
.B(n_990),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_975),
.A2(n_1058),
.B1(n_934),
.B2(n_1012),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_950),
.Y(n_1075)
);

AO31x2_ASAP7_75t_L g1076 ( 
.A1(n_1006),
.A2(n_935),
.A3(n_1042),
.B(n_1041),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_962),
.A2(n_954),
.B1(n_935),
.B2(n_943),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_985),
.A2(n_999),
.B(n_927),
.Y(n_1078)
);

OA21x2_ASAP7_75t_L g1079 ( 
.A1(n_947),
.A2(n_1032),
.B(n_999),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_997),
.A2(n_948),
.B(n_1013),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_992),
.B(n_958),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_993),
.B(n_945),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_988),
.A2(n_998),
.B(n_1006),
.Y(n_1083)
);

NOR2xp67_ASAP7_75t_SL g1084 ( 
.A(n_951),
.B(n_939),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_949),
.Y(n_1085)
);

AOI21x1_ASAP7_75t_L g1086 ( 
.A1(n_942),
.A2(n_996),
.B(n_966),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_998),
.A2(n_932),
.B(n_941),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1043),
.A2(n_1038),
.B(n_960),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_SL g1089 ( 
.A(n_962),
.B(n_929),
.Y(n_1089)
);

NAND3x1_ASAP7_75t_L g1090 ( 
.A(n_938),
.B(n_944),
.C(n_940),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_SL g1091 ( 
.A1(n_930),
.A2(n_976),
.B(n_987),
.C(n_1002),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_969),
.B(n_1020),
.Y(n_1092)
);

AOI21x1_ASAP7_75t_SL g1093 ( 
.A1(n_970),
.A2(n_965),
.B(n_1034),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1001),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_SL g1095 ( 
.A1(n_1052),
.A2(n_970),
.B(n_987),
.Y(n_1095)
);

OR2x6_ASAP7_75t_L g1096 ( 
.A(n_965),
.B(n_1027),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1024),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_976),
.A2(n_984),
.B1(n_977),
.B2(n_1040),
.Y(n_1098)
);

OA21x2_ASAP7_75t_L g1099 ( 
.A1(n_1050),
.A2(n_1049),
.B(n_1044),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_964),
.A2(n_972),
.B(n_984),
.C(n_952),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1016),
.A2(n_1046),
.B(n_1047),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1003),
.B(n_1022),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1016),
.A2(n_1014),
.B(n_1033),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1004),
.B(n_1037),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1009),
.A2(n_1039),
.B(n_1052),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1017),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_SL g1107 ( 
.A(n_1000),
.B(n_1019),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_989),
.B(n_1026),
.Y(n_1108)
);

BUFx2_ASAP7_75t_R g1109 ( 
.A(n_1005),
.Y(n_1109)
);

INVxp67_ASAP7_75t_L g1110 ( 
.A(n_1026),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_1036),
.A2(n_959),
.A3(n_1029),
.B(n_1018),
.Y(n_1111)
);

NAND3xp33_ASAP7_75t_L g1112 ( 
.A(n_1030),
.B(n_1025),
.C(n_933),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1051),
.A2(n_1015),
.B(n_1023),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1028),
.A2(n_963),
.B(n_1019),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1028),
.A2(n_971),
.B(n_957),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_957),
.A2(n_971),
.B(n_1011),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1035),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1010),
.A2(n_989),
.B(n_1035),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_SL g1119 ( 
.A1(n_989),
.A2(n_1035),
.B(n_991),
.C(n_980),
.Y(n_1119)
);

INVx3_ASAP7_75t_SL g1120 ( 
.A(n_956),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_968),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_968),
.A2(n_980),
.B(n_979),
.Y(n_1122)
);

AO31x2_ASAP7_75t_L g1123 ( 
.A1(n_989),
.A2(n_973),
.A3(n_980),
.B(n_979),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_989),
.B(n_973),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_953),
.A2(n_974),
.B1(n_955),
.B2(n_973),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_968),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_978),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_967),
.B(n_978),
.Y(n_1128)
);

INVx4_ASAP7_75t_L g1129 ( 
.A(n_978),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_979),
.B(n_991),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_956),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_981),
.A2(n_762),
.B(n_1055),
.Y(n_1132)
);

AOI221xp5_ASAP7_75t_L g1133 ( 
.A1(n_1056),
.A2(n_641),
.B1(n_419),
.B2(n_900),
.C(n_408),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_928),
.Y(n_1134)
);

NOR2x1_ASAP7_75t_SL g1135 ( 
.A(n_977),
.B(n_817),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1056),
.A2(n_762),
.B(n_995),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1059),
.B(n_1057),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_981),
.A2(n_762),
.B(n_1055),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_SL g1139 ( 
.A1(n_1056),
.A2(n_800),
.B(n_1013),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_967),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_992),
.B(n_602),
.Y(n_1141)
);

AO31x2_ASAP7_75t_L g1142 ( 
.A1(n_1021),
.A2(n_995),
.A3(n_1031),
.B(n_1048),
.Y(n_1142)
);

OR2x2_ASAP7_75t_L g1143 ( 
.A(n_1057),
.B(n_415),
.Y(n_1143)
);

AO21x1_ASAP7_75t_L g1144 ( 
.A1(n_1056),
.A2(n_762),
.B(n_1053),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1059),
.B(n_596),
.Y(n_1145)
);

INVx8_ASAP7_75t_L g1146 ( 
.A(n_968),
.Y(n_1146)
);

AO32x2_ASAP7_75t_L g1147 ( 
.A1(n_1056),
.A2(n_976),
.A3(n_935),
.B1(n_987),
.B2(n_998),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_981),
.A2(n_762),
.B(n_1055),
.Y(n_1148)
);

AOI21x1_ASAP7_75t_L g1149 ( 
.A1(n_983),
.A2(n_1055),
.B(n_982),
.Y(n_1149)
);

AO31x2_ASAP7_75t_L g1150 ( 
.A1(n_1021),
.A2(n_995),
.A3(n_1031),
.B(n_1048),
.Y(n_1150)
);

AOI31xp67_ASAP7_75t_L g1151 ( 
.A1(n_990),
.A2(n_895),
.A3(n_994),
.B(n_1058),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1056),
.A2(n_900),
.B1(n_762),
.B2(n_962),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_928),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1059),
.A2(n_762),
.B(n_913),
.C(n_900),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_936),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_992),
.B(n_602),
.Y(n_1156)
);

CKINVDCx16_ASAP7_75t_R g1157 ( 
.A(n_949),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_931),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1059),
.B(n_596),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_981),
.A2(n_762),
.B(n_1055),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1056),
.A2(n_762),
.B(n_1059),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1045),
.A2(n_856),
.B(n_816),
.Y(n_1162)
);

INVxp67_ASAP7_75t_L g1163 ( 
.A(n_931),
.Y(n_1163)
);

OA21x2_ASAP7_75t_L g1164 ( 
.A1(n_995),
.A2(n_981),
.B(n_1021),
.Y(n_1164)
);

AO32x2_ASAP7_75t_L g1165 ( 
.A1(n_1056),
.A2(n_976),
.A3(n_935),
.B1(n_987),
.B2(n_998),
.Y(n_1165)
);

AO31x2_ASAP7_75t_L g1166 ( 
.A1(n_1021),
.A2(n_995),
.A3(n_1031),
.B(n_1048),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_981),
.A2(n_762),
.B(n_1055),
.Y(n_1167)
);

NAND3x1_ASAP7_75t_L g1168 ( 
.A(n_938),
.B(n_641),
.C(n_596),
.Y(n_1168)
);

NAND3xp33_ASAP7_75t_L g1169 ( 
.A(n_1059),
.B(n_762),
.C(n_900),
.Y(n_1169)
);

NOR2xp67_ASAP7_75t_L g1170 ( 
.A(n_946),
.B(n_769),
.Y(n_1170)
);

BUFx4f_ASAP7_75t_L g1171 ( 
.A(n_956),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1059),
.A2(n_762),
.B(n_913),
.C(n_900),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_961),
.B(n_986),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_981),
.A2(n_762),
.B(n_1055),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_981),
.A2(n_762),
.B(n_1055),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1045),
.A2(n_856),
.B(n_816),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1021),
.A2(n_995),
.A3(n_1031),
.B(n_1048),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_928),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1059),
.A2(n_762),
.B1(n_900),
.B2(n_896),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_981),
.A2(n_762),
.B(n_1055),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_981),
.A2(n_762),
.B(n_1055),
.Y(n_1181)
);

AOI221xp5_ASAP7_75t_SL g1182 ( 
.A1(n_988),
.A2(n_900),
.B1(n_976),
.B2(n_1056),
.C(n_776),
.Y(n_1182)
);

AOI21x1_ASAP7_75t_L g1183 ( 
.A1(n_983),
.A2(n_1055),
.B(n_982),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1059),
.B(n_1057),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_1057),
.B(n_415),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1059),
.A2(n_762),
.B1(n_925),
.B2(n_1057),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_SL g1187 ( 
.A1(n_934),
.A2(n_762),
.B(n_1056),
.C(n_900),
.Y(n_1187)
);

INVxp67_ASAP7_75t_L g1188 ( 
.A(n_1063),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1069),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1133),
.A2(n_1159),
.B1(n_1145),
.B2(n_1089),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1101),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1134),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1089),
.A2(n_1169),
.B1(n_1161),
.B2(n_1179),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1072),
.B(n_1137),
.Y(n_1194)
);

BUFx12f_ASAP7_75t_L g1195 ( 
.A(n_1158),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1184),
.B(n_1186),
.Y(n_1196)
);

OAI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1152),
.A2(n_1169),
.B1(n_1098),
.B2(n_1077),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1146),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1146),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1121),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1152),
.A2(n_1172),
.B1(n_1154),
.B2(n_1098),
.Y(n_1201)
);

CKINVDCx11_ASAP7_75t_R g1202 ( 
.A(n_1140),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1136),
.A2(n_1074),
.B1(n_1083),
.B2(n_1077),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1129),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1153),
.Y(n_1205)
);

BUFx8_ASAP7_75t_L g1206 ( 
.A(n_1128),
.Y(n_1206)
);

INVx6_ASAP7_75t_L g1207 ( 
.A(n_1129),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1083),
.A2(n_1112),
.B1(n_1144),
.B2(n_1087),
.Y(n_1208)
);

BUFx8_ASAP7_75t_L g1209 ( 
.A(n_1085),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1168),
.A2(n_1141),
.B1(n_1156),
.B2(n_1090),
.Y(n_1210)
);

CKINVDCx11_ASAP7_75t_R g1211 ( 
.A(n_1120),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1123),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1143),
.B(n_1185),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1112),
.A2(n_1087),
.B1(n_1088),
.B2(n_1082),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1125),
.A2(n_1157),
.B1(n_1096),
.B2(n_1092),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1178),
.Y(n_1216)
);

BUFx10_ASAP7_75t_L g1217 ( 
.A(n_1067),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1062),
.B(n_1081),
.Y(n_1218)
);

BUFx12f_ASAP7_75t_L g1219 ( 
.A(n_1071),
.Y(n_1219)
);

INVx6_ASAP7_75t_L g1220 ( 
.A(n_1121),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1171),
.Y(n_1221)
);

INVx6_ASAP7_75t_L g1222 ( 
.A(n_1121),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_1131),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_SL g1224 ( 
.A1(n_1107),
.A2(n_1171),
.B1(n_1088),
.B2(n_1164),
.Y(n_1224)
);

BUFx8_ASAP7_75t_SL g1225 ( 
.A(n_1173),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1075),
.Y(n_1226)
);

NAND2x1p5_ASAP7_75t_L g1227 ( 
.A(n_1108),
.B(n_1115),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_SL g1228 ( 
.A1(n_1107),
.A2(n_1164),
.B1(n_1105),
.B2(n_1135),
.Y(n_1228)
);

INVx6_ASAP7_75t_L g1229 ( 
.A(n_1173),
.Y(n_1229)
);

INVx6_ASAP7_75t_L g1230 ( 
.A(n_1070),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1097),
.A2(n_1080),
.B1(n_1106),
.B2(n_1182),
.Y(n_1231)
);

BUFx12f_ASAP7_75t_L g1232 ( 
.A(n_1126),
.Y(n_1232)
);

OAI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1104),
.A2(n_1182),
.B1(n_1094),
.B2(n_1102),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1163),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1068),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1110),
.B(n_1187),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1109),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1155),
.Y(n_1238)
);

BUFx4f_ASAP7_75t_SL g1239 ( 
.A(n_1117),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1130),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1095),
.A2(n_1170),
.B1(n_1100),
.B2(n_1139),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1073),
.A2(n_1079),
.B1(n_1066),
.B2(n_1175),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1079),
.A2(n_1174),
.B1(n_1181),
.B2(n_1132),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1127),
.B(n_1064),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1123),
.Y(n_1245)
);

CKINVDCx16_ASAP7_75t_R g1246 ( 
.A(n_1118),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1138),
.A2(n_1180),
.B1(n_1160),
.B2(n_1148),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1167),
.A2(n_1165),
.B1(n_1147),
.B2(n_1084),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1123),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1124),
.Y(n_1250)
);

INVx6_ASAP7_75t_L g1251 ( 
.A(n_1170),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1091),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1114),
.A2(n_1086),
.B1(n_1113),
.B2(n_1183),
.Y(n_1253)
);

INVx6_ASAP7_75t_L g1254 ( 
.A(n_1093),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1061),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1147),
.A2(n_1165),
.B1(n_1099),
.B2(n_1078),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1122),
.Y(n_1257)
);

BUFx4_ASAP7_75t_SL g1258 ( 
.A(n_1119),
.Y(n_1258)
);

BUFx12f_ASAP7_75t_L g1259 ( 
.A(n_1151),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1116),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_1103),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1149),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1165),
.A2(n_1076),
.B1(n_1111),
.B2(n_1068),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1162),
.A2(n_1176),
.B1(n_1111),
.B2(n_1076),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1076),
.A2(n_1068),
.B1(n_1111),
.B2(n_1142),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1142),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1142),
.A2(n_1150),
.B1(n_1166),
.B2(n_1177),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1150),
.A2(n_1133),
.B1(n_1159),
.B2(n_1145),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_SL g1269 ( 
.A1(n_1166),
.A2(n_1089),
.B1(n_1159),
.B2(n_1145),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1166),
.A2(n_1133),
.B1(n_1159),
.B2(n_1145),
.Y(n_1270)
);

BUFx4f_ASAP7_75t_SL g1271 ( 
.A(n_1177),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1177),
.A2(n_1133),
.B1(n_1159),
.B2(n_1145),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1133),
.A2(n_1159),
.B1(n_1145),
.B2(n_900),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1133),
.A2(n_1159),
.B1(n_1145),
.B2(n_900),
.Y(n_1274)
);

AO22x1_ASAP7_75t_L g1275 ( 
.A1(n_1145),
.A2(n_596),
.B1(n_900),
.B2(n_1159),
.Y(n_1275)
);

INVx6_ASAP7_75t_L g1276 ( 
.A(n_1146),
.Y(n_1276)
);

BUFx2_ASAP7_75t_R g1277 ( 
.A(n_1120),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1140),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1141),
.B(n_1156),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1158),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1133),
.A2(n_1159),
.B1(n_1145),
.B2(n_900),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1065),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1089),
.A2(n_1159),
.B1(n_1145),
.B2(n_762),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_1140),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1158),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1089),
.A2(n_1159),
.B1(n_1145),
.B2(n_762),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1140),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1089),
.A2(n_1159),
.B1(n_1145),
.B2(n_762),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1133),
.A2(n_1159),
.B1(n_1145),
.B2(n_900),
.Y(n_1289)
);

INVx6_ASAP7_75t_L g1290 ( 
.A(n_1146),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1065),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1133),
.A2(n_1159),
.B1(n_1145),
.B2(n_900),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1133),
.A2(n_1159),
.B1(n_1145),
.B2(n_900),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1145),
.A2(n_1159),
.B1(n_1059),
.B2(n_762),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1140),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1133),
.A2(n_1159),
.B1(n_1145),
.B2(n_900),
.Y(n_1296)
);

BUFx12f_ASAP7_75t_L g1297 ( 
.A(n_1158),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1245),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1254),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1249),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1243),
.A2(n_1242),
.B(n_1247),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1243),
.A2(n_1253),
.B(n_1255),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1201),
.A2(n_1294),
.B1(n_1241),
.B2(n_1215),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1259),
.Y(n_1304)
);

AOI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1191),
.A2(n_1196),
.B(n_1262),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1244),
.B(n_1212),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1203),
.B(n_1248),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1273),
.A2(n_1281),
.B(n_1274),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1203),
.B(n_1248),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1208),
.B(n_1250),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1188),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1235),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1208),
.B(n_1266),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1283),
.B(n_1286),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1191),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1271),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1263),
.Y(n_1317)
);

OA21x2_ASAP7_75t_L g1318 ( 
.A1(n_1256),
.A2(n_1267),
.B(n_1265),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1265),
.B(n_1267),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1269),
.B(n_1268),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1273),
.A2(n_1274),
.B1(n_1281),
.B2(n_1293),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1212),
.Y(n_1322)
);

OAI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1210),
.A2(n_1194),
.B1(n_1197),
.B2(n_1237),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1268),
.B(n_1270),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1271),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1189),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1197),
.B(n_1214),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1227),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1192),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1230),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1254),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1264),
.A2(n_1256),
.B(n_1231),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1214),
.B(n_1218),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_1252),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1288),
.B(n_1190),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1190),
.A2(n_1292),
.B1(n_1289),
.B2(n_1293),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1205),
.Y(n_1337)
);

INVx8_ASAP7_75t_L g1338 ( 
.A(n_1232),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1261),
.B(n_1216),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1270),
.B(n_1272),
.Y(n_1340)
);

AOI21xp33_ASAP7_75t_L g1341 ( 
.A1(n_1289),
.A2(n_1296),
.B(n_1292),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1282),
.Y(n_1342)
);

INVxp33_ASAP7_75t_L g1343 ( 
.A(n_1279),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1272),
.B(n_1193),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1291),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1202),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1260),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1240),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_R g1349 ( 
.A(n_1284),
.B(n_1295),
.Y(n_1349)
);

INVx2_ASAP7_75t_SL g1350 ( 
.A(n_1230),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1226),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1240),
.B(n_1238),
.Y(n_1352)
);

INVxp33_ASAP7_75t_L g1353 ( 
.A(n_1213),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1233),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1240),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1233),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1224),
.A2(n_1257),
.B1(n_1234),
.B2(n_1236),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1280),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1230),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1251),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1228),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1258),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1251),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1275),
.A2(n_1204),
.B(n_1285),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_SL g1365 ( 
.A(n_1277),
.B(n_1221),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1251),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1229),
.A2(n_1297),
.B1(n_1195),
.B2(n_1285),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1246),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1258),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1239),
.A2(n_1200),
.B(n_1220),
.Y(n_1370)
);

AND2x2_ASAP7_75t_SL g1371 ( 
.A(n_1225),
.B(n_1206),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1229),
.B(n_1287),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1303),
.B(n_1323),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1368),
.B(n_1278),
.Y(n_1374)
);

BUFx5_ASAP7_75t_L g1375 ( 
.A(n_1322),
.Y(n_1375)
);

O2A1O1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1321),
.A2(n_1198),
.B(n_1199),
.C(n_1223),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1326),
.Y(n_1377)
);

AO22x2_ASAP7_75t_L g1378 ( 
.A1(n_1327),
.A2(n_1198),
.B1(n_1199),
.B2(n_1239),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1308),
.A2(n_1217),
.B(n_1229),
.Y(n_1379)
);

INVx5_ASAP7_75t_SL g1380 ( 
.A(n_1371),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1348),
.B(n_1206),
.Y(n_1381)
);

O2A1O1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1341),
.A2(n_1217),
.B(n_1209),
.C(n_1219),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1336),
.A2(n_1209),
.B(n_1207),
.C(n_1290),
.Y(n_1383)
);

NAND4xp25_ASAP7_75t_L g1384 ( 
.A(n_1335),
.B(n_1211),
.C(n_1222),
.D(n_1207),
.Y(n_1384)
);

NOR2x1p5_ASAP7_75t_L g1385 ( 
.A(n_1333),
.B(n_1276),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1314),
.B(n_1276),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1301),
.A2(n_1290),
.B(n_1347),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1355),
.B(n_1343),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1329),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1313),
.B(n_1352),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1313),
.B(n_1352),
.Y(n_1391)
);

CKINVDCx11_ASAP7_75t_R g1392 ( 
.A(n_1338),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1352),
.B(n_1310),
.Y(n_1393)
);

AOI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1327),
.A2(n_1344),
.B1(n_1320),
.B2(n_1357),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1344),
.A2(n_1356),
.B(n_1354),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1310),
.B(n_1361),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1349),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1305),
.A2(n_1302),
.B(n_1356),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1352),
.B(n_1358),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1360),
.B(n_1363),
.Y(n_1400)
);

AO32x1_ASAP7_75t_L g1401 ( 
.A1(n_1320),
.A2(n_1361),
.A3(n_1354),
.B1(n_1300),
.B2(n_1298),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1353),
.B(n_1364),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1307),
.B(n_1309),
.Y(n_1403)
);

NOR2x1_ASAP7_75t_SL g1404 ( 
.A(n_1305),
.B(n_1299),
.Y(n_1404)
);

INVxp67_ASAP7_75t_L g1405 ( 
.A(n_1315),
.Y(n_1405)
);

AND2x2_ASAP7_75t_SL g1406 ( 
.A(n_1316),
.B(n_1324),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1324),
.A2(n_1340),
.B(n_1347),
.Y(n_1407)
);

O2A1O1Ixp33_ASAP7_75t_SL g1408 ( 
.A1(n_1362),
.A2(n_1369),
.B(n_1334),
.C(n_1330),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1366),
.B(n_1345),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1340),
.A2(n_1309),
.B(n_1307),
.C(n_1332),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1317),
.B(n_1347),
.Y(n_1411)
);

NAND3xp33_ASAP7_75t_L g1412 ( 
.A(n_1347),
.B(n_1311),
.C(n_1366),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1312),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1337),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1393),
.B(n_1332),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1413),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1373),
.A2(n_1304),
.B1(n_1325),
.B2(n_1331),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1377),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1411),
.B(n_1306),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1398),
.B(n_1306),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1411),
.B(n_1312),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1389),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1398),
.B(n_1306),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1403),
.B(n_1342),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1390),
.B(n_1318),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1405),
.Y(n_1426)
);

NOR2x1_ASAP7_75t_L g1427 ( 
.A(n_1412),
.B(n_1328),
.Y(n_1427)
);

INVxp67_ASAP7_75t_L g1428 ( 
.A(n_1402),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1391),
.B(n_1318),
.Y(n_1429)
);

NAND2x1_ASAP7_75t_L g1430 ( 
.A(n_1378),
.B(n_1370),
.Y(n_1430)
);

AO21x2_ASAP7_75t_L g1431 ( 
.A1(n_1387),
.A2(n_1302),
.B(n_1322),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1402),
.A2(n_1304),
.B1(n_1331),
.B2(n_1299),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1384),
.B(n_1372),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1414),
.B(n_1318),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1407),
.B(n_1318),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1407),
.B(n_1319),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1409),
.B(n_1319),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1410),
.B(n_1298),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_L g1439 ( 
.A(n_1394),
.B(n_1299),
.C(n_1351),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1375),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1418),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1425),
.B(n_1406),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1438),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1425),
.B(n_1406),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1419),
.B(n_1387),
.Y(n_1445)
);

AOI221xp5_ASAP7_75t_L g1446 ( 
.A1(n_1428),
.A2(n_1396),
.B1(n_1395),
.B2(n_1376),
.C(n_1379),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1427),
.A2(n_1404),
.B(n_1408),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1439),
.A2(n_1380),
.B1(n_1379),
.B2(n_1396),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1428),
.B(n_1395),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1419),
.B(n_1399),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1418),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1425),
.B(n_1388),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1420),
.B(n_1400),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1416),
.Y(n_1454)
);

INVxp67_ASAP7_75t_L g1455 ( 
.A(n_1438),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1418),
.Y(n_1456)
);

INVxp67_ASAP7_75t_L g1457 ( 
.A(n_1438),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1422),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1426),
.B(n_1421),
.Y(n_1459)
);

OR2x6_ASAP7_75t_L g1460 ( 
.A(n_1430),
.B(n_1378),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1426),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1430),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1421),
.B(n_1339),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1427),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1429),
.B(n_1375),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1429),
.B(n_1415),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1439),
.A2(n_1401),
.B(n_1376),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1460),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1455),
.B(n_1437),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1466),
.B(n_1423),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1443),
.B(n_1421),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1441),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1449),
.B(n_1433),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1441),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1441),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1455),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1451),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1451),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1462),
.B(n_1440),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1465),
.B(n_1435),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1443),
.B(n_1435),
.Y(n_1481)
);

INVxp67_ASAP7_75t_L g1482 ( 
.A(n_1449),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1465),
.B(n_1435),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1457),
.B(n_1429),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1456),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1457),
.B(n_1445),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1447),
.B(n_1436),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1460),
.B(n_1415),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1460),
.B(n_1415),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1456),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1460),
.B(n_1434),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1459),
.B(n_1437),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1447),
.B(n_1436),
.Y(n_1493)
);

INVxp67_ASAP7_75t_SL g1494 ( 
.A(n_1454),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1460),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1448),
.B(n_1436),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1456),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1442),
.B(n_1434),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1442),
.B(n_1434),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1444),
.B(n_1431),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1471),
.B(n_1445),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1495),
.B(n_1468),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1476),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1475),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1471),
.B(n_1463),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1469),
.B(n_1450),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1476),
.Y(n_1507)
);

OAI21xp33_ASAP7_75t_SL g1508 ( 
.A1(n_1487),
.A2(n_1464),
.B(n_1444),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1471),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1487),
.Y(n_1510)
);

AND2x2_ASAP7_75t_SL g1511 ( 
.A(n_1473),
.B(n_1371),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1471),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1469),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1473),
.B(n_1452),
.Y(n_1514)
);

NOR2x1p5_ASAP7_75t_SL g1515 ( 
.A(n_1475),
.B(n_1458),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1494),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1496),
.A2(n_1448),
.B1(n_1446),
.B2(n_1467),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1482),
.B(n_1452),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1494),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1472),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1492),
.B(n_1450),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1482),
.B(n_1453),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1472),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1472),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1496),
.A2(n_1493),
.B1(n_1446),
.B2(n_1467),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1474),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1474),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1486),
.B(n_1453),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1486),
.B(n_1453),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1475),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1474),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1475),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1481),
.B(n_1463),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1485),
.Y(n_1534)
);

NOR2x1p5_ASAP7_75t_L g1535 ( 
.A(n_1468),
.B(n_1397),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1493),
.B(n_1453),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1485),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1468),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1485),
.Y(n_1539)
);

AND2x4_ASAP7_75t_SL g1540 ( 
.A(n_1495),
.B(n_1381),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1481),
.B(n_1461),
.Y(n_1541)
);

OAI21xp33_ASAP7_75t_L g1542 ( 
.A1(n_1500),
.A2(n_1417),
.B(n_1424),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1507),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1507),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1503),
.B(n_1484),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1520),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1525),
.B(n_1484),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1502),
.B(n_1495),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1504),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1516),
.B(n_1481),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1502),
.B(n_1495),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1519),
.B(n_1481),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1540),
.B(n_1495),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1510),
.B(n_1484),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1523),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1540),
.B(n_1495),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1517),
.A2(n_1468),
.B1(n_1488),
.B2(n_1489),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1511),
.B(n_1538),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1511),
.B(n_1488),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1538),
.B(n_1488),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1542),
.B(n_1484),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1515),
.B(n_1488),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1524),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1513),
.B(n_1489),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1514),
.B(n_1498),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1526),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1527),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1541),
.Y(n_1568)
);

NAND2x1_ASAP7_75t_L g1569 ( 
.A(n_1536),
.B(n_1489),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1509),
.B(n_1489),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1504),
.Y(n_1571)
);

AOI221xp5_ASAP7_75t_L g1572 ( 
.A1(n_1508),
.A2(n_1464),
.B1(n_1500),
.B2(n_1491),
.C(n_1382),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1528),
.B(n_1380),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1512),
.B(n_1491),
.Y(n_1574)
);

XNOR2x1_ASAP7_75t_L g1575 ( 
.A(n_1535),
.B(n_1346),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1529),
.B(n_1371),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1518),
.B(n_1492),
.Y(n_1577)
);

NOR3xp33_ASAP7_75t_L g1578 ( 
.A(n_1544),
.B(n_1382),
.C(n_1501),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_1558),
.Y(n_1579)
);

OAI21xp33_ASAP7_75t_L g1580 ( 
.A1(n_1557),
.A2(n_1501),
.B(n_1522),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1547),
.A2(n_1380),
.B1(n_1541),
.B2(n_1500),
.Y(n_1581)
);

A2O1A1Ixp33_ASAP7_75t_L g1582 ( 
.A1(n_1547),
.A2(n_1500),
.B(n_1491),
.C(n_1462),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1559),
.A2(n_1491),
.B1(n_1505),
.B2(n_1506),
.Y(n_1583)
);

AOI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1572),
.A2(n_1539),
.B1(n_1537),
.B2(n_1534),
.C(n_1531),
.Y(n_1584)
);

NOR2x1_ASAP7_75t_L g1585 ( 
.A(n_1544),
.B(n_1462),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1568),
.B(n_1498),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1568),
.B(n_1558),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1559),
.A2(n_1378),
.B1(n_1386),
.B2(n_1480),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1543),
.B(n_1470),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1553),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1543),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1576),
.B(n_1498),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1575),
.B(n_1521),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1553),
.B(n_1498),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1565),
.B(n_1505),
.Y(n_1595)
);

INVxp67_ASAP7_75t_L g1596 ( 
.A(n_1543),
.Y(n_1596)
);

OAI321xp33_ASAP7_75t_L g1597 ( 
.A1(n_1561),
.A2(n_1533),
.A3(n_1386),
.B1(n_1530),
.B2(n_1532),
.C(n_1432),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1560),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1546),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1575),
.A2(n_1338),
.B(n_1533),
.Y(n_1600)
);

OR2x6_ASAP7_75t_L g1601 ( 
.A(n_1556),
.B(n_1338),
.Y(n_1601)
);

AOI321xp33_ASAP7_75t_L g1602 ( 
.A1(n_1561),
.A2(n_1480),
.A3(n_1483),
.B1(n_1383),
.B2(n_1499),
.C(n_1367),
.Y(n_1602)
);

XNOR2xp5_ASAP7_75t_L g1603 ( 
.A(n_1575),
.B(n_1385),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1579),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1579),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1588),
.A2(n_1572),
.B1(n_1569),
.B2(n_1573),
.Y(n_1606)
);

NAND3xp33_ASAP7_75t_L g1607 ( 
.A(n_1584),
.B(n_1551),
.C(n_1548),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1593),
.A2(n_1569),
.B1(n_1562),
.B2(n_1565),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1591),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1589),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1590),
.A2(n_1548),
.B1(n_1551),
.B2(n_1556),
.Y(n_1611)
);

AOI322xp5_ASAP7_75t_L g1612 ( 
.A1(n_1580),
.A2(n_1554),
.A3(n_1562),
.B1(n_1564),
.B2(n_1545),
.C1(n_1570),
.C2(n_1574),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1587),
.B(n_1560),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1589),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1596),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_SL g1616 ( 
.A1(n_1603),
.A2(n_1562),
.B(n_1554),
.Y(n_1616)
);

OAI221xp5_ASAP7_75t_L g1617 ( 
.A1(n_1602),
.A2(n_1545),
.B1(n_1550),
.B2(n_1552),
.C(n_1577),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1598),
.B(n_1564),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1599),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1586),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1594),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1595),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1604),
.Y(n_1623)
);

NOR3xp33_ASAP7_75t_L g1624 ( 
.A(n_1615),
.B(n_1597),
.C(n_1600),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1605),
.B(n_1578),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1610),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1610),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1614),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1614),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1609),
.Y(n_1630)
);

AO22x2_ASAP7_75t_L g1631 ( 
.A1(n_1619),
.A2(n_1608),
.B1(n_1606),
.B2(n_1622),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1618),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1613),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1624),
.A2(n_1616),
.B(n_1597),
.Y(n_1634)
);

OAI211xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1625),
.A2(n_1616),
.B(n_1623),
.C(n_1633),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1631),
.A2(n_1617),
.B1(n_1607),
.B2(n_1581),
.C(n_1620),
.Y(n_1636)
);

NOR3xp33_ASAP7_75t_L g1637 ( 
.A(n_1632),
.B(n_1581),
.C(n_1621),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1626),
.Y(n_1638)
);

CKINVDCx20_ASAP7_75t_R g1639 ( 
.A(n_1633),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1627),
.B(n_1611),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1628),
.B(n_1601),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1629),
.B(n_1631),
.Y(n_1642)
);

AOI211xp5_ASAP7_75t_L g1643 ( 
.A1(n_1635),
.A2(n_1630),
.B(n_1582),
.C(n_1562),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1639),
.A2(n_1601),
.B1(n_1585),
.B2(n_1583),
.Y(n_1644)
);

AOI211xp5_ASAP7_75t_L g1645 ( 
.A1(n_1634),
.A2(n_1592),
.B(n_1552),
.C(n_1550),
.Y(n_1645)
);

OAI211xp5_ASAP7_75t_L g1646 ( 
.A1(n_1636),
.A2(n_1612),
.B(n_1563),
.C(n_1555),
.Y(n_1646)
);

NAND3xp33_ASAP7_75t_L g1647 ( 
.A(n_1642),
.B(n_1601),
.C(n_1555),
.Y(n_1647)
);

NOR4xp25_ASAP7_75t_L g1648 ( 
.A(n_1646),
.B(n_1638),
.C(n_1640),
.D(n_1641),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1643),
.B(n_1644),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1645),
.A2(n_1637),
.B1(n_1577),
.B2(n_1567),
.Y(n_1650)
);

AOI221xp5_ASAP7_75t_L g1651 ( 
.A1(n_1647),
.A2(n_1546),
.B1(n_1563),
.B2(n_1567),
.C(n_1566),
.Y(n_1651)
);

NOR2xp67_ASAP7_75t_L g1652 ( 
.A(n_1647),
.B(n_1566),
.Y(n_1652)
);

XNOR2xp5_ASAP7_75t_L g1653 ( 
.A(n_1644),
.B(n_1381),
.Y(n_1653)
);

XNOR2xp5_ASAP7_75t_L g1654 ( 
.A(n_1648),
.B(n_1574),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1652),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1649),
.B(n_1570),
.Y(n_1656)
);

NAND4xp75_ASAP7_75t_L g1657 ( 
.A(n_1651),
.B(n_1549),
.C(n_1362),
.D(n_1532),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1653),
.B(n_1549),
.Y(n_1658)
);

NAND3xp33_ASAP7_75t_L g1659 ( 
.A(n_1654),
.B(n_1650),
.C(n_1549),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1656),
.Y(n_1660)
);

O2A1O1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1655),
.A2(n_1571),
.B(n_1365),
.C(n_1530),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1660),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1662),
.A2(n_1654),
.B1(n_1658),
.B2(n_1659),
.Y(n_1663)
);

OAI22x1_ASAP7_75t_L g1664 ( 
.A1(n_1663),
.A2(n_1661),
.B1(n_1657),
.B2(n_1571),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1663),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1664),
.Y(n_1666)
);

INVxp33_ASAP7_75t_SL g1667 ( 
.A(n_1665),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1667),
.A2(n_1338),
.B(n_1571),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1666),
.A2(n_1338),
.B(n_1571),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1669),
.A2(n_1392),
.B1(n_1479),
.B2(n_1478),
.Y(n_1670)
);

OAI21xp33_ASAP7_75t_L g1671 ( 
.A1(n_1670),
.A2(n_1668),
.B(n_1374),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1671),
.Y(n_1672)
);

AOI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1672),
.A2(n_1479),
.B1(n_1497),
.B2(n_1490),
.C(n_1477),
.Y(n_1673)
);

AOI211xp5_ASAP7_75t_L g1674 ( 
.A1(n_1673),
.A2(n_1369),
.B(n_1359),
.C(n_1350),
.Y(n_1674)
);


endmodule