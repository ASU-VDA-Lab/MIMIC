module fake_jpeg_9851_n_116 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_116);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_29),
.Y(n_41)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_1),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_1),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_10),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_29),
.B(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_18),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_15),
.C(n_16),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_17),
.B1(n_13),
.B2(n_23),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_36),
.B1(n_31),
.B2(n_32),
.Y(n_67)
);

OR2x4_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_2),
.Y(n_64)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_38),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_47),
.A2(n_28),
.B1(n_26),
.B2(n_21),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_57),
.B1(n_51),
.B2(n_39),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_56),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_15),
.B(n_16),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_50),
.B(n_4),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_47),
.A2(n_24),
.B1(n_20),
.B2(n_22),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_65),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_22),
.B1(n_18),
.B2(n_13),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_67),
.B1(n_48),
.B2(n_39),
.Y(n_79)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_73),
.B1(n_52),
.B2(n_67),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_48),
.A3(n_50),
.B1(n_32),
.B2(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_75),
.B(n_79),
.Y(n_84)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_55),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_6),
.C(n_8),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_81),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_56),
.B(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_88),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_38),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_58),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_78),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_84),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_94),
.A2(n_74),
.B(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_101),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_81),
.C(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_98),
.B(n_96),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_84),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_100),
.C(n_93),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_83),
.C(n_82),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_90),
.B(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_105),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_90),
.B1(n_78),
.B2(n_37),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_105),
.A2(n_37),
.B1(n_49),
.B2(n_45),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_108),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_113),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_106),
.A3(n_107),
.B1(n_109),
.B2(n_11),
.C1(n_45),
.C2(n_3),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_45),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_3),
.Y(n_116)
);


endmodule