module fake_jpeg_31975_n_108 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_2),
.C(n_3),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_15),
.C(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_14),
.B(n_5),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_13),
.B(n_5),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_23),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_19),
.Y(n_34)
);

NAND2x1_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_37),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_22),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_34),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_24),
.B1(n_16),
.B2(n_11),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_11),
.B1(n_16),
.B2(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_52),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_15),
.B(n_13),
.Y(n_51)
);

AO21x1_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_56),
.B(n_22),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_25),
.B(n_21),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_47),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_60),
.A2(n_66),
.B1(n_40),
.B2(n_53),
.Y(n_78)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_70),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_36),
.B1(n_35),
.B2(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_36),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_69),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_46),
.B1(n_43),
.B2(n_47),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_6),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_76),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_22),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_7),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_7),
.C(n_8),
.Y(n_83)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx4f_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_85),
.B(n_88),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_64),
.C(n_67),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_92),
.C(n_83),
.Y(n_99)
);

A2O1A1O1Ixp25_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_73),
.B(n_74),
.C(n_77),
.D(n_75),
.Y(n_92)
);

AOI221xp5_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_73),
.B1(n_77),
.B2(n_68),
.C(n_78),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_79),
.B(n_61),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_77),
.B1(n_59),
.B2(n_61),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_79),
.B1(n_72),
.B2(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_97),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_95),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_98),
.B(n_90),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_102),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_92),
.C(n_63),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_100),
.B(n_82),
.Y(n_105)
);

OAI21x1_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_103),
.B(n_54),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_44),
.B(n_49),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_22),
.Y(n_108)
);


endmodule