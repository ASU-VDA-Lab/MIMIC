module fake_jpeg_29446_n_247 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_4),
.B(n_8),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_43),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_23),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_23),
.B(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_23),
.B(n_25),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_29),
.Y(n_58)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_32),
.Y(n_66)
);

BUFx12f_ASAP7_75t_SL g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_56),
.B(n_27),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_66),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_19),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_65),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_53),
.B1(n_44),
.B2(n_50),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_60),
.A2(n_62),
.B1(n_79),
.B2(n_5),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_21),
.B1(n_25),
.B2(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_70),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_21),
.B1(n_34),
.B2(n_35),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_31),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_31),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_33),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_36),
.B1(n_35),
.B2(n_28),
.Y(n_79)
);

OA22x2_ASAP7_75t_SL g80 ( 
.A1(n_40),
.A2(n_36),
.B1(n_28),
.B2(n_27),
.Y(n_80)
);

AO22x1_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_33),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_38),
.B(n_37),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_6),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_37),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_13),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_54),
.B1(n_30),
.B2(n_5),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_89),
.A2(n_107),
.B1(n_99),
.B2(n_91),
.Y(n_134)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_92),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_94),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_2),
.C(n_3),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_100),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_57),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_96),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_2),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_69),
.C(n_104),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_99),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_5),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_82),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_101),
.Y(n_141)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_104),
.Y(n_125)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_110),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_74),
.B(n_13),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_66),
.A2(n_10),
.B(n_11),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_111),
.A2(n_95),
.B(n_109),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_63),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_115),
.B1(n_119),
.B2(n_107),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_63),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_64),
.B1(n_76),
.B2(n_60),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_116),
.A2(n_61),
.B1(n_72),
.B2(n_78),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_81),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_14),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_110),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_76),
.B1(n_81),
.B2(n_86),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_57),
.B(n_78),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_137),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_96),
.B1(n_113),
.B2(n_94),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_124),
.A2(n_134),
.B1(n_142),
.B2(n_120),
.Y(n_156)
);

AOI32xp33_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_61),
.A3(n_72),
.B1(n_69),
.B2(n_81),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_118),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_133),
.A2(n_143),
.B(n_144),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_105),
.B(n_109),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_140),
.B(n_93),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_105),
.A2(n_101),
.B1(n_90),
.B2(n_114),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_97),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_102),
.B(n_88),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_141),
.A2(n_96),
.B1(n_103),
.B2(n_108),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_147),
.A2(n_159),
.B(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_149),
.A2(n_155),
.B1(n_164),
.B2(n_166),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_125),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_115),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_113),
.B1(n_121),
.B2(n_137),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_145),
.B1(n_146),
.B2(n_151),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_157),
.B(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_122),
.B(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_167),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_123),
.B1(n_124),
.B2(n_133),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_144),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_146),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_125),
.A2(n_143),
.B1(n_128),
.B2(n_129),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_125),
.B(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

NAND2xp33_ASAP7_75t_SL g172 ( 
.A(n_168),
.B(n_131),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_173),
.Y(n_196)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_130),
.C(n_131),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_171),
.B(n_177),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_161),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_130),
.C(n_150),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_175),
.C(n_179),
.Y(n_195)
);

NAND2xp67_ASAP7_75t_SL g174 ( 
.A(n_163),
.B(n_158),
.Y(n_174)
);

OAI322xp33_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_161),
.A3(n_185),
.B1(n_176),
.B2(n_187),
.C1(n_179),
.C2(n_169),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_155),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_188),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_146),
.C(n_156),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_164),
.B1(n_149),
.B2(n_152),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_189),
.A2(n_198),
.B1(n_200),
.B2(n_204),
.Y(n_216)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_181),
.A2(n_148),
.B1(n_160),
.B2(n_168),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_203),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_192),
.A2(n_178),
.B(n_204),
.Y(n_209)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_184),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_183),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_202),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_181),
.C(n_185),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_195),
.C(n_196),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_174),
.B1(n_182),
.B2(n_183),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_186),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_203),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_208),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_195),
.C(n_199),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_201),
.B(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_190),
.B(n_194),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_210),
.B(n_193),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

INVx11_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_221),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_225),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_191),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_214),
.C(n_205),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_192),
.C(n_207),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_215),
.C(n_211),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_215),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_209),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_229),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_210),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_232),
.C(n_205),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_230),
.A2(n_222),
.B(n_224),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_218),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_223),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_231),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_225),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_236),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_232),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_239),
.B(n_237),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_241),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_211),
.C(n_214),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_243),
.A2(n_240),
.B(n_238),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_245),
.A2(n_246),
.B(n_244),
.Y(n_247)
);


endmodule