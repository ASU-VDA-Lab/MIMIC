module fake_jpeg_12918_n_295 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx10_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_43),
.Y(n_102)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_29),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_51),
.Y(n_83)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_31),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_54),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_18),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_60),
.Y(n_61)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

HAxp5_ASAP7_75t_SL g59 ( 
.A(n_18),
.B(n_2),
.CON(n_59),
.SN(n_59)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_2),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_2),
.Y(n_60)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_40),
.B1(n_28),
.B2(n_41),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_67),
.A2(n_82),
.B1(n_89),
.B2(n_99),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_21),
.C(n_18),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_68),
.B(n_72),
.C(n_100),
.Y(n_131)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_90),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_21),
.C(n_18),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_23),
.B1(n_19),
.B2(n_35),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_74),
.A2(n_76),
.B1(n_81),
.B2(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_23),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_29),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_23),
.B1(n_19),
.B2(n_35),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_77),
.Y(n_114)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_41),
.B1(n_40),
.B2(n_19),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_80),
.A2(n_91),
.B1(n_98),
.B2(n_27),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_24),
.B1(n_38),
.B2(n_35),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_41),
.B1(n_40),
.B2(n_21),
.Y(n_82)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_84),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_42),
.A2(n_24),
.B1(n_38),
.B2(n_22),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_42),
.A2(n_24),
.B1(n_38),
.B2(n_21),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_88),
.A2(n_95),
.B1(n_25),
.B2(n_8),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_40),
.B1(n_41),
.B2(n_39),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_21),
.B1(n_39),
.B2(n_33),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_37),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_104),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_52),
.A2(n_21),
.B1(n_37),
.B2(n_36),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_43),
.A2(n_31),
.B1(n_34),
.B2(n_33),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_43),
.A2(n_36),
.B1(n_34),
.B2(n_32),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_60),
.B(n_26),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_32),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

CKINVDCx11_ASAP7_75t_R g154 ( 
.A(n_106),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_108),
.B(n_109),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_61),
.A2(n_75),
.B(n_100),
.C(n_83),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_102),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_3),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_3),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_27),
.B(n_26),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_118),
.A2(n_136),
.B(n_10),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_27),
.B1(n_25),
.B2(n_8),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_119),
.A2(n_135),
.B1(n_122),
.B2(n_116),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_101),
.B1(n_64),
.B2(n_69),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_4),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_128),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_68),
.B(n_4),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_5),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_5),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_63),
.B(n_5),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_65),
.Y(n_159)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_72),
.A2(n_25),
.B(n_8),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_63),
.A2(n_25),
.B(n_10),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_80),
.C(n_65),
.Y(n_150)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_85),
.B1(n_66),
.B2(n_70),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_141),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_144),
.A2(n_145),
.B1(n_155),
.B2(n_166),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_64),
.B1(n_79),
.B2(n_103),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_150),
.A2(n_136),
.B(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_73),
.B1(n_78),
.B2(n_96),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_109),
.A2(n_85),
.B(n_77),
.C(n_62),
.Y(n_156)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_143),
.B(n_144),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_158),
.C(n_161),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_159),
.B(n_168),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_164),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_131),
.A2(n_96),
.B1(n_78),
.B2(n_73),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_163),
.A2(n_111),
.B1(n_124),
.B2(n_134),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g165 ( 
.A(n_126),
.Y(n_165)
);

BUFx24_ASAP7_75t_SL g176 ( 
.A(n_165),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_93),
.B1(n_12),
.B2(n_13),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_110),
.B(n_11),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_128),
.A2(n_93),
.B1(n_12),
.B2(n_14),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_169),
.A2(n_170),
.B1(n_134),
.B2(n_106),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_113),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_170)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_171),
.A2(n_198),
.B(n_199),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_132),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_175),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_174),
.A2(n_198),
.B(n_194),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_108),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_126),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_178),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_162),
.B(n_110),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_112),
.B(n_138),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_192),
.B(n_164),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_123),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_169),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_196),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_123),
.C(n_121),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_151),
.A2(n_114),
.B(n_127),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_142),
.B(n_107),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_195),
.B(n_197),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_153),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_107),
.C(n_117),
.Y(n_197)
);

OR2x6_ASAP7_75t_SL g198 ( 
.A(n_156),
.B(n_115),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_142),
.B(n_115),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_151),
.B1(n_145),
.B2(n_140),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_202),
.A2(n_205),
.B1(n_214),
.B2(n_197),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_204),
.A2(n_206),
.B(n_211),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_140),
.B1(n_158),
.B2(n_147),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_207),
.B(n_183),
.Y(n_223)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_148),
.B(n_161),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_186),
.A2(n_115),
.B1(n_139),
.B2(n_146),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_212),
.A2(n_213),
.B1(n_179),
.B2(n_192),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_171),
.A2(n_170),
.B1(n_152),
.B2(n_146),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_179),
.A2(n_185),
.B1(n_195),
.B2(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_217),
.Y(n_225)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_167),
.Y(n_238)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_226),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_216),
.B(n_178),
.Y(n_224)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

XOR2x2_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_188),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_187),
.C(n_181),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_237),
.C(n_204),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_175),
.Y(n_229)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_203),
.B(n_172),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_230),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_171),
.B1(n_174),
.B2(n_198),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_231),
.A2(n_234),
.B1(n_211),
.B2(n_226),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_154),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_232),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_234),
.A2(n_210),
.B1(n_200),
.B2(n_205),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_206),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_196),
.C(n_193),
.Y(n_237)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_238),
.Y(n_248)
);

OAI22x1_ASAP7_75t_L g257 ( 
.A1(n_241),
.A2(n_231),
.B1(n_202),
.B2(n_233),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_242),
.A2(n_233),
.B(n_246),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_225),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_243),
.B(n_230),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_246),
.C(n_241),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g261 ( 
.A1(n_245),
.A2(n_236),
.B(n_237),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_200),
.C(n_212),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_218),
.Y(n_252)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_220),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_253),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_257),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_224),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_255),
.B(n_260),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_259),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_262),
.C(n_264),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_239),
.B1(n_222),
.B2(n_227),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_176),
.Y(n_260)
);

XOR2x2_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_242),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_228),
.C(n_223),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_239),
.Y(n_264)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_254),
.B(n_251),
.CI(n_245),
.CON(n_266),
.SN(n_266)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_272),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_274),
.Y(n_275)
);

OAI211xp5_ASAP7_75t_L g272 ( 
.A1(n_263),
.A2(n_248),
.B(n_240),
.C(n_252),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_248),
.C(n_253),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_209),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_222),
.B(n_215),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_277),
.Y(n_282)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_274),
.Y(n_277)
);

AND2x6_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_257),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_279),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_265),
.C(n_261),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_273),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_266),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_271),
.C(n_270),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_285),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_276),
.A2(n_269),
.B1(n_266),
.B2(n_235),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_275),
.C(n_278),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_288),
.B(n_289),
.C(n_285),
.Y(n_290)
);

OAI321xp33_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_291),
.A3(n_189),
.B1(n_191),
.B2(n_173),
.C(n_16),
.Y(n_292)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_287),
.A2(n_282),
.A3(n_268),
.B1(n_235),
.B2(n_221),
.C1(n_191),
.C2(n_167),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_173),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_11),
.B(n_15),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_15),
.Y(n_295)
);


endmodule