module fake_netlist_6_608_n_31 (n_7, n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_9, n_8, n_31);

input n_7;
input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;
input n_9;
input n_8;

output n_31;

wire n_16;
wire n_18;
wire n_21;
wire n_10;
wire n_24;
wire n_15;
wire n_27;
wire n_14;
wire n_22;
wire n_26;
wire n_13;
wire n_11;
wire n_28;
wire n_17;
wire n_23;
wire n_12;
wire n_20;
wire n_30;
wire n_19;
wire n_29;
wire n_25;

NAND3x1_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_4),
.C(n_1),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_9),
.B(n_1),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_7),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

OA21x2_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_0),
.B(n_2),
.Y(n_18)
);

OAI21x1_ASAP7_75t_L g19 ( 
.A1(n_15),
.A2(n_2),
.B(n_3),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_12),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_15),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_12),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_14),
.B1(n_18),
.B2(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

AOI222xp33_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_16),
.B1(n_11),
.B2(n_10),
.C1(n_19),
.C2(n_18),
.Y(n_25)
);

AOI221xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_22),
.B1(n_10),
.B2(n_18),
.C(n_4),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_18),
.B1(n_19),
.B2(n_3),
.Y(n_27)
);

NAND4xp25_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_18),
.C(n_6),
.D(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_18),
.B1(n_26),
.B2(n_29),
.Y(n_31)
);


endmodule