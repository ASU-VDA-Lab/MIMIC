module real_jpeg_33024_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_581, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_581;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_578;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_0),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_0),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_0),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_1),
.A2(n_88),
.B1(n_91),
.B2(n_93),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_1),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_1),
.A2(n_93),
.B1(n_324),
.B2(n_326),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_1),
.A2(n_93),
.B1(n_566),
.B2(n_570),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_2),
.A2(n_124),
.B(n_129),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_2),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_2),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_2),
.B(n_187),
.Y(n_472)
);

OAI22xp33_ASAP7_75t_SL g499 ( 
.A1(n_2),
.A2(n_81),
.B1(n_483),
.B2(n_500),
.Y(n_499)
);

OAI32xp33_ASAP7_75t_L g520 ( 
.A1(n_2),
.A2(n_162),
.A3(n_416),
.B1(n_521),
.B2(n_522),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_2),
.A2(n_158),
.B1(n_267),
.B2(n_318),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_3),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_4),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_4),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_4),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_5),
.B(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_5),
.A2(n_41),
.B1(n_240),
.B2(n_242),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_5),
.A2(n_41),
.B1(n_311),
.B2(n_315),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_SL g554 ( 
.A1(n_5),
.A2(n_41),
.B1(n_555),
.B2(n_556),
.Y(n_554)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_6),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_7),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_7),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_7),
.A2(n_148),
.B1(n_195),
.B2(n_198),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_7),
.A2(n_148),
.B1(n_213),
.B2(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_7),
.A2(n_148),
.B1(n_409),
.B2(n_411),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_8),
.A2(n_54),
.B1(n_57),
.B2(n_62),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_8),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_8),
.A2(n_62),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_8),
.A2(n_62),
.B1(n_230),
.B2(n_318),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_8),
.A2(n_62),
.B1(n_212),
.B2(n_367),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_9),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_9),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_9),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_10),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_12),
.A2(n_136),
.B1(n_139),
.B2(n_140),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_12),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_12),
.A2(n_139),
.B1(n_223),
.B2(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_12),
.A2(n_139),
.B1(n_441),
.B2(n_445),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_12),
.A2(n_139),
.B1(n_484),
.B2(n_489),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_13),
.A2(n_151),
.B1(n_152),
.B2(n_158),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_13),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_13),
.A2(n_151),
.B1(n_209),
.B2(n_212),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_13),
.A2(n_151),
.B1(n_350),
.B2(n_476),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_SL g492 ( 
.A1(n_13),
.A2(n_151),
.B1(n_277),
.B2(n_493),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_14),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_14),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_14),
.A2(n_77),
.B1(n_287),
.B2(n_292),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_14),
.A2(n_77),
.B1(n_356),
.B2(n_358),
.Y(n_355)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_15),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_16),
.A2(n_277),
.B1(n_280),
.B2(n_282),
.Y(n_276)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_16),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_16),
.A2(n_57),
.B1(n_282),
.B2(n_349),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_21),
.B(n_578),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_17),
.B(n_579),
.Y(n_578)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_18),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_19),
.A2(n_180),
.B1(n_181),
.B2(n_183),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_19),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_19),
.A2(n_180),
.B1(n_302),
.B2(n_305),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_19),
.A2(n_145),
.B1(n_180),
.B2(n_401),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_19),
.A2(n_180),
.B1(n_463),
.B2(n_466),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_543),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_389),
.B(n_538),
.Y(n_23)
);

NAND4xp25_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_268),
.C(n_371),
.D(n_382),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_244),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_26),
.B(n_244),
.Y(n_540)
);

XNOR2x1_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_189),
.Y(n_26)
);

XNOR2x1_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_97),
.Y(n_27)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_28),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_73),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_29),
.B(n_73),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_40),
.B1(n_53),
.B2(n_63),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_30),
.A2(n_53),
.B1(n_63),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_30),
.A2(n_63),
.B1(n_144),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_30),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_30),
.A2(n_63),
.B1(n_474),
.B2(n_475),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_30),
.B(n_267),
.Y(n_497)
);

AO21x1_ASAP7_75t_L g561 ( 
.A1(n_30),
.A2(n_63),
.B(n_348),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_31),
.Y(n_285)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AO21x2_ASAP7_75t_L g63 ( 
.A1(n_32),
.A2(n_64),
.B(n_69),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_32)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_33),
.Y(n_281)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_34),
.Y(n_261)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_35),
.Y(n_241)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_40),
.A2(n_63),
.B1(n_284),
.B2(n_286),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B(n_47),
.Y(n_40)
);

BUFx2_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_44),
.Y(n_439)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_48),
.Y(n_147)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_52),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_52),
.Y(n_403)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_52),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_56),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_60),
.Y(n_325)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_60),
.Y(n_351)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_61),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_63),
.A2(n_284),
.B1(n_286),
.B2(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_63),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_67),
.Y(n_173)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_68),
.Y(n_291)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_68),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_69),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_81),
.B1(n_87),
.B2(n_94),
.Y(n_73)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_74),
.Y(n_233)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_75),
.Y(n_450)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_76),
.Y(n_242)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_76),
.Y(n_488)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_81),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_81),
.A2(n_87),
.B1(n_274),
.B2(n_276),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_81),
.A2(n_462),
.B1(n_468),
.B2(n_470),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_81),
.A2(n_483),
.B1(n_492),
.B2(n_496),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

BUFx4f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_84),
.Y(n_412)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_86),
.Y(n_264)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_86),
.Y(n_279)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_86),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_86),
.Y(n_467)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_86),
.Y(n_491)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_95),
.Y(n_265)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g414 ( 
.A(n_96),
.Y(n_414)
);

INVx8_ASAP7_75t_L g496 ( 
.A(n_96),
.Y(n_496)
);

INVxp33_ASAP7_75t_L g385 ( 
.A(n_97),
.Y(n_385)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_142),
.C(n_149),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_99),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_123),
.B1(n_134),
.B2(n_135),
.Y(n_99)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_100),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_100),
.A2(n_134),
.B1(n_297),
.B2(n_301),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_100),
.A2(n_134),
.B1(n_208),
.B2(n_301),
.Y(n_336)
);

OAI22xp33_ASAP7_75t_L g376 ( 
.A1(n_100),
.A2(n_134),
.B1(n_208),
.B2(n_301),
.Y(n_376)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_101),
.A2(n_206),
.B1(n_298),
.B2(n_366),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_114),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_107),
.B1(n_109),
.B2(n_111),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_106),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_106),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_106),
.Y(n_304)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_106),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_108),
.Y(n_222)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_109),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

AOI22x1_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_117),
.B1(n_120),
.B2(n_122),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_118),
.Y(n_225)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_118),
.Y(n_423)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_124),
.Y(n_228)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AO21x1_ASAP7_75t_L g217 ( 
.A1(n_129),
.A2(n_218),
.B(n_226),
.Y(n_217)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_132),
.Y(n_558)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_134),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_134),
.B(n_267),
.Y(n_266)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_135),
.Y(n_204)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_142),
.A2(n_143),
.B1(n_149),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_149),
.Y(n_247)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_161),
.B1(n_179),
.B2(n_186),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_150),
.A2(n_161),
.B1(n_186),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_156),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_157),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_157),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_161),
.A2(n_179),
.B1(n_194),
.B2(n_200),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_161),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_161),
.A2(n_194),
.B1(n_200),
.B2(n_317),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_161),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_161),
.A2(n_200),
.B1(n_252),
.B2(n_525),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_161),
.A2(n_200),
.B1(n_564),
.B2(n_565),
.Y(n_563)
);

AO21x2_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_167),
.B(n_172),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g415 ( 
.A1(n_162),
.A2(n_416),
.B(n_422),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_163),
.Y(n_315)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_171),
.Y(n_314)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_171),
.Y(n_357)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_177),
.Y(n_172)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_SL g572 ( 
.A(n_182),
.Y(n_572)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AO22x2_ASAP7_75t_L g309 ( 
.A1(n_187),
.A2(n_310),
.B1(n_316),
.B2(n_319),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_187),
.A2(n_310),
.B1(n_355),
.B2(n_360),
.Y(n_354)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_189),
.B(n_384),
.C(n_385),
.Y(n_383)
);

XNOR2x1_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_216),
.Y(n_189)
);

OAI21x1_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_201),
.B(n_215),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_192),
.B(n_216),
.C(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_203),
.Y(n_215)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_197),
.Y(n_318)
);

INVx3_ASAP7_75t_SL g230 ( 
.A(n_198),
.Y(n_230)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_203),
.Y(n_378)
);

AOI22x1_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_205),
.A2(n_206),
.B1(n_366),
.B2(n_554),
.Y(n_553)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_231),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_217),
.A2(n_231),
.B1(n_232),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_223),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

NOR3xp33_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_227),
.C(n_229),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_239),
.B2(n_243),
.Y(n_232)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_235),
.B(n_267),
.Y(n_502)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_237),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_238),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_239),
.A2(n_243),
.B1(n_259),
.B2(n_265),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OA21x2_ASAP7_75t_L g329 ( 
.A1(n_243),
.A2(n_330),
.B(n_331),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_243),
.A2(n_259),
.B1(n_408),
.B2(n_413),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_243),
.A2(n_507),
.B1(n_508),
.B2(n_509),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.C(n_250),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_245),
.B(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_248),
.B(n_250),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_257),
.C(n_266),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_251),
.B(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_257),
.A2(n_258),
.B1(n_266),
.B2(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_266),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_267),
.B(n_417),
.Y(n_416)
);

NAND3xp33_ASAP7_75t_L g422 ( 
.A(n_267),
.B(n_423),
.C(n_424),
.Y(n_422)
);

OAI21xp33_ASAP7_75t_SL g434 ( 
.A1(n_267),
.A2(n_435),
.B(n_437),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_267),
.B(n_438),
.Y(n_437)
);

A2O1A1O1Ixp25_ASAP7_75t_L g538 ( 
.A1(n_268),
.A2(n_371),
.B(n_539),
.C(n_541),
.D(n_542),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_340),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_269),
.B(n_340),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_320),
.C(n_332),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_271),
.B(n_321),
.Y(n_381)
);

XNOR2x1_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_295),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_272),
.B(n_342),
.C(n_343),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_283),
.Y(n_272)
);

XOR2x2_ASAP7_75t_L g379 ( 
.A(n_273),
.B(n_283),
.Y(n_379)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_276),
.Y(n_331)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_278),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_280),
.Y(n_503)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_285),
.A2(n_347),
.B1(n_352),
.B2(n_353),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_285),
.A2(n_352),
.B1(n_400),
.B2(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_294),
.Y(n_436)
);

XNOR2x1_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_309),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_296),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_300),
.Y(n_299)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_302),
.Y(n_555)
);

INVx11_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx12f_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_309),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_328),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_322),
.B(n_329),
.Y(n_362)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_323),
.Y(n_353)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_327),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_328),
.A2(n_329),
.B1(n_364),
.B2(n_365),
.Y(n_363)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_329),
.A2(n_574),
.B1(n_575),
.B2(n_581),
.Y(n_573)
);

INVx5_ASAP7_75t_L g500 ( 
.A(n_330),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_332),
.B(n_381),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_335),
.C(n_337),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_334),
.B(n_375),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_335),
.A2(n_338),
.B1(n_339),
.B2(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_344),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_341),
.B(n_547),
.C(n_548),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_361),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_345),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_354),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_346),
.B(n_354),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_352),
.A2(n_434),
.B1(n_440),
.B2(n_446),
.Y(n_433)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_355),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_361),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_362),
.Y(n_574)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_365),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_380),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_372),
.B(n_380),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_377),
.C(n_379),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_388),
.Y(n_387)
);

XNOR2x1_ASAP7_75t_L g386 ( 
.A(n_377),
.B(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_379),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_386),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_383),
.B(n_386),
.C(n_540),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_427),
.B(n_537),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_393),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_391),
.B(n_393),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_398),
.C(n_404),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_394),
.A2(n_395),
.B1(n_531),
.B2(n_532),
.Y(n_530)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_398),
.A2(n_404),
.B1(n_405),
.B2(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_398),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_403),
.Y(n_476)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_415),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_406),
.A2(n_407),
.B1(n_415),
.B2(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_408),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_410),
.Y(n_458)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_423),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_424),
.Y(n_522)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_529),
.B(n_536),
.Y(n_427)
);

AOI21x1_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_515),
.B(n_528),
.Y(n_428)
);

OAI21x1_ASAP7_75t_SL g429 ( 
.A1(n_430),
.A2(n_479),
.B(n_514),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_460),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_431),
.B(n_460),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_447),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_432),
.A2(n_433),
.B1(n_447),
.B2(n_448),
.Y(n_512)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_437),
.Y(n_455)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_440),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx3_ASAP7_75t_SL g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_455),
.B1(n_456),
.B2(n_459),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_SL g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_471),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_461),
.B(n_473),
.C(n_477),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_462),
.Y(n_508)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_467),
.Y(n_495)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_472),
.A2(n_473),
.B1(n_477),
.B2(n_478),
.Y(n_471)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_472),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_473),
.Y(n_478)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_475),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_480),
.A2(n_505),
.B(n_513),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_481),
.A2(n_498),
.B(n_504),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_497),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_482),
.B(n_497),
.Y(n_504)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_492),
.Y(n_507)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_501),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_503),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_512),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_506),
.B(n_512),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_517),
.Y(n_515)
);

NOR2x1_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_517),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_523),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_518),
.B(n_526),
.C(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_526),
.Y(n_523)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_524),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_534),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_530),
.B(n_534),
.Y(n_536)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_576),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_546),
.B(n_549),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_546),
.B(n_549),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_550),
.B(n_573),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_551),
.B(n_552),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_553),
.B(n_559),
.Y(n_552)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx3_ASAP7_75t_SL g557 ( 
.A(n_558),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_560),
.A2(n_561),
.B1(n_562),
.B2(n_563),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);


endmodule