module real_jpeg_6936_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_1),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_1),
.B(n_181),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_1),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_1),
.B(n_248),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g296 ( 
.A(n_1),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_1),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_1),
.B(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_1),
.B(n_389),
.Y(n_388)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_2),
.B(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_2),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_2),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_2),
.B(n_239),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_3),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_3),
.Y(n_139)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_3),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_4),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_4),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_4),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_4),
.B(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_4),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_4),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_4),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_4),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_5),
.B(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_5),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_5),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_5),
.B(n_181),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_5),
.B(n_399),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_6),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_6),
.B(n_142),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_6),
.B(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_6),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_6),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_6),
.B(n_406),
.Y(n_405)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_8),
.Y(n_149)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_8),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_8),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_8),
.Y(n_391)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_9),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_9),
.Y(n_171)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_11),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_11),
.Y(n_152)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_11),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_11),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_11),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_12),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_12),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_12),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_12),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_12),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_12),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_12),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_13),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_13),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_13),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_13),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_13),
.B(n_363),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_13),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_13),
.B(n_412),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_14),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_14),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_15),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_15),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_15),
.B(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_15),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_15),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_15),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_15),
.B(n_309),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_15),
.B(n_62),
.Y(n_348)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_104),
.B(n_323),
.C(n_497),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_33),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_24),
.C(n_28),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_20),
.A2(n_28),
.B1(n_74),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_20),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_20),
.A2(n_85),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_20),
.B(n_228),
.Y(n_227)
);

NOR3xp33_ASAP7_75t_L g497 ( 
.A(n_20),
.B(n_44),
.C(n_100),
.Y(n_497)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_23),
.Y(n_203)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_23),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_24),
.A2(n_25),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_24),
.A2(n_25),
.B1(n_330),
.B2(n_336),
.Y(n_329)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_25),
.B(n_331),
.C(n_335),
.Y(n_478)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_27),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_28),
.A2(n_38),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_28),
.A2(n_74),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_28),
.B(n_147),
.C(n_151),
.Y(n_252)
);

OR2x2_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_31),
.Y(n_133)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_31),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_31),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_39),
.Y(n_38)
);

OR2x2_ASAP7_75t_SL g48 ( 
.A(n_32),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_32),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_94),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_80),
.C(n_81),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_35),
.B(n_494),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_60),
.C(n_71),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_36),
.B(n_485),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_51),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_56),
.C(n_58),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_44),
.C(n_47),
.Y(n_37)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_38),
.B(n_74),
.C(n_79),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_38),
.A2(n_75),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_38),
.B(n_115),
.C(n_118),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_38),
.A2(n_75),
.B1(n_473),
.B2(n_474),
.Y(n_472)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_41),
.Y(n_128)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx11_ASAP7_75t_L g217 ( 
.A(n_43),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_43),
.Y(n_251)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_43),
.Y(n_370)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_43),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_44),
.A2(n_97),
.B1(n_98),
.B2(n_102),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_44),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_44),
.A2(n_47),
.B1(n_48),
.B2(n_102),
.Y(n_474)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_47),
.A2(n_48),
.B1(n_129),
.B2(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_47),
.A2(n_48),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_48),
.B(n_125),
.C(n_129),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_48),
.B(n_193),
.C(n_323),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_49),
.B(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_49),
.Y(n_230)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_50),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_52),
.Y(n_58)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_55),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_56),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_60),
.B(n_71),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_63),
.C(n_67),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_61),
.A2(n_63),
.B1(n_64),
.B2(n_468),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_61),
.Y(n_468)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_63),
.A2(n_64),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_64),
.B(n_136),
.C(n_238),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_67),
.B(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_76),
.B2(n_79),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_76),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_76),
.A2(n_79),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_79),
.B(n_193),
.C(n_291),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_80),
.B(n_81),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_86),
.B1(n_87),
.B2(n_93),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_85),
.B(n_229),
.C(n_231),
.Y(n_286)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_90),
.C(n_93),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_103),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_99),
.A2(n_100),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_99),
.A2(n_100),
.B1(n_348),
.B2(n_349),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_99),
.B(n_344),
.C(n_349),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_100),
.B(n_308),
.C(n_311),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_492),
.B(n_496),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_460),
.B(n_489),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_350),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_280),
.B(n_313),
.C(n_314),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_253),
.B(n_279),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_109),
.B(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_221),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_110),
.B(n_221),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_172),
.C(n_204),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_111),
.B(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_143),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_112),
.B(n_144),
.C(n_153),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_124),
.C(n_134),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_113),
.B(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx8_ASAP7_75t_L g360 ( 
.A(n_123),
.Y(n_360)
);

BUFx5_ASAP7_75t_L g418 ( 
.A(n_123),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_124),
.A2(n_134),
.B1(n_135),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_124),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_125),
.B(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_127),
.B(n_168),
.Y(n_267)
);

INVx5_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_129),
.Y(n_262)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_133),
.Y(n_272)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_133),
.Y(n_310)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_136),
.A2(n_237),
.B1(n_238),
.B2(n_240),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_136),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_136),
.A2(n_140),
.B1(n_141),
.B2(n_240),
.Y(n_273)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_139),
.Y(n_386)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_139),
.Y(n_409)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_153),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_148),
.B(n_193),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_161),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_155),
.B(n_156),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_154),
.B(n_162),
.C(n_167),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_160),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_165),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_172),
.B(n_204),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_188),
.C(n_190),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_173),
.A2(n_188),
.B1(n_189),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_173),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_179),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_180),
.C(n_185),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_175),
.B(n_417),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_175),
.B(n_425),
.Y(n_424)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_178),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_184),
.B1(n_185),
.B2(n_187),
.Y(n_179)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_180),
.Y(n_187)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_184),
.A2(n_185),
.B1(n_295),
.B2(n_299),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_185),
.B(n_238),
.C(n_296),
.Y(n_345)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_190),
.B(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_197),
.C(n_200),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_191),
.A2(n_192),
.B1(n_447),
.B2(n_448),
.Y(n_446)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_193),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_193),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_193),
.A2(n_288),
.B1(n_323),
.B2(n_326),
.Y(n_322)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_196),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_448)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_220),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_207),
.C(n_220),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_214),
.C(n_218),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_214),
.A2(n_331),
.B1(n_334),
.B2(n_335),
.Y(n_330)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_214),
.Y(n_335)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_217),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_222),
.B(n_224),
.C(n_241),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_241),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_234),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_226),
.B(n_227),
.C(n_234),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_237),
.A2(n_238),
.B1(n_296),
.B2(n_298),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_237),
.A2(n_238),
.B1(n_358),
.B2(n_359),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_238),
.B(n_358),
.Y(n_357)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_239),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_242),
.B(n_244),
.C(n_245),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_252),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_247),
.B(n_249),
.C(n_304),
.Y(n_303)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_252),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_277),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_254),
.B(n_277),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_259),
.C(n_274),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_255),
.A2(n_256),
.B1(n_452),
.B2(n_453),
.Y(n_451)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_259),
.B(n_274),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.C(n_273),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_260),
.B(n_442),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_263),
.B(n_273),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.C(n_268),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_264),
.A2(n_265),
.B1(n_268),
.B2(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_267),
.B(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_268),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_269),
.B(n_368),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_269),
.B(n_420),
.Y(n_419)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_281),
.B(n_315),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_283),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_316),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g459 ( 
.A(n_283),
.B(n_316),
.Y(n_459)
);

FAx1_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_300),
.CI(n_312),
.CON(n_283),
.SN(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_294),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_286),
.B(n_287),
.C(n_294),
.Y(n_339)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_295),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_296),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_303),
.C(n_305),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_311),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_317),
.B(n_319),
.C(n_337),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_337),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_327),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_320),
.B(n_328),
.C(n_329),
.Y(n_469)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_323),
.Y(n_326)
);

INVx8_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_330),
.Y(n_336)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_331),
.Y(n_334)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_338),
.B(n_342),
.C(n_343),
.Y(n_479)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

AO22x1_ASAP7_75t_SL g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_346),
.B2(n_347),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_348),
.Y(n_349)
);

OAI31xp33_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_456),
.A3(n_457),
.B(n_459),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_450),
.B(n_455),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_353),
.A2(n_437),
.B(n_449),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_393),
.B(n_436),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_378),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_355),
.B(n_378),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_365),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_356),
.B(n_366),
.C(n_375),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_357),
.B(n_361),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_357),
.B(n_362),
.C(n_364),
.Y(n_445)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_375),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_371),
.C(n_373),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_367),
.B(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_371),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_380)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_381),
.C(n_392),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_379),
.B(n_433),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_381),
.A2(n_382),
.B1(n_392),
.B2(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_387),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_383),
.A2(n_384),
.B1(n_387),
.B2(n_388),
.Y(n_402)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_392),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_430),
.B(n_435),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_414),
.B(n_429),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_403),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_396),
.B(n_403),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_402),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_398),
.B(n_400),
.C(n_402),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_410),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_404),
.A2(n_405),
.B1(n_410),
.B2(n_411),
.Y(n_427)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx6_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx8_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_423),
.B(n_428),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_419),
.Y(n_415)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_421),
.Y(n_420)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_427),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_424),
.B(n_427),
.Y(n_428)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_432),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_431),
.B(n_432),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_438),
.B(n_439),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_440),
.A2(n_441),
.B1(n_443),
.B2(n_444),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_440),
.B(n_445),
.C(n_446),
.Y(n_454)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_454),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_451),
.B(n_454),
.Y(n_455)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_452),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_486),
.Y(n_460)
);

OAI21xp33_ASAP7_75t_L g489 ( 
.A1(n_461),
.A2(n_490),
.B(n_491),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_480),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_462),
.B(n_480),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_470),
.C(n_479),
.Y(n_462)
);

FAx1_ASAP7_75t_SL g488 ( 
.A(n_463),
.B(n_470),
.CI(n_479),
.CON(n_488),
.SN(n_488)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_469),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_466),
.C(n_469),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_472),
.B1(n_475),
.B2(n_476),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_477),
.C(n_478),
.Y(n_483)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_482),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_481),
.B(n_483),
.C(n_484),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_487),
.B(n_488),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g498 ( 
.A(n_488),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_495),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_493),
.B(n_495),
.Y(n_496)
);


endmodule