module fake_jpeg_20551_n_336 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_18),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_19),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_20),
.B1(n_33),
.B2(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_58),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_20),
.B1(n_33),
.B2(n_26),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_65),
.B1(n_36),
.B2(n_25),
.Y(n_73)
);

NAND2x1_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_17),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_53),
.B(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_20),
.B1(n_26),
.B2(n_32),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_23),
.B1(n_32),
.B2(n_25),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_67),
.B1(n_25),
.B2(n_27),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_32),
.B1(n_23),
.B2(n_26),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_SL g117 ( 
.A1(n_73),
.A2(n_76),
.B(n_48),
.Y(n_117)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_77),
.B(n_39),
.Y(n_112)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_82),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_71),
.Y(n_119)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_98),
.B(n_121),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_53),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_100),
.A2(n_109),
.B(n_114),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_68),
.C(n_53),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_124),
.C(n_37),
.Y(n_144)
);

MAJx2_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_84),
.C(n_72),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_125),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_108),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_59),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_119),
.Y(n_135)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_59),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_116),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_36),
.B1(n_55),
.B2(n_61),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_58),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_81),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_37),
.C(n_39),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_27),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_94),
.B1(n_79),
.B2(n_75),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_128),
.A2(n_147),
.B1(n_106),
.B2(n_123),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_78),
.B(n_80),
.C(n_55),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_148),
.B(n_110),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_61),
.B1(n_69),
.B2(n_49),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_138),
.B1(n_140),
.B2(n_142),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_88),
.B1(n_74),
.B2(n_96),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_88),
.B1(n_92),
.B2(n_36),
.Y(n_140)
);

OAI32xp33_ASAP7_75t_L g141 ( 
.A1(n_102),
.A2(n_52),
.A3(n_27),
.B1(n_28),
.B2(n_17),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_116),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_109),
.B1(n_100),
.B2(n_125),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_17),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_30),
.B1(n_29),
.B2(n_22),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_153),
.C(n_30),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_114),
.B1(n_104),
.B2(n_107),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_31),
.Y(n_148)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_98),
.A2(n_52),
.B1(n_42),
.B2(n_51),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_152),
.B1(n_97),
.B2(n_17),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_28),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_31),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_99),
.A2(n_52),
.B1(n_42),
.B2(n_51),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_45),
.C(n_39),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_154),
.Y(n_204)
);

AO21x1_ASAP7_75t_L g195 ( 
.A1(n_155),
.A2(n_158),
.B(n_151),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_156),
.A2(n_169),
.B1(n_140),
.B2(n_145),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_135),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_161),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_126),
.A2(n_122),
.B(n_28),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_160),
.B(n_176),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_97),
.B(n_123),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_149),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_163),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_134),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_164),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_137),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_166),
.Y(n_191)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_106),
.Y(n_168)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_139),
.A2(n_111),
.B1(n_107),
.B2(n_118),
.Y(n_169)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_170),
.B(n_173),
.CI(n_150),
.CON(n_190),
.SN(n_190)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_132),
.B(n_111),
.Y(n_173)
);

OAI211xp5_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_17),
.B(n_118),
.C(n_29),
.Y(n_174)
);

OAI31xp33_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_129),
.A3(n_143),
.B(n_152),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_181),
.B1(n_171),
.B2(n_153),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_17),
.B(n_1),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_30),
.Y(n_208)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_133),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_181),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_182),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_187),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_136),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_186),
.B(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_180),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_179),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_193),
.A2(n_205),
.B1(n_166),
.B2(n_164),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_195),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_144),
.C(n_148),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_203),
.C(n_155),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_158),
.B(n_136),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_208),
.Y(n_218)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_202),
.B1(n_207),
.B2(n_210),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_139),
.B1(n_132),
.B2(n_146),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_148),
.C(n_146),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_172),
.A2(n_145),
.B1(n_29),
.B2(n_22),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_29),
.B1(n_22),
.B2(n_21),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_204),
.B(n_173),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_211),
.B(n_220),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_197),
.B(n_159),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_222),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_216),
.C(n_224),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_192),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_217),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_161),
.B(n_154),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_215),
.A2(n_228),
.B(n_234),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_162),
.C(n_163),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_189),
.A2(n_176),
.B1(n_174),
.B2(n_157),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_191),
.B(n_184),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_175),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_223),
.A2(n_206),
.B1(n_207),
.B2(n_193),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_182),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_236),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_194),
.A2(n_182),
.B(n_178),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_192),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_189),
.A2(n_182),
.B1(n_178),
.B2(n_165),
.Y(n_230)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_198),
.B1(n_206),
.B2(n_185),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_188),
.A2(n_167),
.B(n_10),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_188),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_237),
.A2(n_213),
.B1(n_225),
.B2(n_212),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_238),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_229),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_242),
.Y(n_261)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_226),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_254),
.B1(n_256),
.B2(n_219),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_205),
.B(n_190),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_221),
.Y(n_253)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_224),
.A2(n_208),
.B1(n_190),
.B2(n_201),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_216),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_222),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_22),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_218),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_251),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_270),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_264),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_220),
.Y(n_263)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_239),
.B(n_236),
.Y(n_264)
);

XOR2x1_ASAP7_75t_SL g266 ( 
.A(n_237),
.B(n_217),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_267),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_268),
.B(n_269),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_228),
.B(n_9),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_21),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_21),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_277),
.C(n_256),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_248),
.B(n_21),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_245),
.Y(n_279)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_271),
.A2(n_246),
.B1(n_259),
.B2(n_250),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_286),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_244),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_247),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_248),
.C(n_267),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_293),
.C(n_284),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_243),
.B1(n_266),
.B2(n_275),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_288),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_247),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_290),
.Y(n_306)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_238),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_265),
.A2(n_258),
.B(n_254),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_262),
.C(n_264),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_244),
.C(n_258),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_294),
.B(n_296),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_299),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_302),
.B(n_292),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_270),
.B1(n_9),
.B2(n_10),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_15),
.C(n_14),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_294),
.C(n_297),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_15),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_13),
.C(n_12),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_304),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g305 ( 
.A(n_280),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_305),
.B(n_283),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_309),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_281),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_302),
.A2(n_282),
.B1(n_283),
.B2(n_278),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_11),
.B1(n_8),
.B2(n_3),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_314),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_298),
.A2(n_306),
.B(n_278),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_313),
.A2(n_316),
.B1(n_8),
.B2(n_2),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_12),
.Y(n_316)
);

AND2x2_ASAP7_75t_SL g317 ( 
.A(n_308),
.B(n_314),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_318),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_319),
.A2(n_0),
.B(n_3),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_316),
.B(n_11),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_L g325 ( 
.A1(n_320),
.A2(n_307),
.B(n_2),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_324),
.C(n_4),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_0),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_327),
.Y(n_331)
);

NAND4xp25_ASAP7_75t_SL g328 ( 
.A(n_317),
.B(n_0),
.C(n_3),
.D(n_4),
.Y(n_328)
);

O2A1O1Ixp33_ASAP7_75t_SL g330 ( 
.A1(n_328),
.A2(n_329),
.B(n_321),
.C(n_5),
.Y(n_330)
);

O2A1O1Ixp33_ASAP7_75t_SL g332 ( 
.A1(n_330),
.A2(n_326),
.B(n_5),
.C(n_6),
.Y(n_332)
);

A2O1A1O1Ixp25_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_331),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_4),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g335 ( 
.A(n_334),
.B(n_4),
.CI(n_323),
.CON(n_335),
.SN(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_321),
.Y(n_336)
);


endmodule