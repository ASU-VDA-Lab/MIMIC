module fake_jpeg_30445_n_515 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_515);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_515;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_361;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_20),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_53),
.B(n_98),
.Y(n_116)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_54),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_74),
.Y(n_115)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_28),
.B(n_6),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_57),
.B(n_60),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_6),
.Y(n_60)
);

BUFx6f_ASAP7_75t_SL g61 ( 
.A(n_19),
.Y(n_61)
);

INVxp67_ASAP7_75t_SL g136 ( 
.A(n_61),
.Y(n_136)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_8),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_65),
.B(n_71),
.Y(n_129)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_17),
.B(n_0),
.Y(n_70)
);

NAND2x1_ASAP7_75t_SL g149 ( 
.A(n_70),
.B(n_36),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_16),
.B(n_8),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_16),
.B(n_8),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_75),
.B(n_82),
.Y(n_148)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_19),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_23),
.B(n_5),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_83),
.B(n_90),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_19),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_85),
.B(n_97),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_18),
.A2(n_15),
.B(n_1),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_36),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_23),
.B(n_5),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_29),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_34),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_100),
.B(n_121),
.Y(n_176)
);

INVx6_ASAP7_75t_SL g107 ( 
.A(n_61),
.Y(n_107)
);

CKINVDCx9p33_ASAP7_75t_R g204 ( 
.A(n_107),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_113),
.B(n_125),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_70),
.A2(n_17),
.B1(n_44),
.B2(n_36),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_117),
.A2(n_54),
.B1(n_59),
.B2(n_50),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_78),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_89),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_99),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_146),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_131),
.B(n_152),
.Y(n_199)
);

BUFx4f_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

NOR4xp25_ASAP7_75t_SL g146 ( 
.A(n_53),
.B(n_9),
.C(n_1),
.D(n_3),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_85),
.B(n_44),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_80),
.B(n_34),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_155),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_96),
.B(n_40),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_40),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_82),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_50),
.Y(n_207)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_158),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_160),
.B(n_197),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_115),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_161),
.B(n_165),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g217 ( 
.A(n_162),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

INVx3_ASAP7_75t_SL g219 ( 
.A(n_163),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_164),
.A2(n_180),
.B1(n_200),
.B2(n_202),
.Y(n_242)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_167),
.Y(n_221)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

CKINVDCx12_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_169),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_122),
.A2(n_33),
.B1(n_47),
.B2(n_88),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_174),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_147),
.A2(n_33),
.B1(n_47),
.B2(n_58),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_39),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_187),
.Y(n_209)
);

BUFx4f_ASAP7_75t_SL g182 ( 
.A(n_112),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_182),
.B(n_190),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_183),
.Y(n_245)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_185),
.Y(n_235)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_39),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_137),
.B(n_38),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_203),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_118),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_62),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_191),
.B(n_195),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_130),
.Y(n_192)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_119),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_110),
.Y(n_196)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_198),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_117),
.A2(n_84),
.B1(n_93),
.B2(n_67),
.Y(n_200)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_110),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_201),
.A2(n_109),
.B1(n_112),
.B2(n_111),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_105),
.A2(n_47),
.B1(n_63),
.B2(n_64),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_116),
.B(n_38),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_129),
.B(n_46),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_207),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_133),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_206),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_160),
.B(n_114),
.C(n_129),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_213),
.B(n_223),
.C(n_227),
.Y(n_284)
);

AO21x2_ASAP7_75t_L g214 ( 
.A1(n_204),
.A2(n_150),
.B(n_105),
.Y(n_214)
);

OA22x2_ASAP7_75t_L g275 ( 
.A1(n_214),
.A2(n_197),
.B1(n_185),
.B2(n_201),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_114),
.C(n_133),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_113),
.C(n_123),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_172),
.A2(n_95),
.B1(n_86),
.B2(n_72),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_237),
.A2(n_243),
.B1(n_244),
.B2(n_246),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_181),
.A2(n_69),
.B1(n_87),
.B2(n_73),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_203),
.A2(n_51),
.B1(n_150),
.B2(n_142),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_205),
.A2(n_157),
.B1(n_142),
.B2(n_132),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_158),
.B(n_123),
.C(n_91),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_247),
.B(n_179),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_184),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_248),
.B(n_249),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_165),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_251),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_241),
.A2(n_206),
.B1(n_204),
.B2(n_109),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_252),
.A2(n_196),
.B1(n_233),
.B2(n_245),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_253),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_176),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_254),
.B(n_276),
.Y(n_309)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_255),
.Y(n_293)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_256),
.Y(n_290)
);

AND2x6_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_199),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_259),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_231),
.Y(n_258)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_258),
.Y(n_297)
);

AND2x6_ASAP7_75t_L g259 ( 
.A(n_213),
.B(n_223),
.Y(n_259)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_218),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_260),
.Y(n_304)
);

OR2x2_ASAP7_75t_SL g261 ( 
.A(n_209),
.B(n_224),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g316 ( 
.A(n_261),
.B(n_279),
.CI(n_94),
.CON(n_316),
.SN(n_316)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_234),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_262),
.B(n_269),
.Y(n_303)
);

AND2x6_ASAP7_75t_L g263 ( 
.A(n_208),
.B(n_56),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_271),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_241),
.A2(n_166),
.B(n_175),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_264),
.A2(n_265),
.B(n_215),
.Y(n_288)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_212),
.Y(n_266)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_266),
.Y(n_299)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_210),
.Y(n_268)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_268),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_224),
.B(n_198),
.Y(n_269)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_218),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_270),
.Y(n_305)
);

INVx13_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_242),
.A2(n_171),
.B1(n_132),
.B2(n_130),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_291)
);

NOR3xp33_ASAP7_75t_L g273 ( 
.A(n_209),
.B(n_167),
.C(n_46),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_273),
.B(n_274),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_222),
.B(n_168),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_275),
.A2(n_214),
.B1(n_215),
.B2(n_235),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_227),
.B(n_173),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_222),
.B(n_159),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_277),
.B(n_282),
.Y(n_311)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_210),
.Y(n_278)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_278),
.Y(n_301)
);

NAND2x1p5_ASAP7_75t_L g279 ( 
.A(n_214),
.B(n_76),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_225),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_283),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_244),
.A2(n_157),
.B1(n_159),
.B2(n_188),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_217),
.B1(n_219),
.B2(n_238),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_186),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_239),
.B(n_182),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_237),
.C(n_226),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_259),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_249),
.B(n_246),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_286),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_288),
.B(n_248),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_291),
.A2(n_292),
.B1(n_302),
.B2(n_281),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_267),
.A2(n_214),
.B1(n_243),
.B2(n_228),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_296),
.A2(n_310),
.B1(n_255),
.B2(n_253),
.Y(n_344)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_251),
.Y(n_308)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_308),
.Y(n_342)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_256),
.Y(n_312)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_312),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_254),
.A2(n_214),
.B(n_182),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_313),
.A2(n_264),
.B(n_250),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_240),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_314),
.B(n_316),
.Y(n_334)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_266),
.Y(n_315)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_315),
.Y(n_347)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_268),
.Y(n_317)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_278),
.Y(n_318)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_318),
.Y(n_329)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_258),
.Y(n_319)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_319),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_303),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_320),
.B(n_321),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_306),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_322),
.A2(n_325),
.B(n_336),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_284),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_323),
.B(n_350),
.C(n_297),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_311),
.A2(n_267),
.B1(n_272),
.B2(n_282),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_324),
.A2(n_233),
.B1(n_235),
.B2(n_178),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_316),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_326),
.B(n_135),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_289),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_328),
.B(n_335),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_330),
.A2(n_331),
.B1(n_341),
.B2(n_296),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_302),
.A2(n_265),
.B1(n_276),
.B2(n_250),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_333),
.B(n_280),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_295),
.B(n_262),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_313),
.A2(n_279),
.B(n_275),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_289),
.Y(n_337)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_337),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_286),
.B(n_314),
.Y(n_338)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_338),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_309),
.B(n_257),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_340),
.B(n_353),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_292),
.A2(n_279),
.B1(n_275),
.B2(n_263),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_344),
.A2(n_304),
.B1(n_305),
.B2(n_298),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_311),
.B(n_275),
.Y(n_345)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_345),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_298),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_346),
.Y(n_354)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_290),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_349),
.Y(n_362)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_290),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_287),
.B(n_285),
.C(n_288),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_308),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_299),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_295),
.B(n_307),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_211),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_316),
.B(n_261),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_333),
.B(n_294),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_355),
.B(n_373),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_339),
.A2(n_291),
.B1(n_312),
.B2(n_319),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_356),
.A2(n_361),
.B1(n_370),
.B2(n_386),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_322),
.A2(n_304),
.B(n_305),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_358),
.A2(n_104),
.B(n_270),
.Y(n_400)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_363),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_365),
.A2(n_366),
.B1(n_369),
.B2(n_374),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_345),
.A2(n_299),
.B1(n_315),
.B2(n_317),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_381),
.C(n_347),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_368),
.B(n_342),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_331),
.A2(n_318),
.B1(n_301),
.B2(n_300),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_326),
.A2(n_293),
.B1(n_297),
.B2(n_300),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_338),
.B(n_301),
.Y(n_371)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_371),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_334),
.B(n_293),
.Y(n_372)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_372),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_323),
.B(n_240),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_330),
.A2(n_341),
.B1(n_350),
.B2(n_334),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_332),
.Y(n_375)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_375),
.Y(n_414)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_379),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_340),
.B(n_221),
.Y(n_380)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_380),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_211),
.C(n_221),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_324),
.B(n_271),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_382),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_336),
.B(n_332),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_383),
.B(n_343),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_337),
.A2(n_351),
.B1(n_349),
.B2(n_348),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_384),
.A2(n_163),
.B1(n_162),
.B2(n_170),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_385),
.A2(n_141),
.B(n_144),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_387),
.B(n_388),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_394),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_367),
.B(n_329),
.C(n_327),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_393),
.B(n_401),
.C(n_405),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_329),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_346),
.Y(n_395)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_395),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_364),
.B(n_327),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_410),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_398),
.A2(n_377),
.B1(n_356),
.B2(n_354),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_400),
.A2(n_402),
.B(n_358),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_135),
.C(n_111),
.Y(n_401)
);

OAI21xp33_ASAP7_75t_L g402 ( 
.A1(n_371),
.A2(n_177),
.B(n_144),
.Y(n_402)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_403),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_368),
.B(n_101),
.C(n_141),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_364),
.B(n_104),
.C(n_68),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_412),
.C(n_365),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_359),
.B(n_271),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_376),
.B(n_43),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_411),
.B(n_363),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_381),
.B(n_192),
.C(n_183),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_386),
.A2(n_43),
.B1(n_30),
.B2(n_29),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_413),
.A2(n_385),
.B1(n_30),
.B2(n_366),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_393),
.B(n_357),
.Y(n_415)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_415),
.Y(n_444)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_418),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_260),
.Y(n_445)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_421),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_392),
.B(n_374),
.C(n_383),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_430),
.C(n_431),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_391),
.A2(n_359),
.B(n_400),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_425),
.A2(n_387),
.B(n_396),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_407),
.B(n_369),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_426),
.B(n_434),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_399),
.A2(n_372),
.B1(n_357),
.B2(n_360),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_427),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_406),
.A2(n_360),
.B1(n_389),
.B2(n_390),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_428),
.A2(n_429),
.B1(n_402),
.B2(n_409),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_407),
.B(n_394),
.C(n_397),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_412),
.B(n_385),
.C(n_362),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_414),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_433),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_410),
.B(n_362),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_435),
.B(n_408),
.Y(n_441)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_404),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_436),
.B(n_10),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_384),
.C(n_270),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_437),
.B(n_260),
.C(n_35),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_438),
.A2(n_11),
.B(n_4),
.Y(n_473)
);

BUFx12_ASAP7_75t_L g439 ( 
.A(n_425),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_451),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_440),
.B(n_441),
.Y(n_460)
);

NOR3xp33_ASAP7_75t_SL g443 ( 
.A(n_418),
.B(n_405),
.C(n_388),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_443),
.A2(n_42),
.B1(n_26),
.B2(n_5),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_454),
.C(n_424),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_447),
.B(n_42),
.Y(n_470)
);

FAx1_ASAP7_75t_L g449 ( 
.A(n_434),
.B(n_138),
.CI(n_140),
.CON(n_449),
.SN(n_449)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_449),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_428),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_453),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_423),
.B(n_35),
.C(n_140),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_419),
.A2(n_138),
.B(n_64),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_456),
.A2(n_11),
.B(n_1),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_446),
.A2(n_426),
.B1(n_432),
.B2(n_424),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_457),
.A2(n_471),
.B1(n_450),
.B2(n_449),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_455),
.A2(n_417),
.B1(n_437),
.B2(n_420),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_458),
.B(n_459),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_444),
.A2(n_431),
.B1(n_419),
.B2(n_430),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_463),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_422),
.C(n_416),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_462),
.B(n_442),
.C(n_448),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_448),
.B(n_416),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_452),
.A2(n_422),
.B1(n_63),
.B2(n_177),
.Y(n_466)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_466),
.Y(n_480)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_467),
.Y(n_485)
);

OA21x2_ASAP7_75t_L g468 ( 
.A1(n_439),
.A2(n_136),
.B(n_4),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_469),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_470),
.B(n_473),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_450),
.A2(n_15),
.B1(n_4),
.B2(n_5),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_451),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_476),
.B(n_477),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_439),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_483),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_461),
.B(n_442),
.C(n_454),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_479),
.B(n_484),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_464),
.A2(n_443),
.B(n_449),
.Y(n_481)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_481),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_447),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_462),
.B(n_50),
.C(n_45),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_487),
.B(n_468),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_481),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_491),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_486),
.A2(n_464),
.B(n_468),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_490),
.A2(n_494),
.B(n_496),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_477),
.B(n_457),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_493),
.B(n_482),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_479),
.A2(n_473),
.B(n_463),
.Y(n_494)
);

BUFx24_ASAP7_75t_SL g496 ( 
.A(n_474),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_501),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_492),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_474),
.C(n_495),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_45),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_497),
.B(n_487),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_503),
.Y(n_507)
);

AOI322xp5_ASAP7_75t_L g504 ( 
.A1(n_488),
.A2(n_480),
.A3(n_482),
.B1(n_475),
.B2(n_485),
.C1(n_470),
.C2(n_50),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_504),
.A2(n_136),
.B(n_26),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_508),
.Y(n_510)
);

HAxp5_ASAP7_75t_SL g509 ( 
.A(n_505),
.B(n_499),
.CON(n_509),
.SN(n_509)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_509),
.A2(n_500),
.B(n_507),
.Y(n_511)
);

AOI322xp5_ASAP7_75t_L g512 ( 
.A1(n_511),
.A2(n_510),
.A3(n_504),
.B1(n_4),
.B2(n_9),
.C1(n_10),
.C2(n_42),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_512),
.A2(n_9),
.B(n_0),
.Y(n_513)
);

BUFx24_ASAP7_75t_SL g514 ( 
.A(n_513),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_26),
.C(n_0),
.Y(n_515)
);


endmodule