module fake_jpeg_23784_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_4),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx16f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx10_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_5),
.B(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_1),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_13),
.B(n_15),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_7),
.Y(n_15)
);

NOR3xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_2),
.C(n_7),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_14),
.A2(n_10),
.B1(n_12),
.B2(n_11),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_19),
.B(n_9),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_24),
.Y(n_28)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_11),
.Y(n_25)
);

BUFx24_ASAP7_75t_SL g27 ( 
.A(n_25),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_27),
.B(n_20),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_31),
.B1(n_10),
.B2(n_12),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_34),
.B(n_35),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_13),
.B(n_8),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_19),
.C(n_8),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_9),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_38),
.B(n_2),
.Y(n_39)
);


endmodule