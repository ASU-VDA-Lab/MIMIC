module fake_jpeg_13859_n_565 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_565);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_565;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_12),
.B(n_13),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_62),
.B(n_64),
.Y(n_175)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_16),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_66),
.Y(n_161)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_68),
.Y(n_191)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_69),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_70),
.Y(n_158)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_71),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_73),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_74),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_33),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_75),
.B(n_83),
.Y(n_131)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_78),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_79),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_30),
.B(n_1),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_33),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_96),
.Y(n_133)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_86),
.Y(n_182)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_89),
.Y(n_183)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_90),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_91),
.Y(n_206)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g196 ( 
.A(n_92),
.Y(n_196)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_93),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_27),
.B(n_1),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_94),
.B(n_95),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_27),
.B(n_1),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_45),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_29),
.B(n_15),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_99),
.B(n_109),
.Y(n_150)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_101),
.Y(n_207)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

BUFx10_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_57),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_103),
.B(n_108),
.Y(n_163)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

INVx6_ASAP7_75t_SL g108 ( 
.A(n_57),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_29),
.B(n_43),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_20),
.Y(n_110)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_110),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

INVx3_ASAP7_75t_SL g112 ( 
.A(n_36),
.Y(n_112)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_47),
.B(n_3),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_115),
.B(n_117),
.Y(n_171)
);

BUFx8_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_46),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_19),
.Y(n_118)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_118),
.Y(n_208)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_121),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_120),
.B(n_122),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_19),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_126),
.Y(n_155)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_20),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_124),
.B(n_125),
.Y(n_186)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_23),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_62),
.A2(n_32),
.B1(n_31),
.B2(n_43),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_129),
.A2(n_187),
.B1(n_192),
.B2(n_198),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_61),
.A2(n_32),
.B1(n_31),
.B2(n_53),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_130),
.A2(n_134),
.B1(n_136),
.B2(n_139),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_25),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_132),
.B(n_204),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_65),
.A2(n_70),
.B1(n_121),
.B2(n_72),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_74),
.A2(n_39),
.B1(n_41),
.B2(n_46),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_74),
.A2(n_41),
.B1(n_39),
.B2(n_51),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_41),
.B1(n_39),
.B2(n_51),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_144),
.A2(n_152),
.B1(n_157),
.B2(n_165),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_85),
.A2(n_51),
.B1(n_32),
.B2(n_55),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_73),
.A2(n_55),
.B1(n_23),
.B2(n_25),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_113),
.A2(n_51),
.B1(n_49),
.B2(n_44),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_90),
.A2(n_49),
.B1(n_44),
.B2(n_40),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_167),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_64),
.B(n_40),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_170),
.B(n_190),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_123),
.A2(n_126),
.B1(n_100),
.B2(n_120),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_89),
.A2(n_38),
.B1(n_54),
.B2(n_48),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_102),
.A2(n_38),
.B1(n_54),
.B2(n_5),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_115),
.A2(n_54),
.B1(n_4),
.B2(n_5),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_83),
.B(n_3),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_79),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_104),
.B(n_6),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_193),
.B(n_205),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_107),
.B(n_6),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_194),
.B(n_201),
.Y(n_266)
);

OA22x2_ASAP7_75t_L g197 ( 
.A1(n_80),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_197)
);

OA21x2_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_12),
.B(n_156),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_91),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_107),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_199),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_110),
.B(n_10),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_116),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_110),
.B(n_10),
.Y(n_205)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

BUFx2_ASAP7_75t_SL g327 ( 
.A(n_209),
.Y(n_327)
);

INVx11_ASAP7_75t_L g210 ( 
.A(n_137),
.Y(n_210)
);

INVx11_ASAP7_75t_L g298 ( 
.A(n_210),
.Y(n_298)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_211),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_134),
.A2(n_101),
.B1(n_105),
.B2(n_111),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_213),
.A2(n_263),
.B1(n_254),
.B2(n_271),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_195),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_215),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_217),
.Y(n_289)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_138),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_218),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_219),
.A2(n_241),
.B1(n_242),
.B2(n_252),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_145),
.Y(n_220)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_135),
.Y(n_221)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_221),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_171),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_222),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_131),
.B(n_175),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_223),
.B(n_234),
.Y(n_283)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_145),
.Y(n_224)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_224),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_147),
.B(n_150),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_225),
.B(n_227),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_185),
.A2(n_203),
.B1(n_191),
.B2(n_178),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_226),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_132),
.A2(n_133),
.B(n_172),
.C(n_197),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_168),
.Y(n_228)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_228),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_163),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_229),
.B(n_236),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_143),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_230),
.B(n_240),
.Y(n_316)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_140),
.Y(n_231)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_231),
.Y(n_280)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_146),
.Y(n_232)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_142),
.Y(n_233)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_233),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_156),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_160),
.Y(n_235)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_235),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_196),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_151),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_153),
.B(n_155),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_L g241 ( 
.A1(n_152),
.A2(n_177),
.B1(n_144),
.B2(n_167),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_157),
.A2(n_139),
.B1(n_136),
.B2(n_165),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_178),
.B(n_151),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_243),
.B(n_251),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_166),
.B(n_184),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_244),
.B(n_246),
.C(n_247),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_196),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_245),
.B(n_259),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_149),
.B(n_161),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_164),
.B(n_182),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_174),
.Y(n_248)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_248),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_154),
.Y(n_250)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_250),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_197),
.B(n_180),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_199),
.A2(n_181),
.B1(n_159),
.B2(n_189),
.Y(n_252)
);

BUFx6f_ASAP7_75t_SL g253 ( 
.A(n_137),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_253),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_127),
.A2(n_207),
.B1(n_206),
.B2(n_173),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_254),
.A2(n_261),
.B(n_268),
.Y(n_325)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_174),
.Y(n_255)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_255),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_173),
.Y(n_256)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_176),
.Y(n_257)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_257),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_179),
.B(n_188),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_258),
.B(n_262),
.Y(n_313)
);

BUFx4f_ASAP7_75t_SL g259 ( 
.A(n_137),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_127),
.Y(n_260)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_260),
.Y(n_328)
);

NAND2xp33_ASAP7_75t_SL g261 ( 
.A(n_179),
.B(n_188),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_196),
.B(n_128),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_189),
.A2(n_141),
.B1(n_159),
.B2(n_169),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_128),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_148),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_265),
.B(n_269),
.Y(n_317)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_141),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_267),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_148),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_268),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_154),
.B(n_158),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_158),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_270),
.Y(n_301)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_162),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_271),
.B(n_274),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_162),
.B(n_208),
.C(n_143),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_273),
.B(n_246),
.C(n_247),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_169),
.B(n_131),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_138),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_275),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_133),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_277),
.Y(n_314)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_135),
.Y(n_278)
);

NAND2x1_ASAP7_75t_SL g305 ( 
.A(n_278),
.B(n_279),
.Y(n_305)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_135),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_249),
.A2(n_251),
.B1(n_240),
.B2(n_216),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_287),
.A2(n_332),
.B1(n_321),
.B2(n_300),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_242),
.A2(n_252),
.B1(n_241),
.B2(n_238),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_295),
.Y(n_353)
);

AND2x2_ASAP7_75t_SL g300 ( 
.A(n_230),
.B(n_273),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_300),
.B(n_325),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_212),
.A2(n_219),
.B1(n_249),
.B2(n_227),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_306),
.A2(n_322),
.B1(n_214),
.B2(n_260),
.Y(n_338)
);

FAx1_ASAP7_75t_SL g312 ( 
.A(n_225),
.B(n_222),
.CI(n_261),
.CON(n_312),
.SN(n_312)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_312),
.B(n_321),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_318),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_219),
.A2(n_222),
.B1(n_266),
.B2(n_244),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_246),
.A2(n_247),
.B1(n_260),
.B2(n_267),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_323),
.A2(n_268),
.B(n_264),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_324),
.B(n_239),
.C(n_253),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_244),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_329),
.B(n_312),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_276),
.A2(n_272),
.B1(n_278),
.B2(n_279),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_328),
.Y(n_333)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_328),
.Y(n_335)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_335),
.Y(n_380)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_330),
.Y(n_337)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_337),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_338),
.A2(n_343),
.B1(n_367),
.B2(n_374),
.Y(n_405)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_330),
.Y(n_339)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_339),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_316),
.B(n_235),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_340),
.B(n_346),
.Y(n_377)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_319),
.Y(n_341)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_341),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_342),
.B(n_369),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_306),
.A2(n_224),
.B1(n_231),
.B2(n_221),
.Y(n_343)
);

OA21x2_ASAP7_75t_L g344 ( 
.A1(n_281),
.A2(n_215),
.B(n_210),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_344),
.A2(n_350),
.B(n_357),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_233),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_345),
.B(n_348),
.C(n_301),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_297),
.B(n_237),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_325),
.A2(n_292),
.B(n_281),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_347),
.A2(n_356),
.B(n_296),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_304),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_354),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_287),
.A2(n_265),
.B1(n_256),
.B2(n_257),
.Y(n_350)
);

A2O1A1Ixp33_ASAP7_75t_L g351 ( 
.A1(n_315),
.A2(n_209),
.B(n_259),
.C(n_211),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_351),
.B(n_368),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_292),
.A2(n_220),
.B1(n_250),
.B2(n_259),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_352),
.A2(n_371),
.B1(n_319),
.B2(n_298),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_305),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_330),
.Y(n_355)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_355),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_323),
.A2(n_228),
.B(n_211),
.Y(n_356)
);

NOR2x1_ASAP7_75t_L g357 ( 
.A(n_315),
.B(n_322),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_305),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_358),
.B(n_360),
.Y(n_384)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_359),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_314),
.B(n_283),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_314),
.B(n_332),
.Y(n_361)
);

NAND3xp33_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_285),
.C(n_310),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_327),
.Y(n_362)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_362),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_363),
.B(n_365),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_305),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_364),
.B(n_370),
.Y(n_399)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_291),
.Y(n_366)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_366),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_329),
.A2(n_324),
.B1(n_289),
.B2(n_312),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_300),
.B(n_326),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_291),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_282),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_308),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_372),
.B(n_373),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_317),
.B(n_307),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_296),
.A2(n_289),
.B1(n_313),
.B2(n_318),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_375),
.A2(n_387),
.B(n_358),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_SL g425 ( 
.A1(n_378),
.A2(n_298),
.B1(n_299),
.B2(n_293),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_365),
.A2(n_307),
.B1(n_301),
.B2(n_290),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_381),
.A2(n_385),
.B1(n_398),
.B2(n_409),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_334),
.A2(n_347),
.B1(n_353),
.B2(n_350),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_354),
.B(n_293),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_373),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_389),
.B(n_370),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_368),
.B(n_285),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_390),
.B(n_396),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_340),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_403),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_334),
.A2(n_290),
.B1(n_303),
.B2(n_294),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_342),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_401),
.B(n_407),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_336),
.B(n_310),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_406),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_336),
.B(n_280),
.Y(n_406)
);

OAI32xp33_ASAP7_75t_L g407 ( 
.A1(n_363),
.A2(n_280),
.A3(n_286),
.B1(n_288),
.B2(n_320),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_334),
.A2(n_303),
.B1(n_294),
.B2(n_302),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_410),
.Y(n_444)
);

AO22x1_ASAP7_75t_L g411 ( 
.A1(n_401),
.A2(n_357),
.B1(n_364),
.B2(n_344),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_411),
.A2(n_412),
.B(n_437),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_375),
.A2(n_379),
.B(n_394),
.Y(n_412)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_415),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_405),
.A2(n_353),
.B1(n_338),
.B2(n_344),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_416),
.A2(n_438),
.B1(n_383),
.B2(n_387),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_395),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_418),
.B(n_424),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_385),
.A2(n_344),
.B1(n_374),
.B2(n_343),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_419),
.A2(n_425),
.B1(n_432),
.B2(n_379),
.Y(n_447)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_376),
.Y(n_421)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_421),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_392),
.B(n_345),
.Y(n_423)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_423),
.Y(n_441)
);

CKINVDCx14_ASAP7_75t_R g424 ( 
.A(n_399),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_388),
.Y(n_426)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_426),
.Y(n_446)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_376),
.Y(n_427)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_427),
.Y(n_452)
);

A2O1A1Ixp33_ASAP7_75t_L g428 ( 
.A1(n_408),
.A2(n_336),
.B(n_357),
.C(n_346),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_428),
.B(n_433),
.Y(n_453)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_380),
.Y(n_429)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_429),
.Y(n_458)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_380),
.Y(n_430)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_430),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_377),
.B(n_335),
.Y(n_431)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_431),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_381),
.A2(n_367),
.B1(n_383),
.B2(n_398),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_377),
.B(n_333),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_395),
.B(n_369),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_434),
.B(n_436),
.Y(n_461)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_402),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_435),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_393),
.B(n_366),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_394),
.A2(n_356),
.B(n_351),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_405),
.A2(n_348),
.B1(n_355),
.B2(n_337),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_390),
.B(n_286),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_439),
.B(n_396),
.C(n_384),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_443),
.B(n_460),
.C(n_412),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_447),
.A2(n_438),
.B1(n_411),
.B2(n_437),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_448),
.A2(n_462),
.B1(n_411),
.B2(n_428),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_404),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_454),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_419),
.A2(n_432),
.B1(n_417),
.B2(n_414),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_450),
.A2(n_455),
.B1(n_465),
.B2(n_429),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_436),
.Y(n_451)
);

CKINVDCx14_ASAP7_75t_R g470 ( 
.A(n_451),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_413),
.B(n_408),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_417),
.A2(n_383),
.B1(n_382),
.B2(n_397),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_422),
.A2(n_391),
.B1(n_382),
.B2(n_397),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_456),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_420),
.B(n_406),
.C(n_387),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_416),
.A2(n_409),
.B1(n_402),
.B2(n_407),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_414),
.A2(n_386),
.B1(n_388),
.B2(n_400),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_420),
.B(n_400),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_439),
.Y(n_474)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_461),
.Y(n_467)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_467),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_462),
.A2(n_448),
.B1(n_464),
.B2(n_453),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_468),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_469),
.B(n_474),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_464),
.A2(n_433),
.B1(n_431),
.B2(n_434),
.Y(n_471)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_471),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_423),
.Y(n_472)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_472),
.Y(n_498)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_440),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_475),
.B(n_484),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_441),
.B(n_427),
.Y(n_476)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_476),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_477),
.A2(n_481),
.B1(n_482),
.B2(n_459),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_478),
.A2(n_483),
.B1(n_458),
.B2(n_459),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_441),
.B(n_457),
.Y(n_479)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_479),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_443),
.B(n_410),
.C(n_435),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_460),
.C(n_466),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_450),
.A2(n_426),
.B1(n_386),
.B2(n_341),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_453),
.A2(n_339),
.B1(n_371),
.B2(n_284),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_452),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_372),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_485),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_465),
.B(n_288),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_487),
.B(n_489),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_454),
.B(n_320),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_488),
.B(n_449),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_455),
.B(n_331),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_444),
.A2(n_311),
.B(n_309),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_490),
.A2(n_458),
.B(n_452),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_495),
.B(n_496),
.Y(n_515)
);

INVx13_ASAP7_75t_L g501 ( 
.A(n_470),
.Y(n_501)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_501),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_468),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_502),
.B(n_504),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_469),
.B(n_444),
.C(n_445),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_505),
.A2(n_445),
.B(n_490),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_507),
.B(n_482),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_471),
.B(n_442),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_487),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_509),
.A2(n_478),
.B1(n_486),
.B2(n_483),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_492),
.B(n_475),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_511),
.B(n_512),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_508),
.B(n_481),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_506),
.C(n_504),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_513),
.B(n_521),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_506),
.B(n_473),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_514),
.B(n_522),
.C(n_524),
.Y(n_525)
);

FAx1_ASAP7_75t_SL g516 ( 
.A(n_498),
.B(n_472),
.CI(n_480),
.CON(n_516),
.SN(n_516)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_516),
.B(n_520),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_518),
.A2(n_497),
.B1(n_489),
.B2(n_499),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_519),
.A2(n_507),
.B(n_503),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_473),
.C(n_474),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_494),
.B(n_477),
.C(n_488),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_523),
.B(n_505),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_479),
.C(n_476),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_510),
.A2(n_492),
.B(n_516),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_527),
.B(n_528),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_529),
.B(n_530),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_518),
.A2(n_493),
.B1(n_500),
.B2(n_503),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_513),
.B(n_493),
.C(n_500),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_532),
.B(n_534),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_524),
.A2(n_493),
.B1(n_491),
.B2(n_498),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_522),
.A2(n_491),
.B1(n_497),
.B2(n_467),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_535),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_536),
.B(n_520),
.Y(n_543)
);

AOI21xp33_ASAP7_75t_L g539 ( 
.A1(n_533),
.A2(n_517),
.B(n_501),
.Y(n_539)
);

AOI31xp33_ASAP7_75t_L g552 ( 
.A1(n_539),
.A2(n_542),
.A3(n_545),
.B(n_485),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_531),
.B(n_515),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_543),
.B(n_535),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_526),
.B(n_515),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_544),
.B(n_525),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_532),
.B(n_521),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_525),
.B(n_514),
.C(n_446),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_546),
.B(n_540),
.Y(n_551)
);

NOR3xp33_ASAP7_75t_L g547 ( 
.A(n_537),
.B(n_529),
.C(n_528),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_547),
.B(n_549),
.Y(n_554)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_548),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_541),
.A2(n_534),
.B1(n_530),
.B2(n_536),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_550),
.B(n_551),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_552),
.A2(n_553),
.B(n_539),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_546),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_555),
.B(n_557),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_547),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_556),
.B(n_558),
.C(n_554),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_560),
.B(n_561),
.C(n_446),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_556),
.B(n_538),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_562),
.B(n_559),
.C(n_463),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_563),
.A2(n_484),
.B(n_499),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_564),
.A2(n_309),
.B(n_308),
.Y(n_565)
);


endmodule