module fake_netlist_1_7013_n_1698 (n_117, n_44, n_361, n_185, n_22, n_57, n_26, n_407, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_383, n_6, n_400, n_296, n_157, n_79, n_202, n_386, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_389, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_387, n_163, n_105, n_227, n_384, n_231, n_298, n_411, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_401, n_28, n_48, n_100, n_305, n_228, n_345, n_360, n_236, n_340, n_150, n_373, n_3, n_18, n_301, n_66, n_222, n_234, n_366, n_286, n_15, n_190, n_246, n_321, n_324, n_392, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_367, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_393, n_24, n_247, n_381, n_304, n_399, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_402, n_32, n_413, n_391, n_235, n_243, n_394, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_404, n_54, n_369, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_362, n_153, n_61, n_259, n_308, n_93, n_412, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_403, n_254, n_262, n_10, n_239, n_87, n_379, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_370, n_34, n_5, n_23, n_8, n_217, n_139, n_388, n_193, n_273, n_390, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_4, n_374, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_365, n_179, n_315, n_363, n_409, n_86, n_143, n_295, n_263, n_166, n_186, n_364, n_75, n_376, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_396, n_168, n_398, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_378, n_359, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_397, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_410, n_63, n_14, n_71, n_56, n_188, n_377, n_343, n_127, n_291, n_170, n_380, n_356, n_281, n_341, n_58, n_122, n_187, n_375, n_138, n_371, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_368, n_355, n_226, n_382, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_372, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_408, n_290, n_405, n_280, n_21, n_99, n_109, n_132, n_395, n_406, n_151, n_385, n_257, n_269, n_1698);
input n_117;
input n_44;
input n_361;
input n_185;
input n_22;
input n_57;
input n_26;
input n_407;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_383;
input n_6;
input n_400;
input n_296;
input n_157;
input n_79;
input n_202;
input n_386;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_389;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_387;
input n_163;
input n_105;
input n_227;
input n_384;
input n_231;
input n_298;
input n_411;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_401;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_360;
input n_236;
input n_340;
input n_150;
input n_373;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_366;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_392;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_367;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_393;
input n_24;
input n_247;
input n_381;
input n_304;
input n_399;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_402;
input n_32;
input n_413;
input n_391;
input n_235;
input n_243;
input n_394;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_404;
input n_54;
input n_369;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_362;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_412;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_403;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_379;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_370;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_388;
input n_193;
input n_273;
input n_390;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_374;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_365;
input n_179;
input n_315;
input n_363;
input n_409;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_364;
input n_75;
input n_376;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_396;
input n_168;
input n_398;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_378;
input n_359;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_397;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_410;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_377;
input n_343;
input n_127;
input n_291;
input n_170;
input n_380;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_375;
input n_138;
input n_371;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_368;
input n_355;
input n_226;
input n_382;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_372;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_408;
input n_290;
input n_405;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_395;
input n_406;
input n_151;
input n_385;
input n_257;
input n_269;
output n_1698;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_1671;
wire n_646;
wire n_1334;
wire n_1627;
wire n_829;
wire n_1603;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1618;
wire n_1477;
wire n_1363;
wire n_1594;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_1646;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_1667;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_1663;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_452;
wire n_518;
wire n_1336;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1672;
wire n_1342;
wire n_1619;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1598;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_1631;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_1661;
wire n_999;
wire n_769;
wire n_624;
wire n_1597;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1683;
wire n_1349;
wire n_1573;
wire n_1580;
wire n_1605;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_1656;
wire n_571;
wire n_1595;
wire n_1604;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_1654;
wire n_551;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_1620;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_1623;
wire n_556;
wire n_1214;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_1438;
wire n_514;
wire n_1693;
wire n_1690;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_1613;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_1582;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_1662;
wire n_790;
wire n_761;
wire n_1660;
wire n_1287;
wire n_472;
wire n_1100;
wire n_1648;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_1695;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1682;
wire n_1213;
wire n_1452;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_1639;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_774;
wire n_1207;
wire n_1463;
wire n_510;
wire n_1075;
wire n_1615;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1590;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1628;
wire n_1533;
wire n_1611;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_1694;
wire n_1563;
wire n_1642;
wire n_824;
wire n_793;
wire n_753;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1600;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_992;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1681;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1602;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_1557;
wire n_911;
wire n_980;
wire n_1675;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_1606;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1625;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_1629;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1670;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_1581;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_1643;
wire n_1687;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_550;
wire n_826;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1608;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_478;
wire n_482;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1427;
wire n_1050;
wire n_1593;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_1647;
wire n_1621;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1668;
wire n_1692;
wire n_1153;
wire n_1657;
wire n_1655;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_733;
wire n_894;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_1665;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1696;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_1638;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1645;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_1633;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1626;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_688;
wire n_515;
wire n_1577;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1641;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_1583;
wire n_606;
wire n_1585;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_1586;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_1697;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_1599;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1679;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_1688;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_1634;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_1455;
wire n_659;
wire n_432;
wire n_1329;
wire n_1572;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_436;
wire n_1653;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1640;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_1579;
wire n_609;
wire n_909;
wire n_1273;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1658;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_1575;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_1659;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_1635;
wire n_871;
wire n_803;
wire n_1429;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_516;
wire n_549;
wire n_1576;
wire n_1609;
wire n_832;
wire n_996;
wire n_1578;
wire n_420;
wire n_1684;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1610;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_1678;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1674;
wire n_1351;
wire n_1318;
wire n_956;
wire n_1622;
wire n_1614;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_495;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1612;
wire n_1636;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1587;
wire n_1489;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1689;
wire n_1592;
wire n_1168;
wire n_1574;
wire n_458;
wire n_1084;
wire n_1624;
wire n_618;
wire n_1596;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_1616;
wire n_1378;
wire n_1570;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_757;
wire n_1568;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_1676;
wire n_678;
wire n_1200;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_481;
wire n_443;
wire n_694;
wire n_1601;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_1666;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1680;
wire n_1644;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1518;
wire n_945;
wire n_1669;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1673;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_1589;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_1630;
wire n_784;
wire n_1491;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1637;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1617;
wire n_1632;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_1664;
wire n_682;
wire n_1607;
wire n_906;
wire n_1650;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1591;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_1685;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1335;
wire n_1239;
wire n_924;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1677;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1649;
wire n_1143;
wire n_629;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_1691;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_1686;
wire n_600;
wire n_1531;
wire n_1548;
wire n_1651;
wire n_1584;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_1588;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_1652;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_1398;
wire n_491;
wire n_1291;
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_227), .Y(n_414) );
INVx4_ASAP7_75t_R g415 ( .A(n_37), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_366), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_410), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_393), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_10), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_17), .Y(n_420) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_294), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_50), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_29), .Y(n_423) );
CKINVDCx14_ASAP7_75t_R g424 ( .A(n_265), .Y(n_424) );
INVxp67_ASAP7_75t_SL g425 ( .A(n_408), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_217), .Y(n_426) );
INVx2_ASAP7_75t_SL g427 ( .A(n_214), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_158), .B(n_166), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_18), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_4), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_259), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_162), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_40), .Y(n_433) );
INVxp67_ASAP7_75t_SL g434 ( .A(n_361), .Y(n_434) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_43), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_35), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_35), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_92), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_306), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_45), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_189), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_151), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_187), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_360), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_107), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_236), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_177), .Y(n_447) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_305), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_132), .Y(n_449) );
INVxp67_ASAP7_75t_L g450 ( .A(n_19), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_271), .Y(n_451) );
CKINVDCx16_ASAP7_75t_R g452 ( .A(n_375), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_183), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_71), .Y(n_454) );
CKINVDCx16_ASAP7_75t_R g455 ( .A(n_44), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_209), .Y(n_456) );
CKINVDCx16_ASAP7_75t_R g457 ( .A(n_330), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_32), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_291), .Y(n_459) );
INVxp67_ASAP7_75t_SL g460 ( .A(n_200), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_221), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_147), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_91), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_274), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_204), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_145), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_94), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_402), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_353), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_395), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_287), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_129), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_280), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_186), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_278), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_254), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_67), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_301), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_237), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_332), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_12), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_356), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_290), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_93), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_295), .Y(n_485) );
INVxp67_ASAP7_75t_L g486 ( .A(n_336), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_197), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_136), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_285), .Y(n_489) );
INVx2_ASAP7_75t_SL g490 ( .A(n_303), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_81), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_173), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_47), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_26), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_0), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_193), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_78), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_131), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_2), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_30), .Y(n_500) );
INVx2_ASAP7_75t_SL g501 ( .A(n_138), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_401), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_143), .Y(n_503) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_213), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_399), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_230), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_59), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_235), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_53), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_203), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_86), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_144), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_329), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_110), .Y(n_514) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_226), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g516 ( .A(n_211), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_222), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_325), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_277), .Y(n_519) );
INVxp33_ASAP7_75t_L g520 ( .A(n_334), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_157), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_122), .Y(n_522) );
BUFx3_ASAP7_75t_L g523 ( .A(n_299), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_153), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_148), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_154), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_205), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_11), .Y(n_528) );
BUFx5_ASAP7_75t_L g529 ( .A(n_263), .Y(n_529) );
CKINVDCx16_ASAP7_75t_R g530 ( .A(n_286), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_267), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_215), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_121), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_270), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_99), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_381), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_249), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_78), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_312), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_201), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_3), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_93), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_170), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_155), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_98), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_169), .Y(n_546) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_252), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_99), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_146), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_92), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_164), .Y(n_551) );
BUFx3_ASAP7_75t_L g552 ( .A(n_335), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_279), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_324), .Y(n_554) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_239), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_218), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_390), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_405), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_135), .Y(n_559) );
BUFx3_ASAP7_75t_L g560 ( .A(n_308), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_319), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_128), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_117), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_413), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_191), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_380), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_242), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_185), .Y(n_568) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_89), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_384), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_135), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_316), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_296), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_192), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_409), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_8), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_269), .B(n_387), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_37), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_33), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_46), .Y(n_580) );
NOR2xp67_ASAP7_75t_L g581 ( .A(n_121), .B(n_292), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_179), .Y(n_582) );
XNOR2xp5_ASAP7_75t_L g583 ( .A(n_302), .B(n_36), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_127), .Y(n_584) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_273), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_317), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_262), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_412), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_98), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_394), .Y(n_590) );
BUFx3_ASAP7_75t_L g591 ( .A(n_379), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_161), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_261), .Y(n_593) );
CKINVDCx16_ASAP7_75t_R g594 ( .A(n_310), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_10), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_300), .Y(n_596) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_234), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_126), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_398), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_293), .Y(n_600) );
CKINVDCx16_ASAP7_75t_R g601 ( .A(n_43), .Y(n_601) );
BUFx10_ASAP7_75t_L g602 ( .A(n_272), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_133), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_314), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_365), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_309), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_66), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_69), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_59), .Y(n_609) );
INVxp33_ASAP7_75t_SL g610 ( .A(n_11), .Y(n_610) );
BUFx2_ASAP7_75t_L g611 ( .A(n_102), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_255), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_529), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_421), .Y(n_614) );
AND2x4_ASAP7_75t_L g615 ( .A(n_421), .B(n_0), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_454), .B(n_1), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_529), .Y(n_617) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_448), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_452), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_468), .B(n_1), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_468), .Y(n_621) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_448), .Y(n_622) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_448), .Y(n_623) );
XOR2xp5_ASAP7_75t_L g624 ( .A(n_437), .B(n_2), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_445), .B(n_3), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_487), .Y(n_626) );
AND2x4_ASAP7_75t_L g627 ( .A(n_487), .B(n_5), .Y(n_627) );
OA21x2_ASAP7_75t_L g628 ( .A1(n_447), .A2(n_140), .B(n_139), .Y(n_628) );
INVxp67_ASAP7_75t_L g629 ( .A(n_445), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_430), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_430), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_529), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_484), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_484), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_529), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_529), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_611), .B(n_6), .Y(n_637) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_450), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_455), .A2(n_8), .B1(n_6), .B2(n_7), .Y(n_639) );
INVx3_ASAP7_75t_L g640 ( .A(n_602), .Y(n_640) );
NOR2x1_ASAP7_75t_L g641 ( .A(n_581), .B(n_7), .Y(n_641) );
INVx4_ASAP7_75t_L g642 ( .A(n_523), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_497), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_529), .Y(n_644) );
OA21x2_ASAP7_75t_L g645 ( .A1(n_447), .A2(n_142), .B(n_141), .Y(n_645) );
AND2x4_ASAP7_75t_L g646 ( .A(n_497), .B(n_9), .Y(n_646) );
INVx4_ASAP7_75t_L g647 ( .A(n_523), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_559), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_501), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_427), .B(n_9), .Y(n_650) );
INVx3_ASAP7_75t_L g651 ( .A(n_602), .Y(n_651) );
AND2x2_ASAP7_75t_SL g652 ( .A(n_577), .B(n_149), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_559), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_457), .Y(n_654) );
BUFx2_ASAP7_75t_L g655 ( .A(n_629), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_615), .A2(n_423), .B1(n_429), .B2(n_419), .Y(n_656) );
INVx1_ASAP7_75t_SL g657 ( .A(n_619), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_613), .Y(n_658) );
NAND2xp33_ASAP7_75t_L g659 ( .A(n_614), .B(n_414), .Y(n_659) );
INVx4_ASAP7_75t_L g660 ( .A(n_615), .Y(n_660) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_625), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_640), .B(n_520), .Y(n_662) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_618), .Y(n_663) );
INVx2_ASAP7_75t_SL g664 ( .A(n_640), .Y(n_664) );
NAND2xp33_ASAP7_75t_L g665 ( .A(n_614), .B(n_418), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_618), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_621), .B(n_601), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_618), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_613), .Y(n_669) );
BUFx3_ASAP7_75t_L g670 ( .A(n_628), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_621), .B(n_626), .Y(n_671) );
INVx5_ASAP7_75t_L g672 ( .A(n_642), .Y(n_672) );
AND2x6_ASAP7_75t_L g673 ( .A(n_615), .B(n_552), .Y(n_673) );
OR2x2_ASAP7_75t_L g674 ( .A(n_626), .B(n_638), .Y(n_674) );
INVx1_ASAP7_75t_SL g675 ( .A(n_654), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_640), .B(n_530), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_640), .B(n_520), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_642), .B(n_490), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_642), .B(n_453), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_642), .B(n_453), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_613), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_618), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_617), .Y(n_683) );
INVx3_ASAP7_75t_L g684 ( .A(n_646), .Y(n_684) );
BUFx8_ASAP7_75t_SL g685 ( .A(n_651), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_618), .Y(n_686) );
INVx3_ASAP7_75t_L g687 ( .A(n_646), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_618), .Y(n_688) );
INVx5_ASAP7_75t_L g689 ( .A(n_647), .Y(n_689) );
BUFx3_ASAP7_75t_L g690 ( .A(n_628), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_622), .Y(n_691) );
INVx4_ASAP7_75t_L g692 ( .A(n_615), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_617), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_664), .Y(n_694) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_655), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_684), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_684), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_664), .Y(n_698) );
INVx3_ASAP7_75t_L g699 ( .A(n_660), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_660), .B(n_652), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_662), .B(n_651), .Y(n_701) );
CKINVDCx5p33_ASAP7_75t_R g702 ( .A(n_655), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_660), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_660), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_661), .B(n_625), .Y(n_705) );
NOR3xp33_ASAP7_75t_L g706 ( .A(n_667), .B(n_639), .C(n_637), .Y(n_706) );
INVx2_ASAP7_75t_SL g707 ( .A(n_674), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_671), .B(n_651), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_692), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_684), .A2(n_652), .B1(n_646), .B2(n_627), .Y(n_710) );
NOR2xp67_ASAP7_75t_L g711 ( .A(n_667), .B(n_651), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_671), .B(n_620), .Y(n_712) );
AND2x4_ASAP7_75t_SL g713 ( .A(n_692), .B(n_466), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_677), .B(n_620), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_692), .B(n_620), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_692), .B(n_652), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_687), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_673), .B(n_620), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_673), .B(n_656), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_687), .Y(n_720) );
A2O1A1Ixp33_ASAP7_75t_SL g721 ( .A1(n_687), .A2(n_650), .B(n_617), .C(n_635), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_687), .A2(n_646), .B1(n_627), .B2(n_635), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_673), .A2(n_627), .B1(n_635), .B2(n_632), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_679), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_673), .B(n_627), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_676), .B(n_649), .Y(n_726) );
BUFx5_ASAP7_75t_L g727 ( .A(n_673), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_673), .A2(n_632), .B1(n_636), .B2(n_644), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_659), .B(n_616), .Y(n_729) );
INVx2_ASAP7_75t_SL g730 ( .A(n_674), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_665), .B(n_647), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_673), .B(n_647), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_678), .B(n_547), .Y(n_733) );
AND2x6_ASAP7_75t_L g734 ( .A(n_670), .B(n_552), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_658), .A2(n_632), .B1(n_636), .B2(n_644), .Y(n_735) );
INVxp67_ASAP7_75t_L g736 ( .A(n_657), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_658), .A2(n_636), .B1(n_610), .B2(n_631), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_678), .B(n_594), .Y(n_738) );
AND2x2_ASAP7_75t_SL g739 ( .A(n_679), .B(n_628), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_669), .B(n_424), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_669), .B(n_424), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_681), .B(n_653), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_680), .Y(n_743) );
NOR2xp67_ASAP7_75t_L g744 ( .A(n_680), .B(n_583), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_681), .B(n_630), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_675), .B(n_420), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_683), .A2(n_610), .B1(n_631), .B2(n_630), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_683), .B(n_633), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_693), .Y(n_749) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_675), .A2(n_624), .B1(n_493), .B2(n_437), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_672), .B(n_634), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_672), .B(n_634), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_672), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_672), .B(n_653), .Y(n_754) );
OR2x2_ASAP7_75t_L g755 ( .A(n_685), .B(n_624), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_672), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_670), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_672), .B(n_648), .Y(n_758) );
INVx5_ASAP7_75t_L g759 ( .A(n_672), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_670), .A2(n_648), .B1(n_643), .B2(n_438), .Y(n_760) );
A2O1A1Ixp33_ASAP7_75t_L g761 ( .A1(n_690), .A2(n_643), .B(n_440), .C(n_463), .Y(n_761) );
INVx1_ASAP7_75t_SL g762 ( .A(n_689), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_689), .B(n_439), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_690), .A2(n_472), .B1(n_477), .B2(n_433), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_689), .B(n_442), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_689), .B(n_456), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_690), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_689), .A2(n_471), .B1(n_475), .B2(n_466), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_666), .A2(n_481), .B1(n_494), .B2(n_488), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_703), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_705), .B(n_422), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_715), .A2(n_645), .B(n_628), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g773 ( .A1(n_739), .A2(n_645), .B(n_428), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_708), .B(n_436), .Y(n_774) );
INVxp67_ASAP7_75t_L g775 ( .A(n_695), .Y(n_775) );
INVx3_ASAP7_75t_L g776 ( .A(n_699), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g777 ( .A1(n_739), .A2(n_645), .B(n_434), .Y(n_777) );
NAND2xp5_ASAP7_75t_SL g778 ( .A(n_736), .B(n_503), .Y(n_778) );
BUFx12f_ASAP7_75t_L g779 ( .A(n_702), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_708), .B(n_449), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_712), .B(n_458), .Y(n_781) );
NAND2xp5_ASAP7_75t_SL g782 ( .A(n_727), .B(n_503), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_710), .A2(n_532), .B1(n_539), .B2(n_518), .Y(n_783) );
AOI21xp5_ASAP7_75t_L g784 ( .A1(n_714), .A2(n_645), .B(n_460), .Y(n_784) );
A2O1A1Ixp33_ASAP7_75t_L g785 ( .A1(n_712), .A2(n_500), .B(n_507), .C(n_498), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g786 ( .A1(n_718), .A2(n_515), .B(n_425), .Y(n_786) );
NAND2xp5_ASAP7_75t_SL g787 ( .A(n_727), .B(n_518), .Y(n_787) );
AOI21xp5_ASAP7_75t_L g788 ( .A1(n_725), .A2(n_417), .B(n_416), .Y(n_788) );
INVx3_ASAP7_75t_L g789 ( .A(n_699), .Y(n_789) );
NAND2xp5_ASAP7_75t_SL g790 ( .A(n_727), .B(n_532), .Y(n_790) );
O2A1O1Ixp5_ASAP7_75t_L g791 ( .A1(n_716), .A2(n_496), .B(n_508), .C(n_464), .Y(n_791) );
AOI22x1_ASAP7_75t_L g792 ( .A1(n_757), .A2(n_623), .B1(n_622), .B2(n_508), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_716), .A2(n_574), .B1(n_582), .B2(n_539), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_707), .B(n_467), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_696), .Y(n_795) );
AO21x1_ASAP7_75t_L g796 ( .A1(n_767), .A2(n_431), .B(n_426), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_732), .A2(n_441), .B(n_432), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_730), .B(n_491), .Y(n_798) );
AOI21xp5_ASAP7_75t_L g799 ( .A1(n_721), .A2(n_444), .B(n_443), .Y(n_799) );
INVx5_ASAP7_75t_L g800 ( .A(n_734), .Y(n_800) );
BUFx6f_ASAP7_75t_L g801 ( .A(n_759), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_711), .B(n_495), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_704), .Y(n_803) );
AOI21xp5_ASAP7_75t_L g804 ( .A1(n_721), .A2(n_451), .B(n_446), .Y(n_804) );
BUFx2_ASAP7_75t_L g805 ( .A(n_768), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_724), .B(n_499), .Y(n_806) );
NAND2xp5_ASAP7_75t_SL g807 ( .A(n_727), .B(n_723), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_726), .B(n_574), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_701), .A2(n_741), .B(n_740), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_743), .B(n_511), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_750), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_710), .A2(n_722), .B1(n_713), .B2(n_764), .Y(n_812) );
BUFx12f_ASAP7_75t_L g813 ( .A(n_755), .Y(n_813) );
OAI21xp33_ASAP7_75t_L g814 ( .A1(n_733), .A2(n_533), .B(n_528), .Y(n_814) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_746), .Y(n_815) );
AND2x2_ASAP7_75t_L g816 ( .A(n_744), .B(n_550), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_738), .B(n_538), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_737), .B(n_571), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_747), .B(n_580), .Y(n_819) );
A2O1A1Ixp33_ASAP7_75t_L g820 ( .A1(n_729), .A2(n_514), .B(n_522), .C(n_509), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_747), .B(n_584), .Y(n_821) );
BUFx3_ASAP7_75t_L g822 ( .A(n_751), .Y(n_822) );
INVx5_ASAP7_75t_L g823 ( .A(n_734), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_729), .B(n_598), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g825 ( .A1(n_697), .A2(n_465), .B(n_461), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_726), .B(n_582), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_717), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_706), .B(n_608), .Y(n_828) );
AOI21x1_ASAP7_75t_L g829 ( .A1(n_719), .A2(n_668), .B(n_666), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_720), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_764), .B(n_535), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_709), .B(n_727), .Y(n_832) );
BUFx12f_ASAP7_75t_L g833 ( .A(n_734), .Y(n_833) );
BUFx12f_ASAP7_75t_L g834 ( .A(n_734), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_742), .Y(n_835) );
INVxp67_ASAP7_75t_L g836 ( .A(n_745), .Y(n_836) );
BUFx2_ASAP7_75t_L g837 ( .A(n_734), .Y(n_837) );
OAI21xp5_ASAP7_75t_L g838 ( .A1(n_760), .A2(n_641), .B(n_476), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_731), .A2(n_478), .B(n_473), .Y(n_839) );
AO21x2_ASAP7_75t_L g840 ( .A1(n_748), .A2(n_483), .B(n_480), .Y(n_840) );
AO21x1_ASAP7_75t_L g841 ( .A1(n_731), .A2(n_492), .B(n_485), .Y(n_841) );
AO22x1_ASAP7_75t_L g842 ( .A1(n_749), .A2(n_641), .B1(n_459), .B2(n_470), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_727), .B(n_541), .Y(n_843) );
A2O1A1Ixp33_ASAP7_75t_L g844 ( .A1(n_722), .A2(n_545), .B(n_548), .C(n_542), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_694), .Y(n_845) );
AND2x4_ASAP7_75t_L g846 ( .A(n_723), .B(n_562), .Y(n_846) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_698), .B(n_563), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_728), .B(n_576), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_728), .A2(n_595), .B1(n_603), .B2(n_579), .Y(n_849) );
AOI21xp5_ASAP7_75t_L g850 ( .A1(n_763), .A2(n_505), .B(n_502), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_762), .B(n_607), .Y(n_851) );
AO21x1_ASAP7_75t_L g852 ( .A1(n_752), .A2(n_510), .B(n_506), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g853 ( .A1(n_765), .A2(n_517), .B(n_513), .Y(n_853) );
AOI21xp5_ASAP7_75t_L g854 ( .A1(n_766), .A2(n_521), .B(n_519), .Y(n_854) );
BUFx6f_ASAP7_75t_L g855 ( .A(n_759), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_769), .B(n_609), .Y(n_856) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_753), .B(n_469), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g858 ( .A(n_756), .B(n_486), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_735), .A2(n_589), .B1(n_578), .B2(n_525), .Y(n_859) );
BUFx2_ASAP7_75t_L g860 ( .A(n_754), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_735), .B(n_589), .Y(n_861) );
NAND2xp5_ASAP7_75t_SL g862 ( .A(n_759), .B(n_758), .Y(n_862) );
AOI221xp5_ASAP7_75t_L g863 ( .A1(n_759), .A2(n_569), .B1(n_435), .B2(n_587), .C(n_526), .Y(n_863) );
INVx1_ASAP7_75t_SL g864 ( .A(n_713), .Y(n_864) );
BUFx2_ASAP7_75t_L g865 ( .A(n_702), .Y(n_865) );
AOI33xp33_ASAP7_75t_L g866 ( .A1(n_707), .A2(n_534), .A3(n_527), .B1(n_536), .B2(n_531), .B3(n_524), .Y(n_866) );
AOI21xp5_ASAP7_75t_L g867 ( .A1(n_715), .A2(n_546), .B(n_540), .Y(n_867) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_707), .B(n_462), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_705), .B(n_474), .Y(n_869) );
NAND2xp5_ASAP7_75t_SL g870 ( .A(n_736), .B(n_479), .Y(n_870) );
NAND2xp5_ASAP7_75t_SL g871 ( .A(n_736), .B(n_482), .Y(n_871) );
A2O1A1Ixp33_ASAP7_75t_L g872 ( .A1(n_712), .A2(n_553), .B(n_554), .C(n_551), .Y(n_872) );
NAND2xp5_ASAP7_75t_SL g873 ( .A(n_736), .B(n_489), .Y(n_873) );
INVx2_ASAP7_75t_SL g874 ( .A(n_713), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_700), .A2(n_558), .B1(n_561), .B2(n_556), .Y(n_875) );
NOR2xp33_ASAP7_75t_R g876 ( .A(n_702), .B(n_516), .Y(n_876) );
OAI21xp5_ASAP7_75t_L g877 ( .A1(n_739), .A2(n_565), .B(n_564), .Y(n_877) );
O2A1O1Ixp33_ASAP7_75t_L g878 ( .A1(n_761), .A2(n_567), .B(n_568), .C(n_566), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_705), .B(n_537), .Y(n_879) );
INVx5_ASAP7_75t_L g880 ( .A(n_734), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_705), .B(n_543), .Y(n_881) );
AO21x1_ASAP7_75t_L g882 ( .A1(n_700), .A2(n_575), .B(n_572), .Y(n_882) );
NAND2xp5_ASAP7_75t_SL g883 ( .A(n_736), .B(n_544), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_707), .B(n_435), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_705), .B(n_570), .Y(n_885) );
INVx2_ASAP7_75t_L g886 ( .A(n_703), .Y(n_886) );
INVx4_ASAP7_75t_L g887 ( .A(n_713), .Y(n_887) );
AOI21xp5_ASAP7_75t_L g888 ( .A1(n_772), .A2(n_588), .B(n_586), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_836), .B(n_435), .Y(n_889) );
OAI22x1_ASAP7_75t_L g890 ( .A1(n_805), .A2(n_590), .B1(n_593), .B2(n_592), .Y(n_890) );
NAND2xp5_ASAP7_75t_SL g891 ( .A(n_864), .B(n_573), .Y(n_891) );
OAI21xp5_ASAP7_75t_L g892 ( .A1(n_777), .A2(n_600), .B(n_596), .Y(n_892) );
AOI21xp5_ASAP7_75t_L g893 ( .A1(n_773), .A2(n_606), .B(n_605), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_770), .Y(n_894) );
AO31x2_ASAP7_75t_L g895 ( .A1(n_852), .A2(n_464), .A3(n_549), .B(n_512), .Y(n_895) );
AO32x2_ASAP7_75t_L g896 ( .A1(n_859), .A2(n_623), .A3(n_622), .B1(n_569), .B2(n_435), .Y(n_896) );
AOI21xp5_ASAP7_75t_L g897 ( .A1(n_809), .A2(n_612), .B(n_668), .Y(n_897) );
INVx4_ASAP7_75t_L g898 ( .A(n_779), .Y(n_898) );
INVx4_ASAP7_75t_L g899 ( .A(n_887), .Y(n_899) );
OAI21xp5_ASAP7_75t_L g900 ( .A1(n_784), .A2(n_549), .B(n_512), .Y(n_900) );
OAI21x1_ASAP7_75t_L g901 ( .A1(n_829), .A2(n_792), .B(n_799), .Y(n_901) );
INVx3_ASAP7_75t_L g902 ( .A(n_887), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_835), .B(n_569), .Y(n_903) );
INVxp67_ASAP7_75t_SL g904 ( .A(n_783), .Y(n_904) );
AOI21xp5_ASAP7_75t_L g905 ( .A1(n_807), .A2(n_691), .B(n_682), .Y(n_905) );
AOI21x1_ASAP7_75t_L g906 ( .A1(n_804), .A2(n_682), .B(n_668), .Y(n_906) );
OA21x2_ASAP7_75t_L g907 ( .A1(n_877), .A2(n_599), .B(n_557), .Y(n_907) );
OAI21x1_ASAP7_75t_L g908 ( .A1(n_791), .A2(n_599), .B(n_557), .Y(n_908) );
INVxp67_ASAP7_75t_SL g909 ( .A(n_812), .Y(n_909) );
AOI21xp5_ASAP7_75t_L g910 ( .A1(n_806), .A2(n_686), .B(n_682), .Y(n_910) );
NOR2xp33_ASAP7_75t_L g911 ( .A(n_808), .B(n_585), .Y(n_911) );
OAI21x1_ASAP7_75t_L g912 ( .A1(n_877), .A2(n_688), .B(n_686), .Y(n_912) );
AOI221x1_ASAP7_75t_L g913 ( .A1(n_838), .A2(n_623), .B1(n_622), .B2(n_504), .C(n_555), .Y(n_913) );
A2O1A1Ixp33_ASAP7_75t_L g914 ( .A1(n_878), .A2(n_591), .B(n_560), .C(n_569), .Y(n_914) );
AND2x4_ASAP7_75t_L g915 ( .A(n_874), .B(n_560), .Y(n_915) );
AOI21xp5_ASAP7_75t_L g916 ( .A1(n_810), .A2(n_688), .B(n_686), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_828), .B(n_597), .Y(n_917) );
AO21x2_ASAP7_75t_L g918 ( .A1(n_882), .A2(n_691), .B(n_688), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_884), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_846), .B(n_604), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_846), .B(n_12), .Y(n_921) );
BUFx6f_ASAP7_75t_L g922 ( .A(n_801), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_851), .Y(n_923) );
A2O1A1Ixp33_ASAP7_75t_L g924 ( .A1(n_843), .A2(n_448), .B(n_555), .C(n_504), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_793), .A2(n_504), .B1(n_555), .B2(n_415), .Y(n_925) );
BUFx12f_ASAP7_75t_L g926 ( .A(n_813), .Y(n_926) );
AO31x2_ASAP7_75t_L g927 ( .A1(n_841), .A2(n_623), .A3(n_622), .B(n_555), .Y(n_927) );
INVx2_ASAP7_75t_L g928 ( .A(n_803), .Y(n_928) );
NOR2xp33_ASAP7_75t_L g929 ( .A(n_826), .B(n_775), .Y(n_929) );
AOI21xp5_ASAP7_75t_L g930 ( .A1(n_797), .A2(n_663), .B(n_623), .Y(n_930) );
CKINVDCx20_ASAP7_75t_R g931 ( .A(n_865), .Y(n_931) );
AOI21xp5_ASAP7_75t_L g932 ( .A1(n_839), .A2(n_663), .B(n_623), .Y(n_932) );
NAND3xp33_ASAP7_75t_SL g933 ( .A(n_876), .B(n_811), .C(n_864), .Y(n_933) );
A2O1A1Ixp33_ASAP7_75t_L g934 ( .A1(n_867), .A2(n_663), .B(n_15), .C(n_13), .Y(n_934) );
AO21x2_ASAP7_75t_L g935 ( .A1(n_796), .A2(n_840), .B(n_838), .Y(n_935) );
BUFx6f_ASAP7_75t_L g936 ( .A(n_801), .Y(n_936) );
INVx5_ASAP7_75t_L g937 ( .A(n_801), .Y(n_937) );
AOI21xp5_ASAP7_75t_L g938 ( .A1(n_832), .A2(n_663), .B(n_152), .Y(n_938) );
CKINVDCx6p67_ASAP7_75t_R g939 ( .A(n_778), .Y(n_939) );
NOR2x1_ASAP7_75t_SL g940 ( .A(n_833), .B(n_13), .Y(n_940) );
OR2x6_ASAP7_75t_L g941 ( .A(n_834), .B(n_815), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_849), .A2(n_16), .B1(n_14), .B2(n_15), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_845), .Y(n_943) );
AOI21xp5_ASAP7_75t_L g944 ( .A1(n_788), .A2(n_156), .B(n_150), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_785), .B(n_14), .Y(n_945) );
AO31x2_ASAP7_75t_L g946 ( .A1(n_859), .A2(n_21), .A3(n_19), .B(n_20), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_844), .B(n_20), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_795), .Y(n_948) );
AOI21xp5_ASAP7_75t_L g949 ( .A1(n_850), .A2(n_160), .B(n_159), .Y(n_949) );
AOI21xp5_ASAP7_75t_L g950 ( .A1(n_853), .A2(n_165), .B(n_163), .Y(n_950) );
AOI21xp5_ASAP7_75t_L g951 ( .A1(n_854), .A2(n_817), .B(n_824), .Y(n_951) );
AO21x2_ASAP7_75t_L g952 ( .A1(n_840), .A2(n_168), .B(n_167), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_827), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_830), .Y(n_954) );
AOI221xp5_ASAP7_75t_L g955 ( .A1(n_771), .A2(n_24), .B1(n_22), .B2(n_23), .C(n_25), .Y(n_955) );
AOI21x1_ASAP7_75t_L g956 ( .A1(n_861), .A2(n_172), .B(n_171), .Y(n_956) );
AOI21xp5_ASAP7_75t_L g957 ( .A1(n_781), .A2(n_175), .B(n_174), .Y(n_957) );
OAI21x1_ASAP7_75t_L g958 ( .A1(n_862), .A2(n_178), .B(n_176), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_820), .B(n_24), .Y(n_959) );
AO31x2_ASAP7_75t_L g960 ( .A1(n_872), .A2(n_28), .A3(n_26), .B(n_27), .Y(n_960) );
AOI21xp5_ASAP7_75t_L g961 ( .A1(n_774), .A2(n_181), .B(n_180), .Y(n_961) );
NAND2x1p5_ASAP7_75t_L g962 ( .A(n_855), .B(n_28), .Y(n_962) );
OA21x2_ASAP7_75t_L g963 ( .A1(n_825), .A2(n_184), .B(n_182), .Y(n_963) );
CKINVDCx20_ASAP7_75t_R g964 ( .A(n_794), .Y(n_964) );
INVx5_ASAP7_75t_L g965 ( .A(n_855), .Y(n_965) );
BUFx6f_ASAP7_75t_L g966 ( .A(n_855), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_831), .A2(n_34), .B1(n_31), .B2(n_32), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_866), .B(n_34), .Y(n_968) );
INVx2_ASAP7_75t_L g969 ( .A(n_886), .Y(n_969) );
NOR2xp67_ASAP7_75t_L g970 ( .A(n_798), .B(n_36), .Y(n_970) );
BUFx6f_ASAP7_75t_L g971 ( .A(n_822), .Y(n_971) );
BUFx6f_ASAP7_75t_L g972 ( .A(n_860), .Y(n_972) );
HB1xp67_ASAP7_75t_L g973 ( .A(n_782), .Y(n_973) );
NAND2xp5_ASAP7_75t_SL g974 ( .A(n_868), .B(n_38), .Y(n_974) );
AND2x4_ASAP7_75t_L g975 ( .A(n_800), .B(n_38), .Y(n_975) );
AO31x2_ASAP7_75t_L g976 ( .A1(n_837), .A2(n_41), .A3(n_39), .B(n_40), .Y(n_976) );
A2O1A1Ixp33_ASAP7_75t_L g977 ( .A1(n_875), .A2(n_42), .B(n_39), .C(n_41), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_800), .A2(n_45), .B1(n_42), .B2(n_44), .Y(n_978) );
OR2x2_ASAP7_75t_L g979 ( .A(n_869), .B(n_46), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_819), .B(n_47), .Y(n_980) );
AO31x2_ASAP7_75t_L g981 ( .A1(n_848), .A2(n_50), .A3(n_48), .B(n_49), .Y(n_981) );
INVx2_ASAP7_75t_L g982 ( .A(n_776), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_776), .Y(n_983) );
AO31x2_ASAP7_75t_L g984 ( .A1(n_847), .A2(n_51), .A3(n_48), .B(n_49), .Y(n_984) );
OAI21xp5_ASAP7_75t_L g985 ( .A1(n_786), .A2(n_190), .B(n_188), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_821), .B(n_51), .Y(n_986) );
AO31x2_ASAP7_75t_L g987 ( .A1(n_856), .A2(n_55), .A3(n_52), .B(n_54), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_789), .Y(n_988) );
OAI21xp5_ASAP7_75t_L g989 ( .A1(n_780), .A2(n_195), .B(n_194), .Y(n_989) );
OAI21x1_ASAP7_75t_L g990 ( .A1(n_789), .A2(n_198), .B(n_196), .Y(n_990) );
AO31x2_ASAP7_75t_L g991 ( .A1(n_857), .A2(n_57), .A3(n_55), .B(n_56), .Y(n_991) );
CKINVDCx16_ASAP7_75t_R g992 ( .A(n_816), .Y(n_992) );
OR2x2_ASAP7_75t_L g993 ( .A(n_879), .B(n_56), .Y(n_993) );
BUFx2_ASAP7_75t_L g994 ( .A(n_800), .Y(n_994) );
INVx3_ASAP7_75t_SL g995 ( .A(n_870), .Y(n_995) );
NOR2xp33_ASAP7_75t_L g996 ( .A(n_814), .B(n_57), .Y(n_996) );
AO31x2_ASAP7_75t_L g997 ( .A1(n_858), .A2(n_61), .A3(n_58), .B(n_60), .Y(n_997) );
CKINVDCx11_ASAP7_75t_R g998 ( .A(n_842), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_881), .B(n_58), .Y(n_999) );
CKINVDCx5p33_ASAP7_75t_R g1000 ( .A(n_871), .Y(n_1000) );
CKINVDCx11_ASAP7_75t_R g1001 ( .A(n_873), .Y(n_1001) );
AO31x2_ASAP7_75t_L g1002 ( .A1(n_802), .A2(n_62), .A3(n_60), .B(n_61), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_885), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_818), .Y(n_1004) );
NAND2x1p5_ASAP7_75t_L g1005 ( .A(n_800), .B(n_62), .Y(n_1005) );
NAND2xp5_ASAP7_75t_SL g1006 ( .A(n_823), .B(n_63), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_823), .A2(n_880), .B1(n_790), .B2(n_787), .Y(n_1007) );
AO32x2_ASAP7_75t_L g1008 ( .A1(n_863), .A2(n_63), .A3(n_64), .B1(n_65), .B2(n_66), .Y(n_1008) );
NOR2xp33_ASAP7_75t_L g1009 ( .A(n_883), .B(n_65), .Y(n_1009) );
NAND2x1p5_ASAP7_75t_L g1010 ( .A(n_823), .B(n_67), .Y(n_1010) );
AOI21xp5_ASAP7_75t_L g1011 ( .A1(n_823), .A2(n_202), .B(n_199), .Y(n_1011) );
BUFx10_ASAP7_75t_L g1012 ( .A(n_880), .Y(n_1012) );
INVx2_ASAP7_75t_L g1013 ( .A(n_880), .Y(n_1013) );
AOI21xp5_ASAP7_75t_L g1014 ( .A1(n_880), .A2(n_207), .B(n_206), .Y(n_1014) );
CKINVDCx11_ASAP7_75t_R g1015 ( .A(n_779), .Y(n_1015) );
AOI21xp5_ASAP7_75t_L g1016 ( .A1(n_772), .A2(n_210), .B(n_208), .Y(n_1016) );
A2O1A1Ixp33_ASAP7_75t_L g1017 ( .A1(n_809), .A2(n_68), .B(n_69), .C(n_70), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_836), .Y(n_1018) );
OAI21x1_ASAP7_75t_L g1019 ( .A1(n_829), .A2(n_216), .B(n_212), .Y(n_1019) );
CKINVDCx6p67_ASAP7_75t_R g1020 ( .A(n_779), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_836), .Y(n_1021) );
OAI21x1_ASAP7_75t_L g1022 ( .A1(n_829), .A2(n_220), .B(n_219), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_836), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_836), .B(n_72), .Y(n_1024) );
A2O1A1Ixp33_ASAP7_75t_L g1025 ( .A1(n_809), .A2(n_73), .B(n_74), .C(n_75), .Y(n_1025) );
AOI21xp5_ASAP7_75t_L g1026 ( .A1(n_772), .A2(n_224), .B(n_223), .Y(n_1026) );
OA21x2_ASAP7_75t_L g1027 ( .A1(n_773), .A2(n_228), .B(n_225), .Y(n_1027) );
BUFx3_ASAP7_75t_L g1028 ( .A(n_779), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_836), .B(n_74), .Y(n_1029) );
OR2x2_ASAP7_75t_L g1030 ( .A(n_783), .B(n_75), .Y(n_1030) );
AO21x1_ASAP7_75t_L g1031 ( .A1(n_777), .A2(n_231), .B(n_229), .Y(n_1031) );
BUFx12f_ASAP7_75t_L g1032 ( .A(n_779), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_836), .Y(n_1033) );
AND2x4_ASAP7_75t_L g1034 ( .A(n_887), .B(n_76), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_836), .B(n_76), .Y(n_1035) );
CKINVDCx20_ASAP7_75t_R g1036 ( .A(n_865), .Y(n_1036) );
OAI21x1_ASAP7_75t_L g1037 ( .A1(n_829), .A2(n_233), .B(n_232), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_836), .Y(n_1038) );
INVx2_ASAP7_75t_L g1039 ( .A(n_948), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1018), .Y(n_1040) );
BUFx2_ASAP7_75t_L g1041 ( .A(n_931), .Y(n_1041) );
CKINVDCx20_ASAP7_75t_R g1042 ( .A(n_1015), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1021), .Y(n_1043) );
OAI21xp5_ASAP7_75t_L g1044 ( .A1(n_893), .A2(n_77), .B(n_79), .Y(n_1044) );
AOI21x1_ASAP7_75t_L g1045 ( .A1(n_913), .A2(n_240), .B(n_238), .Y(n_1045) );
OAI21x1_ASAP7_75t_L g1046 ( .A1(n_901), .A2(n_906), .B(n_912), .Y(n_1046) );
INVx4_ASAP7_75t_L g1047 ( .A(n_937), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1023), .Y(n_1048) );
AOI21x1_ASAP7_75t_L g1049 ( .A1(n_913), .A2(n_243), .B(n_241), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_909), .B(n_77), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_923), .B(n_79), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1033), .Y(n_1052) );
AOI21xp5_ASAP7_75t_L g1053 ( .A1(n_951), .A2(n_245), .B(n_244), .Y(n_1053) );
OAI21x1_ASAP7_75t_L g1054 ( .A1(n_906), .A2(n_247), .B(n_246), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_904), .B(n_80), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1038), .Y(n_1056) );
AND2x4_ASAP7_75t_L g1057 ( .A(n_937), .B(n_81), .Y(n_1057) );
OA21x2_ASAP7_75t_L g1058 ( .A1(n_900), .A2(n_250), .B(n_248), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_1003), .B(n_82), .Y(n_1059) );
NAND2x1p5_ASAP7_75t_L g1060 ( .A(n_899), .B(n_82), .Y(n_1060) );
AOI21x1_ASAP7_75t_L g1061 ( .A1(n_956), .A2(n_253), .B(n_251), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_929), .A2(n_83), .B1(n_84), .B2(n_85), .Y(n_1062) );
OAI21x1_ASAP7_75t_L g1063 ( .A1(n_1019), .A2(n_257), .B(n_256), .Y(n_1063) );
INVx2_ASAP7_75t_L g1064 ( .A(n_953), .Y(n_1064) );
BUFx12f_ASAP7_75t_L g1065 ( .A(n_1032), .Y(n_1065) );
OAI21x1_ASAP7_75t_L g1066 ( .A1(n_1022), .A2(n_260), .B(n_258), .Y(n_1066) );
AOI21x1_ASAP7_75t_L g1067 ( .A1(n_956), .A2(n_266), .B(n_264), .Y(n_1067) );
INVx2_ASAP7_75t_L g1068 ( .A(n_954), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_1004), .B(n_84), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1029), .B(n_85), .Y(n_1070) );
AOI21xp33_ASAP7_75t_SL g1071 ( .A1(n_1030), .A2(n_941), .B(n_1034), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_943), .Y(n_1072) );
OR2x2_ASAP7_75t_L g1073 ( .A(n_992), .B(n_86), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1074 ( .A(n_1035), .B(n_87), .Y(n_1074) );
AND2x4_ASAP7_75t_L g1075 ( .A(n_937), .B(n_87), .Y(n_1075) );
AOI221xp5_ASAP7_75t_SL g1076 ( .A1(n_1017), .A2(n_88), .B1(n_89), .B2(n_90), .C(n_91), .Y(n_1076) );
INVx2_ASAP7_75t_L g1077 ( .A(n_894), .Y(n_1077) );
AO31x2_ASAP7_75t_L g1078 ( .A1(n_1031), .A2(n_90), .A3(n_94), .B(n_95), .Y(n_1078) );
AO21x2_ASAP7_75t_L g1079 ( .A1(n_892), .A2(n_275), .B(n_268), .Y(n_1079) );
INVx2_ASAP7_75t_SL g1080 ( .A(n_972), .Y(n_1080) );
INVx3_ASAP7_75t_L g1081 ( .A(n_965), .Y(n_1081) );
INVx2_ASAP7_75t_L g1082 ( .A(n_928), .Y(n_1082) );
AOI21xp5_ASAP7_75t_L g1083 ( .A1(n_888), .A2(n_281), .B(n_276), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_968), .Y(n_1084) );
AO31x2_ASAP7_75t_L g1085 ( .A1(n_924), .A2(n_95), .A3(n_96), .B(n_97), .Y(n_1085) );
OAI21xp5_ASAP7_75t_L g1086 ( .A1(n_897), .A2(n_96), .B(n_97), .Y(n_1086) );
BUFx2_ASAP7_75t_L g1087 ( .A(n_1036), .Y(n_1087) );
AOI22xp33_ASAP7_75t_SL g1088 ( .A1(n_1034), .A2(n_100), .B1(n_101), .B2(n_102), .Y(n_1088) );
AO21x2_ASAP7_75t_L g1089 ( .A1(n_935), .A2(n_326), .B(n_407), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_903), .Y(n_1090) );
AOI21xp5_ASAP7_75t_L g1091 ( .A1(n_930), .A2(n_323), .B(n_406), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_999), .B(n_101), .Y(n_1092) );
BUFx2_ASAP7_75t_L g1093 ( .A(n_971), .Y(n_1093) );
OA21x2_ASAP7_75t_L g1094 ( .A1(n_1037), .A2(n_327), .B(n_404), .Y(n_1094) );
OA21x2_ASAP7_75t_L g1095 ( .A1(n_908), .A2(n_322), .B(n_403), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_964), .A2(n_103), .B1(n_104), .B2(n_105), .Y(n_1096) );
OAI21x1_ASAP7_75t_L g1097 ( .A1(n_905), .A2(n_321), .B(n_400), .Y(n_1097) );
AO21x2_ASAP7_75t_L g1098 ( .A1(n_989), .A2(n_320), .B(n_397), .Y(n_1098) );
AO31x2_ASAP7_75t_L g1099 ( .A1(n_1016), .A2(n_103), .A3(n_104), .B(n_105), .Y(n_1099) );
INVx1_ASAP7_75t_L g1100 ( .A(n_889), .Y(n_1100) );
HB1xp67_ASAP7_75t_L g1101 ( .A(n_971), .Y(n_1101) );
AOI21xp5_ASAP7_75t_L g1102 ( .A1(n_932), .A2(n_328), .B(n_396), .Y(n_1102) );
AOI22xp5_ASAP7_75t_L g1103 ( .A1(n_942), .A2(n_106), .B1(n_107), .B2(n_108), .Y(n_1103) );
AOI21xp5_ASAP7_75t_L g1104 ( .A1(n_1026), .A2(n_331), .B(n_392), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_960), .Y(n_1105) );
AND2x4_ASAP7_75t_L g1106 ( .A(n_965), .B(n_106), .Y(n_1106) );
AOI21xp5_ASAP7_75t_L g1107 ( .A1(n_910), .A2(n_318), .B(n_391), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_960), .Y(n_1108) );
BUFx3_ASAP7_75t_L g1109 ( .A(n_926), .Y(n_1109) );
NAND2x1p5_ASAP7_75t_L g1110 ( .A(n_965), .B(n_108), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1024), .Y(n_1111) );
INVx2_ASAP7_75t_L g1112 ( .A(n_969), .Y(n_1112) );
INVx3_ASAP7_75t_L g1113 ( .A(n_922), .Y(n_1113) );
OAI21x1_ASAP7_75t_L g1114 ( .A1(n_990), .A2(n_333), .B(n_389), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_946), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_946), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_959), .Y(n_1117) );
AO21x2_ASAP7_75t_L g1118 ( .A1(n_918), .A2(n_315), .B(n_388), .Y(n_1118) );
HB1xp67_ASAP7_75t_L g1119 ( .A(n_975), .Y(n_1119) );
OAI22xp5_ASAP7_75t_L g1120 ( .A1(n_921), .A2(n_109), .B1(n_110), .B2(n_111), .Y(n_1120) );
OR2x2_ASAP7_75t_L g1121 ( .A(n_939), .B(n_111), .Y(n_1121) );
AO22x2_ASAP7_75t_L g1122 ( .A1(n_975), .A2(n_112), .B1(n_113), .B2(n_114), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_987), .Y(n_1123) );
AOI21xp33_ASAP7_75t_SL g1124 ( .A1(n_995), .A2(n_112), .B(n_113), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_979), .B(n_115), .Y(n_1125) );
INVx1_ASAP7_75t_L g1126 ( .A(n_987), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_993), .Y(n_1127) );
AO21x1_ASAP7_75t_L g1128 ( .A1(n_1005), .A2(n_116), .B(n_118), .Y(n_1128) );
BUFx2_ASAP7_75t_L g1129 ( .A(n_1020), .Y(n_1129) );
INVx3_ASAP7_75t_L g1130 ( .A(n_922), .Y(n_1130) );
OA21x2_ASAP7_75t_L g1131 ( .A1(n_985), .A2(n_338), .B(n_386), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_984), .Y(n_1132) );
AO31x2_ASAP7_75t_L g1133 ( .A1(n_1025), .A2(n_116), .A3(n_119), .B(n_120), .Y(n_1133) );
OAI21xp5_ASAP7_75t_L g1134 ( .A1(n_914), .A2(n_119), .B(n_120), .Y(n_1134) );
INVx2_ASAP7_75t_L g1135 ( .A(n_927), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_984), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_981), .Y(n_1137) );
NOR2x1_ASAP7_75t_SL g1138 ( .A(n_936), .B(n_122), .Y(n_1138) );
NOR2xp33_ASAP7_75t_L g1139 ( .A(n_933), .B(n_123), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_973), .A2(n_123), .B1(n_124), .B2(n_125), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_890), .B(n_124), .Y(n_1141) );
BUFx8_ASAP7_75t_L g1142 ( .A(n_1028), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_920), .B(n_125), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_991), .Y(n_1144) );
AOI21xp5_ASAP7_75t_L g1145 ( .A1(n_916), .A2(n_341), .B(n_385), .Y(n_1145) );
NOR2xp33_ASAP7_75t_L g1146 ( .A(n_917), .B(n_126), .Y(n_1146) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_915), .B(n_127), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_998), .B(n_128), .Y(n_1148) );
CKINVDCx5p33_ASAP7_75t_R g1149 ( .A(n_898), .Y(n_1149) );
CKINVDCx20_ASAP7_75t_R g1150 ( .A(n_1001), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_911), .B(n_129), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_991), .Y(n_1152) );
AND2x4_ASAP7_75t_L g1153 ( .A(n_902), .B(n_130), .Y(n_1153) );
AND2x4_ASAP7_75t_L g1154 ( .A(n_936), .B(n_130), .Y(n_1154) );
NAND2x1_ASAP7_75t_L g1155 ( .A(n_966), .B(n_282), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_925), .A2(n_131), .B1(n_132), .B2(n_133), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_997), .Y(n_1157) );
NOR2xp67_ASAP7_75t_L g1158 ( .A(n_966), .B(n_346), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_919), .B(n_134), .Y(n_1159) );
AO21x2_ASAP7_75t_L g1160 ( .A1(n_952), .A2(n_345), .B(n_383), .Y(n_1160) );
OAI21x1_ASAP7_75t_L g1161 ( .A1(n_958), .A2(n_344), .B(n_382), .Y(n_1161) );
INVx11_ASAP7_75t_L g1162 ( .A(n_940), .Y(n_1162) );
OAI21x1_ASAP7_75t_L g1163 ( .A1(n_938), .A2(n_343), .B(n_378), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_980), .B(n_134), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_945), .B(n_136), .Y(n_1165) );
OR2x6_ASAP7_75t_L g1166 ( .A(n_1010), .B(n_137), .Y(n_1166) );
AOI21x1_ASAP7_75t_L g1167 ( .A1(n_907), .A2(n_347), .B(n_377), .Y(n_1167) );
CKINVDCx5p33_ASAP7_75t_R g1168 ( .A(n_1000), .Y(n_1168) );
AO21x2_ASAP7_75t_L g1169 ( .A1(n_934), .A2(n_342), .B(n_376), .Y(n_1169) );
OAI21xp5_ASAP7_75t_L g1170 ( .A1(n_947), .A2(n_137), .B(n_138), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_915), .B(n_283), .Y(n_1171) );
AO21x2_ASAP7_75t_L g1172 ( .A1(n_1006), .A2(n_284), .B(n_288), .Y(n_1172) );
INVx2_ASAP7_75t_L g1173 ( .A(n_927), .Y(n_1173) );
NAND2xp5_ASAP7_75t_L g1174 ( .A(n_970), .B(n_289), .Y(n_1174) );
INVx1_ASAP7_75t_SL g1175 ( .A(n_962), .Y(n_1175) );
INVx2_ASAP7_75t_L g1176 ( .A(n_927), .Y(n_1176) );
OAI21x1_ASAP7_75t_L g1177 ( .A1(n_1027), .A2(n_297), .B(n_298), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_986), .B(n_411), .Y(n_1178) );
INVxp67_ASAP7_75t_L g1179 ( .A(n_1009), .Y(n_1179) );
BUFx3_ASAP7_75t_L g1180 ( .A(n_1012), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_982), .B(n_304), .Y(n_1181) );
AOI21xp33_ASAP7_75t_L g1182 ( .A1(n_1007), .A2(n_307), .B(n_311), .Y(n_1182) );
OR2x2_ASAP7_75t_L g1183 ( .A(n_891), .B(n_313), .Y(n_1183) );
BUFx3_ASAP7_75t_L g1184 ( .A(n_994), .Y(n_1184) );
AOI21xp5_ASAP7_75t_L g1185 ( .A1(n_957), .A2(n_337), .B(n_339), .Y(n_1185) );
NOR2xp33_ASAP7_75t_L g1186 ( .A(n_974), .B(n_340), .Y(n_1186) );
INVx4_ASAP7_75t_L g1187 ( .A(n_994), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_997), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_955), .B(n_374), .Y(n_1189) );
NOR2x1p5_ASAP7_75t_L g1190 ( .A(n_1013), .B(n_348), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_996), .B(n_988), .Y(n_1191) );
A2O1A1Ixp33_ASAP7_75t_L g1192 ( .A1(n_977), .A2(n_349), .B(n_350), .C(n_351), .Y(n_1192) );
BUFx2_ASAP7_75t_L g1193 ( .A(n_983), .Y(n_1193) );
NOR2xp67_ASAP7_75t_L g1194 ( .A(n_961), .B(n_352), .Y(n_1194) );
HB1xp67_ASAP7_75t_L g1195 ( .A(n_967), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1002), .Y(n_1196) );
OA21x2_ASAP7_75t_L g1197 ( .A1(n_944), .A2(n_354), .B(n_355), .Y(n_1197) );
INVx8_ASAP7_75t_L g1198 ( .A(n_1065), .Y(n_1198) );
BUFx3_ASAP7_75t_L g1199 ( .A(n_1081), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1040), .Y(n_1200) );
INVx2_ASAP7_75t_L g1201 ( .A(n_1135), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1043), .Y(n_1202) );
OR2x6_ASAP7_75t_L g1203 ( .A(n_1166), .B(n_978), .Y(n_1203) );
OR2x6_ASAP7_75t_L g1204 ( .A(n_1166), .B(n_1011), .Y(n_1204) );
AO21x2_ASAP7_75t_L g1205 ( .A1(n_1196), .A2(n_949), .B(n_950), .Y(n_1205) );
INVx2_ASAP7_75t_L g1206 ( .A(n_1173), .Y(n_1206) );
INVx2_ASAP7_75t_L g1207 ( .A(n_1176), .Y(n_1207) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1084), .B(n_895), .Y(n_1208) );
INVx2_ASAP7_75t_SL g1209 ( .A(n_1142), .Y(n_1209) );
OR2x6_ASAP7_75t_L g1210 ( .A(n_1166), .B(n_1014), .Y(n_1210) );
OR2x2_ASAP7_75t_L g1211 ( .A(n_1147), .B(n_1002), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1048), .Y(n_1212) );
AOI221xp5_ASAP7_75t_L g1213 ( .A1(n_1071), .A2(n_1008), .B1(n_976), .B2(n_896), .C(n_963), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1052), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1117), .B(n_896), .Y(n_1215) );
AND2x4_ASAP7_75t_L g1216 ( .A(n_1081), .B(n_357), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1056), .Y(n_1217) );
INVx2_ASAP7_75t_L g1218 ( .A(n_1039), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1064), .Y(n_1219) );
INVx2_ASAP7_75t_L g1220 ( .A(n_1068), .Y(n_1220) );
INVx2_ASAP7_75t_L g1221 ( .A(n_1072), .Y(n_1221) );
INVx3_ASAP7_75t_L g1222 ( .A(n_1047), .Y(n_1222) );
OR2x6_ASAP7_75t_L g1223 ( .A(n_1110), .B(n_358), .Y(n_1223) );
NOR2xp33_ASAP7_75t_L g1224 ( .A(n_1071), .B(n_359), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1051), .Y(n_1225) );
INVxp67_ASAP7_75t_SL g1226 ( .A(n_1119), .Y(n_1226) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1077), .Y(n_1227) );
AO21x2_ASAP7_75t_L g1228 ( .A1(n_1123), .A2(n_1137), .B(n_1126), .Y(n_1228) );
INVx3_ASAP7_75t_L g1229 ( .A(n_1047), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1051), .Y(n_1230) );
INVx2_ASAP7_75t_L g1231 ( .A(n_1082), .Y(n_1231) );
OR2x2_ASAP7_75t_L g1232 ( .A(n_1041), .B(n_362), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1122), .B(n_363), .Y(n_1233) );
INVx2_ASAP7_75t_L g1234 ( .A(n_1112), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1159), .Y(n_1235) );
OR2x6_ASAP7_75t_L g1236 ( .A(n_1057), .B(n_364), .Y(n_1236) );
NOR2xp33_ASAP7_75t_L g1237 ( .A(n_1179), .B(n_367), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1195), .B(n_368), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1111), .B(n_369), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1159), .Y(n_1240) );
BUFx2_ASAP7_75t_L g1241 ( .A(n_1180), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1122), .Y(n_1242) );
OR2x2_ASAP7_75t_L g1243 ( .A(n_1087), .B(n_370), .Y(n_1243) );
A2O1A1Ixp33_ASAP7_75t_L g1244 ( .A1(n_1044), .A2(n_373), .B(n_371), .C(n_372), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1153), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1059), .Y(n_1246) );
OAI21x1_ASAP7_75t_L g1247 ( .A1(n_1177), .A2(n_1067), .B(n_1061), .Y(n_1247) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1141), .Y(n_1248) );
INVx2_ASAP7_75t_L g1249 ( .A(n_1054), .Y(n_1249) );
HB1xp67_ASAP7_75t_L g1250 ( .A(n_1187), .Y(n_1250) );
BUFx2_ASAP7_75t_L g1251 ( .A(n_1093), .Y(n_1251) );
HB1xp67_ASAP7_75t_L g1252 ( .A(n_1187), .Y(n_1252) );
HB1xp67_ASAP7_75t_L g1253 ( .A(n_1184), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1075), .Y(n_1254) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1106), .Y(n_1255) );
AO21x2_ASAP7_75t_L g1256 ( .A1(n_1132), .A2(n_1136), .B(n_1188), .Y(n_1256) );
OAI21xp5_ASAP7_75t_L g1257 ( .A1(n_1055), .A2(n_1050), .B(n_1044), .Y(n_1257) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1080), .B(n_1073), .Y(n_1258) );
OA21x2_ASAP7_75t_L g1259 ( .A1(n_1115), .A2(n_1116), .B(n_1108), .Y(n_1259) );
OR2x6_ASAP7_75t_L g1260 ( .A(n_1106), .B(n_1060), .Y(n_1260) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1127), .Y(n_1261) );
INVx4_ASAP7_75t_L g1262 ( .A(n_1109), .Y(n_1262) );
AND2x4_ASAP7_75t_SL g1263 ( .A(n_1101), .B(n_1154), .Y(n_1263) );
AO21x2_ASAP7_75t_L g1264 ( .A1(n_1144), .A2(n_1152), .B(n_1157), .Y(n_1264) );
AND2x4_ASAP7_75t_L g1265 ( .A(n_1113), .B(n_1130), .Y(n_1265) );
INVx2_ASAP7_75t_L g1266 ( .A(n_1167), .Y(n_1266) );
AO21x2_ASAP7_75t_L g1267 ( .A1(n_1105), .A2(n_1045), .B(n_1049), .Y(n_1267) );
OR2x6_ASAP7_75t_L g1268 ( .A(n_1129), .B(n_1190), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1148), .B(n_1096), .Y(n_1269) );
INVx3_ASAP7_75t_L g1270 ( .A(n_1162), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1069), .Y(n_1271) );
BUFx2_ASAP7_75t_L g1272 ( .A(n_1142), .Y(n_1272) );
OA21x2_ASAP7_75t_L g1273 ( .A1(n_1076), .A2(n_1063), .B(n_1066), .Y(n_1273) );
BUFx3_ASAP7_75t_L g1274 ( .A(n_1113), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1193), .B(n_1088), .Y(n_1275) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1050), .Y(n_1276) );
HB1xp67_ASAP7_75t_L g1277 ( .A(n_1154), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1055), .Y(n_1278) );
OR2x6_ASAP7_75t_L g1279 ( .A(n_1171), .B(n_1086), .Y(n_1279) );
HB1xp67_ASAP7_75t_L g1280 ( .A(n_1175), .Y(n_1280) );
BUFx3_ASAP7_75t_L g1281 ( .A(n_1130), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1092), .B(n_1139), .Y(n_1282) );
OR2x2_ASAP7_75t_L g1283 ( .A(n_1092), .B(n_1125), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1120), .Y(n_1284) );
HB1xp67_ASAP7_75t_L g1285 ( .A(n_1175), .Y(n_1285) );
BUFx12f_ASAP7_75t_L g1286 ( .A(n_1149), .Y(n_1286) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1120), .Y(n_1287) );
AO21x2_ASAP7_75t_L g1288 ( .A1(n_1118), .A2(n_1134), .B(n_1089), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1121), .B(n_1146), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1168), .B(n_1070), .Y(n_1290) );
OAI21x1_ASAP7_75t_L g1291 ( .A1(n_1114), .A2(n_1161), .B(n_1097), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1103), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1103), .Y(n_1293) );
NOR2xp33_ASAP7_75t_L g1294 ( .A(n_1074), .B(n_1143), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1124), .B(n_1062), .Y(n_1295) );
INVx3_ASAP7_75t_L g1296 ( .A(n_1183), .Y(n_1296) );
AO21x2_ASAP7_75t_L g1297 ( .A1(n_1118), .A2(n_1134), .B(n_1089), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1128), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1170), .B(n_1140), .Y(n_1299) );
NOR2xp33_ASAP7_75t_L g1300 ( .A(n_1151), .B(n_1165), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1164), .B(n_1191), .Y(n_1301) );
AOI21xp5_ASAP7_75t_SL g1302 ( .A1(n_1138), .A2(n_1131), .B(n_1192), .Y(n_1302) );
OAI21x1_ASAP7_75t_L g1303 ( .A1(n_1053), .A2(n_1163), .B(n_1095), .Y(n_1303) );
NAND2x1_ASAP7_75t_L g1304 ( .A(n_1158), .B(n_1058), .Y(n_1304) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1164), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1133), .B(n_1076), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1133), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1133), .Y(n_1308) );
INVx4_ASAP7_75t_SL g1309 ( .A(n_1085), .Y(n_1309) );
AO21x2_ASAP7_75t_L g1310 ( .A1(n_1160), .A2(n_1098), .B(n_1182), .Y(n_1310) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1099), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1099), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1085), .B(n_1150), .Y(n_1313) );
AO21x2_ASAP7_75t_L g1314 ( .A1(n_1160), .A2(n_1098), .B(n_1182), .Y(n_1314) );
HB1xp67_ASAP7_75t_L g1315 ( .A(n_1090), .Y(n_1315) );
INVxp67_ASAP7_75t_L g1316 ( .A(n_1181), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1078), .Y(n_1317) );
OR2x2_ASAP7_75t_L g1318 ( .A(n_1078), .B(n_1156), .Y(n_1318) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1078), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1181), .Y(n_1320) );
INVx2_ASAP7_75t_L g1321 ( .A(n_1094), .Y(n_1321) );
INVx5_ASAP7_75t_SL g1322 ( .A(n_1042), .Y(n_1322) );
AO21x2_ASAP7_75t_L g1323 ( .A1(n_1194), .A2(n_1169), .B(n_1079), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1186), .B(n_1189), .Y(n_1324) );
BUFx12f_ASAP7_75t_L g1325 ( .A(n_1158), .Y(n_1325) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1100), .Y(n_1326) );
AO21x2_ASAP7_75t_L g1327 ( .A1(n_1169), .A2(n_1079), .B(n_1178), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1174), .Y(n_1328) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1172), .Y(n_1329) );
OA21x2_ASAP7_75t_L g1330 ( .A1(n_1091), .A2(n_1104), .B(n_1102), .Y(n_1330) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1155), .Y(n_1331) );
INVx3_ASAP7_75t_L g1332 ( .A(n_1197), .Y(n_1332) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1083), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1107), .B(n_1145), .Y(n_1334) );
AO21x2_ASAP7_75t_L g1335 ( .A1(n_1185), .A2(n_1196), .B(n_1046), .Y(n_1335) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1200), .Y(n_1336) );
OR2x2_ASAP7_75t_L g1337 ( .A(n_1253), .B(n_1315), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1220), .B(n_1221), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1220), .B(n_1221), .Y(n_1339) );
NAND2xp5_ASAP7_75t_L g1340 ( .A(n_1261), .B(n_1282), .Y(n_1340) );
INVx2_ASAP7_75t_L g1341 ( .A(n_1201), .Y(n_1341) );
INVx2_ASAP7_75t_L g1342 ( .A(n_1201), .Y(n_1342) );
INVx2_ASAP7_75t_SL g1343 ( .A(n_1250), .Y(n_1343) );
INVx3_ASAP7_75t_L g1344 ( .A(n_1206), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1276), .B(n_1278), .Y(n_1345) );
INVx2_ASAP7_75t_L g1346 ( .A(n_1207), .Y(n_1346) );
INVx2_ASAP7_75t_L g1347 ( .A(n_1207), .Y(n_1347) );
INVx4_ASAP7_75t_L g1348 ( .A(n_1236), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1227), .B(n_1231), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1202), .B(n_1212), .Y(n_1350) );
INVx2_ASAP7_75t_L g1351 ( .A(n_1259), .Y(n_1351) );
INVxp67_ASAP7_75t_SL g1352 ( .A(n_1252), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1231), .B(n_1234), .Y(n_1353) );
BUFx2_ASAP7_75t_L g1354 ( .A(n_1252), .Y(n_1354) );
HB1xp67_ASAP7_75t_L g1355 ( .A(n_1315), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_1234), .B(n_1307), .Y(n_1356) );
HB1xp67_ASAP7_75t_L g1357 ( .A(n_1280), .Y(n_1357) );
HB1xp67_ASAP7_75t_L g1358 ( .A(n_1280), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1214), .Y(n_1359) );
OR2x2_ASAP7_75t_L g1360 ( .A(n_1219), .B(n_1218), .Y(n_1360) );
OR2x6_ASAP7_75t_L g1361 ( .A(n_1236), .B(n_1203), .Y(n_1361) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1217), .Y(n_1362) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1308), .B(n_1311), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1312), .B(n_1306), .Y(n_1364) );
AND2x4_ASAP7_75t_L g1365 ( .A(n_1309), .B(n_1256), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1317), .B(n_1319), .Y(n_1366) );
INVx1_ASAP7_75t_SL g1367 ( .A(n_1241), .Y(n_1367) );
NAND2x1_ASAP7_75t_L g1368 ( .A(n_1268), .B(n_1236), .Y(n_1368) );
OR2x2_ASAP7_75t_L g1369 ( .A(n_1285), .B(n_1242), .Y(n_1369) );
HB1xp67_ASAP7_75t_L g1370 ( .A(n_1285), .Y(n_1370) );
OR2x2_ASAP7_75t_L g1371 ( .A(n_1226), .B(n_1248), .Y(n_1371) );
OR2x2_ASAP7_75t_L g1372 ( .A(n_1226), .B(n_1251), .Y(n_1372) );
BUFx3_ASAP7_75t_L g1373 ( .A(n_1199), .Y(n_1373) );
OR2x2_ASAP7_75t_L g1374 ( .A(n_1258), .B(n_1313), .Y(n_1374) );
NAND3xp33_ASAP7_75t_L g1375 ( .A(n_1298), .B(n_1300), .C(n_1294), .Y(n_1375) );
INVx2_ASAP7_75t_SL g1376 ( .A(n_1199), .Y(n_1376) );
NAND2xp5_ASAP7_75t_L g1377 ( .A(n_1292), .B(n_1293), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1256), .B(n_1264), .Y(n_1378) );
INVx3_ASAP7_75t_L g1379 ( .A(n_1268), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_1264), .B(n_1326), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_1257), .B(n_1228), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1257), .B(n_1228), .Y(n_1382) );
HB1xp67_ASAP7_75t_L g1383 ( .A(n_1277), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1208), .B(n_1305), .Y(n_1384) );
BUFx6f_ASAP7_75t_L g1385 ( .A(n_1204), .Y(n_1385) );
NAND2x1p5_ASAP7_75t_L g1386 ( .A(n_1270), .B(n_1262), .Y(n_1386) );
INVx2_ASAP7_75t_SL g1387 ( .A(n_1222), .Y(n_1387) );
HB1xp67_ASAP7_75t_L g1388 ( .A(n_1277), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1389 ( .A(n_1208), .B(n_1225), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1289), .B(n_1290), .Y(n_1390) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1245), .Y(n_1391) );
AND2x2_ASAP7_75t_L g1392 ( .A(n_1230), .B(n_1309), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1309), .B(n_1235), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_1240), .B(n_1275), .Y(n_1394) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1301), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1284), .B(n_1287), .Y(n_1396) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1215), .B(n_1316), .Y(n_1397) );
AND2x4_ASAP7_75t_SL g1398 ( .A(n_1270), .B(n_1260), .Y(n_1398) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_1203), .A2(n_1299), .B1(n_1295), .B2(n_1300), .Y(n_1399) );
NOR2xp33_ASAP7_75t_L g1400 ( .A(n_1269), .B(n_1283), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1215), .B(n_1316), .Y(n_1401) );
INVx1_ASAP7_75t_SL g1402 ( .A(n_1272), .Y(n_1402) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1254), .Y(n_1403) );
OR2x2_ASAP7_75t_L g1404 ( .A(n_1211), .B(n_1279), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1279), .B(n_1318), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1246), .B(n_1271), .Y(n_1406) );
INVx2_ASAP7_75t_L g1407 ( .A(n_1321), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1279), .B(n_1320), .Y(n_1408) );
INVx2_ASAP7_75t_SL g1409 ( .A(n_1222), .Y(n_1409) );
OR2x2_ASAP7_75t_L g1410 ( .A(n_1232), .B(n_1243), .Y(n_1410) );
NAND2xp5_ASAP7_75t_L g1411 ( .A(n_1294), .B(n_1203), .Y(n_1411) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1255), .Y(n_1412) );
NAND2xp5_ASAP7_75t_L g1413 ( .A(n_1296), .B(n_1263), .Y(n_1413) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1229), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1415 ( .A(n_1233), .B(n_1296), .Y(n_1415) );
NOR2x1_ASAP7_75t_L g1416 ( .A(n_1260), .B(n_1223), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1213), .B(n_1288), .Y(n_1417) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1213), .B(n_1288), .Y(n_1418) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1216), .Y(n_1419) );
AND2x2_ASAP7_75t_L g1420 ( .A(n_1297), .B(n_1328), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1421 ( .A(n_1297), .B(n_1335), .Y(n_1421) );
INVx3_ASAP7_75t_L g1422 ( .A(n_1304), .Y(n_1422) );
AND2x4_ASAP7_75t_SL g1423 ( .A(n_1260), .B(n_1223), .Y(n_1423) );
INVx2_ASAP7_75t_SL g1424 ( .A(n_1263), .Y(n_1424) );
AND2x2_ASAP7_75t_L g1425 ( .A(n_1335), .B(n_1329), .Y(n_1425) );
NAND2xp5_ASAP7_75t_L g1426 ( .A(n_1324), .B(n_1265), .Y(n_1426) );
NOR2xp33_ASAP7_75t_L g1427 ( .A(n_1237), .B(n_1239), .Y(n_1427) );
AOI22xp33_ASAP7_75t_L g1428 ( .A1(n_1204), .A2(n_1210), .B1(n_1223), .B2(n_1224), .Y(n_1428) );
NOR2xp33_ASAP7_75t_L g1429 ( .A(n_1237), .B(n_1239), .Y(n_1429) );
INVx1_ASAP7_75t_SL g1430 ( .A(n_1209), .Y(n_1430) );
HB1xp67_ASAP7_75t_L g1431 ( .A(n_1274), .Y(n_1431) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1238), .Y(n_1432) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1238), .Y(n_1433) );
AND2x4_ASAP7_75t_L g1434 ( .A(n_1204), .B(n_1210), .Y(n_1434) );
NAND2xp5_ASAP7_75t_L g1435 ( .A(n_1265), .B(n_1224), .Y(n_1435) );
NAND2xp5_ASAP7_75t_L g1436 ( .A(n_1281), .B(n_1210), .Y(n_1436) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1325), .Y(n_1437) );
INVx2_ASAP7_75t_L g1438 ( .A(n_1351), .Y(n_1438) );
NAND2xp5_ASAP7_75t_L g1439 ( .A(n_1395), .B(n_1322), .Y(n_1439) );
AND3x1_ASAP7_75t_L g1440 ( .A(n_1416), .B(n_1198), .C(n_1322), .Y(n_1440) );
AND2x4_ASAP7_75t_L g1441 ( .A(n_1434), .B(n_1331), .Y(n_1441) );
INVx2_ASAP7_75t_L g1442 ( .A(n_1351), .Y(n_1442) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1336), .Y(n_1443) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1359), .Y(n_1444) );
NAND2xp5_ASAP7_75t_L g1445 ( .A(n_1400), .B(n_1333), .Y(n_1445) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1362), .Y(n_1446) );
AND2x4_ASAP7_75t_L g1447 ( .A(n_1434), .B(n_1332), .Y(n_1447) );
INVx2_ASAP7_75t_SL g1448 ( .A(n_1343), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1449 ( .A(n_1364), .B(n_1332), .Y(n_1449) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1350), .Y(n_1450) );
OR2x2_ASAP7_75t_L g1451 ( .A(n_1355), .B(n_1267), .Y(n_1451) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1363), .Y(n_1452) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1363), .Y(n_1453) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1366), .Y(n_1454) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1364), .B(n_1267), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_1400), .B(n_1244), .Y(n_1456) );
AOI22xp33_ASAP7_75t_L g1457 ( .A1(n_1361), .A2(n_1334), .B1(n_1205), .B2(n_1327), .Y(n_1457) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1366), .Y(n_1458) );
INVx2_ASAP7_75t_L g1459 ( .A(n_1407), .Y(n_1459) );
NAND2xp5_ASAP7_75t_SL g1460 ( .A(n_1348), .B(n_1244), .Y(n_1460) );
NAND2xp5_ASAP7_75t_L g1461 ( .A(n_1340), .B(n_1273), .Y(n_1461) );
AND2x4_ASAP7_75t_SL g1462 ( .A(n_1348), .B(n_1198), .Y(n_1462) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1396), .B(n_1384), .Y(n_1463) );
OAI21xp33_ASAP7_75t_L g1464 ( .A1(n_1399), .A2(n_1302), .B(n_1266), .Y(n_1464) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_1396), .B(n_1205), .Y(n_1465) );
NAND2xp5_ASAP7_75t_L g1466 ( .A(n_1384), .B(n_1327), .Y(n_1466) );
AND2x2_ASAP7_75t_L g1467 ( .A(n_1389), .B(n_1323), .Y(n_1467) );
NAND2xp5_ASAP7_75t_L g1468 ( .A(n_1394), .B(n_1314), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1405), .B(n_1314), .Y(n_1469) );
INVx4_ASAP7_75t_L g1470 ( .A(n_1348), .Y(n_1470) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1337), .Y(n_1471) );
AND2x2_ASAP7_75t_L g1472 ( .A(n_1420), .B(n_1310), .Y(n_1472) );
INVx4_ASAP7_75t_L g1473 ( .A(n_1361), .Y(n_1473) );
AND2x2_ASAP7_75t_L g1474 ( .A(n_1420), .B(n_1310), .Y(n_1474) );
INVxp67_ASAP7_75t_L g1475 ( .A(n_1354), .Y(n_1475) );
AND3x1_ASAP7_75t_L g1476 ( .A(n_1379), .B(n_1286), .C(n_1249), .Y(n_1476) );
BUFx2_ASAP7_75t_L g1477 ( .A(n_1361), .Y(n_1477) );
AND2x4_ASAP7_75t_L g1478 ( .A(n_1385), .B(n_1291), .Y(n_1478) );
NAND2xp5_ASAP7_75t_L g1479 ( .A(n_1345), .B(n_1330), .Y(n_1479) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1360), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1481 ( .A(n_1381), .B(n_1330), .Y(n_1481) );
INVxp33_ASAP7_75t_L g1482 ( .A(n_1368), .Y(n_1482) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1371), .Y(n_1483) );
OR2x2_ASAP7_75t_L g1484 ( .A(n_1374), .B(n_1303), .Y(n_1484) );
AND2x4_ASAP7_75t_L g1485 ( .A(n_1385), .B(n_1247), .Y(n_1485) );
OR2x2_ASAP7_75t_SL g1486 ( .A(n_1385), .B(n_1372), .Y(n_1486) );
HB1xp67_ASAP7_75t_L g1487 ( .A(n_1343), .Y(n_1487) );
CKINVDCx16_ASAP7_75t_R g1488 ( .A(n_1361), .Y(n_1488) );
AND2x2_ASAP7_75t_L g1489 ( .A(n_1381), .B(n_1382), .Y(n_1489) );
BUFx3_ASAP7_75t_L g1490 ( .A(n_1386), .Y(n_1490) );
OR2x2_ASAP7_75t_L g1491 ( .A(n_1369), .B(n_1404), .Y(n_1491) );
HB1xp67_ASAP7_75t_L g1492 ( .A(n_1352), .Y(n_1492) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1382), .B(n_1356), .Y(n_1493) );
NAND2xp5_ASAP7_75t_L g1494 ( .A(n_1406), .B(n_1377), .Y(n_1494) );
INVx1_ASAP7_75t_SL g1495 ( .A(n_1367), .Y(n_1495) );
BUFx2_ASAP7_75t_L g1496 ( .A(n_1373), .Y(n_1496) );
AND2x2_ASAP7_75t_L g1497 ( .A(n_1397), .B(n_1401), .Y(n_1497) );
AND2x2_ASAP7_75t_L g1498 ( .A(n_1397), .B(n_1401), .Y(n_1498) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1380), .Y(n_1499) );
AND2x2_ASAP7_75t_L g1500 ( .A(n_1380), .B(n_1338), .Y(n_1500) );
OR2x2_ASAP7_75t_L g1501 ( .A(n_1357), .B(n_1358), .Y(n_1501) );
AND2x2_ASAP7_75t_L g1502 ( .A(n_1338), .B(n_1339), .Y(n_1502) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1370), .Y(n_1503) );
AND2x2_ASAP7_75t_L g1504 ( .A(n_1339), .B(n_1417), .Y(n_1504) );
AND2x2_ASAP7_75t_L g1505 ( .A(n_1417), .B(n_1418), .Y(n_1505) );
NAND2xp5_ASAP7_75t_L g1506 ( .A(n_1399), .B(n_1411), .Y(n_1506) );
AND2x2_ASAP7_75t_L g1507 ( .A(n_1418), .B(n_1344), .Y(n_1507) );
AND2x2_ASAP7_75t_L g1508 ( .A(n_1344), .B(n_1408), .Y(n_1508) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1391), .Y(n_1509) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_1344), .B(n_1408), .Y(n_1510) );
NAND2xp5_ASAP7_75t_L g1511 ( .A(n_1375), .B(n_1403), .Y(n_1511) );
NAND2xp5_ASAP7_75t_SL g1512 ( .A(n_1423), .B(n_1409), .Y(n_1512) );
NOR2xp33_ASAP7_75t_L g1513 ( .A(n_1495), .B(n_1390), .Y(n_1513) );
INVx2_ASAP7_75t_L g1514 ( .A(n_1438), .Y(n_1514) );
AND2x4_ASAP7_75t_L g1515 ( .A(n_1473), .B(n_1477), .Y(n_1515) );
INVx4_ASAP7_75t_L g1516 ( .A(n_1462), .Y(n_1516) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1443), .Y(n_1517) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1444), .Y(n_1518) );
OR2x2_ASAP7_75t_L g1519 ( .A(n_1463), .B(n_1383), .Y(n_1519) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1446), .Y(n_1520) );
INVx2_ASAP7_75t_SL g1521 ( .A(n_1496), .Y(n_1521) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1501), .Y(n_1522) );
AND2x2_ASAP7_75t_L g1523 ( .A(n_1497), .B(n_1415), .Y(n_1523) );
AND2x4_ASAP7_75t_L g1524 ( .A(n_1473), .B(n_1365), .Y(n_1524) );
AND2x2_ASAP7_75t_L g1525 ( .A(n_1497), .B(n_1498), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1498), .B(n_1415), .Y(n_1526) );
OR2x2_ASAP7_75t_L g1527 ( .A(n_1463), .B(n_1388), .Y(n_1527) );
OAI22xp5_ASAP7_75t_L g1528 ( .A1(n_1488), .A2(n_1428), .B1(n_1423), .B2(n_1427), .Y(n_1528) );
OR2x2_ASAP7_75t_L g1529 ( .A(n_1502), .B(n_1346), .Y(n_1529) );
AND2x2_ASAP7_75t_L g1530 ( .A(n_1500), .B(n_1392), .Y(n_1530) );
AOI211xp5_ASAP7_75t_L g1531 ( .A1(n_1482), .A2(n_1402), .B(n_1430), .C(n_1379), .Y(n_1531) );
AND2x2_ASAP7_75t_L g1532 ( .A(n_1504), .B(n_1393), .Y(n_1532) );
NAND2xp5_ASAP7_75t_L g1533 ( .A(n_1505), .B(n_1378), .Y(n_1533) );
INVx2_ASAP7_75t_L g1534 ( .A(n_1438), .Y(n_1534) );
NAND2xp5_ASAP7_75t_L g1535 ( .A(n_1505), .B(n_1378), .Y(n_1535) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1501), .Y(n_1536) );
INVx2_ASAP7_75t_L g1537 ( .A(n_1442), .Y(n_1537) );
INVx4_ASAP7_75t_L g1538 ( .A(n_1462), .Y(n_1538) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_1504), .B(n_1393), .Y(n_1539) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1509), .Y(n_1540) );
AND2x2_ASAP7_75t_L g1541 ( .A(n_1493), .B(n_1431), .Y(n_1541) );
INVxp67_ASAP7_75t_SL g1542 ( .A(n_1492), .Y(n_1542) );
OR2x2_ASAP7_75t_L g1543 ( .A(n_1491), .B(n_1341), .Y(n_1543) );
NAND2xp5_ASAP7_75t_L g1544 ( .A(n_1499), .B(n_1432), .Y(n_1544) );
NAND2xp5_ASAP7_75t_L g1545 ( .A(n_1499), .B(n_1433), .Y(n_1545) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1503), .Y(n_1546) );
NAND4xp25_ASAP7_75t_L g1547 ( .A(n_1506), .B(n_1428), .C(n_1429), .D(n_1427), .Y(n_1547) );
OR2x2_ASAP7_75t_L g1548 ( .A(n_1491), .B(n_1346), .Y(n_1548) );
OR2x2_ASAP7_75t_L g1549 ( .A(n_1493), .B(n_1347), .Y(n_1549) );
OR2x2_ASAP7_75t_L g1550 ( .A(n_1471), .B(n_1347), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1551 ( .A(n_1508), .B(n_1349), .Y(n_1551) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1452), .Y(n_1552) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1452), .Y(n_1553) );
AND2x2_ASAP7_75t_L g1554 ( .A(n_1508), .B(n_1349), .Y(n_1554) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1453), .Y(n_1555) );
OR2x6_ASAP7_75t_L g1556 ( .A(n_1473), .B(n_1379), .Y(n_1556) );
AND2x2_ASAP7_75t_L g1557 ( .A(n_1510), .B(n_1353), .Y(n_1557) );
AND2x2_ASAP7_75t_L g1558 ( .A(n_1510), .B(n_1353), .Y(n_1558) );
NAND2xp5_ASAP7_75t_L g1559 ( .A(n_1489), .B(n_1425), .Y(n_1559) );
AND2x2_ASAP7_75t_L g1560 ( .A(n_1489), .B(n_1376), .Y(n_1560) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1453), .Y(n_1561) );
AND2x2_ASAP7_75t_L g1562 ( .A(n_1487), .B(n_1376), .Y(n_1562) );
AND2x4_ASAP7_75t_L g1563 ( .A(n_1477), .B(n_1365), .Y(n_1563) );
AND2x2_ASAP7_75t_L g1564 ( .A(n_1448), .B(n_1436), .Y(n_1564) );
INVxp67_ASAP7_75t_SL g1565 ( .A(n_1451), .Y(n_1565) );
NAND2xp5_ASAP7_75t_L g1566 ( .A(n_1454), .B(n_1425), .Y(n_1566) );
OR2x2_ASAP7_75t_L g1567 ( .A(n_1483), .B(n_1342), .Y(n_1567) );
OR2x2_ASAP7_75t_L g1568 ( .A(n_1458), .B(n_1342), .Y(n_1568) );
NOR2xp67_ASAP7_75t_L g1569 ( .A(n_1470), .B(n_1409), .Y(n_1569) );
AND2x2_ASAP7_75t_L g1570 ( .A(n_1448), .B(n_1373), .Y(n_1570) );
AND2x2_ASAP7_75t_L g1571 ( .A(n_1480), .B(n_1387), .Y(n_1571) );
INVx2_ASAP7_75t_SL g1572 ( .A(n_1496), .Y(n_1572) );
HB1xp67_ASAP7_75t_L g1573 ( .A(n_1459), .Y(n_1573) );
NAND3xp33_ASAP7_75t_L g1574 ( .A(n_1547), .B(n_1531), .C(n_1542), .Y(n_1574) );
HB1xp67_ASAP7_75t_L g1575 ( .A(n_1542), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1576 ( .A(n_1525), .B(n_1469), .Y(n_1576) );
NAND2xp5_ASAP7_75t_L g1577 ( .A(n_1522), .B(n_1450), .Y(n_1577) );
INVx2_ASAP7_75t_L g1578 ( .A(n_1514), .Y(n_1578) );
AND2x4_ASAP7_75t_L g1579 ( .A(n_1524), .B(n_1478), .Y(n_1579) );
AOI211xp5_ASAP7_75t_L g1580 ( .A1(n_1528), .A2(n_1482), .B(n_1512), .C(n_1460), .Y(n_1580) );
INVxp67_ASAP7_75t_SL g1581 ( .A(n_1573), .Y(n_1581) );
NAND2xp5_ASAP7_75t_L g1582 ( .A(n_1536), .B(n_1511), .Y(n_1582) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1552), .Y(n_1583) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1553), .Y(n_1584) );
NAND2xp5_ASAP7_75t_L g1585 ( .A(n_1533), .B(n_1445), .Y(n_1585) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1555), .Y(n_1586) );
NOR2x1p5_ASAP7_75t_SL g1587 ( .A(n_1514), .B(n_1451), .Y(n_1587) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1561), .Y(n_1588) );
AND2x2_ASAP7_75t_L g1589 ( .A(n_1551), .B(n_1469), .Y(n_1589) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1554), .B(n_1507), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1557), .B(n_1507), .Y(n_1591) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1517), .Y(n_1592) );
OR2x2_ASAP7_75t_L g1593 ( .A(n_1559), .B(n_1466), .Y(n_1593) );
HB1xp67_ASAP7_75t_L g1594 ( .A(n_1521), .Y(n_1594) );
NAND3xp33_ASAP7_75t_L g1595 ( .A(n_1546), .B(n_1457), .C(n_1475), .Y(n_1595) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1518), .Y(n_1596) );
INVx1_ASAP7_75t_L g1597 ( .A(n_1520), .Y(n_1597) );
AND2x4_ASAP7_75t_L g1598 ( .A(n_1563), .B(n_1447), .Y(n_1598) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1540), .Y(n_1599) );
INVx1_ASAP7_75t_SL g1600 ( .A(n_1516), .Y(n_1600) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1565), .Y(n_1601) );
INVx2_ASAP7_75t_L g1602 ( .A(n_1534), .Y(n_1602) );
NAND2xp5_ASAP7_75t_L g1603 ( .A(n_1533), .B(n_1465), .Y(n_1603) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1558), .B(n_1530), .Y(n_1604) );
INVxp67_ASAP7_75t_L g1605 ( .A(n_1513), .Y(n_1605) );
INVx2_ASAP7_75t_SL g1606 ( .A(n_1516), .Y(n_1606) );
INVx3_ASAP7_75t_L g1607 ( .A(n_1516), .Y(n_1607) );
INVx2_ASAP7_75t_L g1608 ( .A(n_1534), .Y(n_1608) );
INVx2_ASAP7_75t_L g1609 ( .A(n_1537), .Y(n_1609) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1565), .Y(n_1610) );
AND2x2_ASAP7_75t_L g1611 ( .A(n_1532), .B(n_1455), .Y(n_1611) );
INVx2_ASAP7_75t_L g1612 ( .A(n_1537), .Y(n_1612) );
AOI222xp33_ASAP7_75t_L g1613 ( .A1(n_1574), .A2(n_1528), .B1(n_1513), .B2(n_1535), .C1(n_1494), .C2(n_1456), .Y(n_1613) );
AOI221xp5_ASAP7_75t_L g1614 ( .A1(n_1605), .A2(n_1535), .B1(n_1526), .B2(n_1523), .C(n_1559), .Y(n_1614) );
INVx2_ASAP7_75t_L g1615 ( .A(n_1578), .Y(n_1615) );
INVx2_ASAP7_75t_L g1616 ( .A(n_1578), .Y(n_1616) );
NOR2x1_ASAP7_75t_L g1617 ( .A(n_1607), .B(n_1538), .Y(n_1617) );
NOR3xp33_ASAP7_75t_L g1618 ( .A(n_1595), .B(n_1439), .C(n_1437), .Y(n_1618) );
INVx1_ASAP7_75t_L g1619 ( .A(n_1592), .Y(n_1619) );
OR2x2_ASAP7_75t_L g1620 ( .A(n_1593), .B(n_1549), .Y(n_1620) );
OAI21xp5_ASAP7_75t_L g1621 ( .A1(n_1600), .A2(n_1538), .B(n_1440), .Y(n_1621) );
INVx2_ASAP7_75t_L g1622 ( .A(n_1602), .Y(n_1622) );
OAI22xp33_ASAP7_75t_L g1623 ( .A1(n_1607), .A2(n_1470), .B1(n_1569), .B2(n_1556), .Y(n_1623) );
NAND3xp33_ASAP7_75t_L g1624 ( .A(n_1580), .B(n_1572), .C(n_1521), .Y(n_1624) );
OAI221xp5_ASAP7_75t_L g1625 ( .A1(n_1606), .A2(n_1464), .B1(n_1572), .B2(n_1545), .C(n_1544), .Y(n_1625) );
XNOR2x2_ASAP7_75t_L g1626 ( .A(n_1601), .B(n_1410), .Y(n_1626) );
INVx2_ASAP7_75t_L g1627 ( .A(n_1602), .Y(n_1627) );
INVx2_ASAP7_75t_L g1628 ( .A(n_1608), .Y(n_1628) );
INVx2_ASAP7_75t_L g1629 ( .A(n_1608), .Y(n_1629) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1592), .Y(n_1630) );
AND2x2_ASAP7_75t_L g1631 ( .A(n_1576), .B(n_1541), .Y(n_1631) );
O2A1O1Ixp33_ASAP7_75t_L g1632 ( .A1(n_1606), .A2(n_1386), .B(n_1490), .C(n_1426), .Y(n_1632) );
AOI221xp5_ASAP7_75t_L g1633 ( .A1(n_1585), .A2(n_1571), .B1(n_1545), .B2(n_1566), .C(n_1539), .Y(n_1633) );
INVx3_ASAP7_75t_L g1634 ( .A(n_1579), .Y(n_1634) );
OA21x2_ASAP7_75t_L g1635 ( .A1(n_1610), .A2(n_1468), .B(n_1481), .Y(n_1635) );
AOI221xp5_ASAP7_75t_L g1636 ( .A1(n_1582), .A2(n_1560), .B1(n_1564), .B2(n_1527), .C(n_1519), .Y(n_1636) );
NAND2xp5_ASAP7_75t_L g1637 ( .A(n_1576), .B(n_1465), .Y(n_1637) );
AOI21xp33_ASAP7_75t_SL g1638 ( .A1(n_1575), .A2(n_1556), .B(n_1515), .Y(n_1638) );
OAI21xp33_ASAP7_75t_L g1639 ( .A1(n_1613), .A2(n_1587), .B(n_1593), .Y(n_1639) );
AOI221xp5_ASAP7_75t_L g1640 ( .A1(n_1614), .A2(n_1577), .B1(n_1599), .B2(n_1596), .C(n_1597), .Y(n_1640) );
OAI221xp5_ASAP7_75t_L g1641 ( .A1(n_1621), .A2(n_1594), .B1(n_1610), .B2(n_1581), .C(n_1599), .Y(n_1641) );
AOI211x1_ASAP7_75t_L g1642 ( .A1(n_1624), .A2(n_1604), .B(n_1591), .C(n_1590), .Y(n_1642) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1620), .Y(n_1643) );
AOI21xp33_ASAP7_75t_SL g1644 ( .A1(n_1632), .A2(n_1556), .B(n_1598), .Y(n_1644) );
AOI22xp5_ASAP7_75t_L g1645 ( .A1(n_1618), .A2(n_1579), .B1(n_1598), .B2(n_1563), .Y(n_1645) );
AOI22xp5_ASAP7_75t_L g1646 ( .A1(n_1633), .A2(n_1579), .B1(n_1598), .B2(n_1563), .Y(n_1646) );
AOI22xp5_ASAP7_75t_L g1647 ( .A1(n_1617), .A2(n_1579), .B1(n_1562), .B2(n_1603), .Y(n_1647) );
OAI22xp5_ASAP7_75t_L g1648 ( .A1(n_1636), .A2(n_1486), .B1(n_1529), .B2(n_1604), .Y(n_1648) );
AOI221xp5_ASAP7_75t_L g1649 ( .A1(n_1625), .A2(n_1586), .B1(n_1583), .B2(n_1588), .C(n_1584), .Y(n_1649) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1634), .B(n_1589), .Y(n_1650) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1619), .Y(n_1651) );
AOI221xp5_ASAP7_75t_L g1652 ( .A1(n_1638), .A2(n_1586), .B1(n_1583), .B2(n_1588), .C(n_1584), .Y(n_1652) );
AOI211xp5_ASAP7_75t_L g1653 ( .A1(n_1623), .A2(n_1570), .B(n_1515), .C(n_1524), .Y(n_1653) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1630), .Y(n_1654) );
OAI221xp5_ASAP7_75t_L g1655 ( .A1(n_1635), .A2(n_1476), .B1(n_1484), .B2(n_1548), .C(n_1543), .Y(n_1655) );
AOI21xp5_ASAP7_75t_L g1656 ( .A1(n_1635), .A2(n_1524), .B(n_1387), .Y(n_1656) );
XOR2x2_ASAP7_75t_L g1657 ( .A(n_1626), .B(n_1611), .Y(n_1657) );
AOI21xp5_ASAP7_75t_L g1658 ( .A1(n_1635), .A2(n_1398), .B(n_1609), .Y(n_1658) );
O2A1O1Ixp33_ASAP7_75t_L g1659 ( .A1(n_1626), .A2(n_1419), .B(n_1429), .C(n_1413), .Y(n_1659) );
AOI211xp5_ASAP7_75t_L g1660 ( .A1(n_1631), .A2(n_1424), .B(n_1441), .C(n_1435), .Y(n_1660) );
INVx1_ASAP7_75t_L g1661 ( .A(n_1615), .Y(n_1661) );
OAI211xp5_ASAP7_75t_L g1662 ( .A1(n_1637), .A2(n_1424), .B(n_1484), .C(n_1481), .Y(n_1662) );
OAI221xp5_ASAP7_75t_L g1663 ( .A1(n_1616), .A2(n_1550), .B1(n_1567), .B2(n_1568), .C(n_1461), .Y(n_1663) );
NAND4xp75_ASAP7_75t_L g1664 ( .A(n_1642), .B(n_1646), .C(n_1645), .D(n_1649), .Y(n_1664) );
NOR3xp33_ASAP7_75t_L g1665 ( .A(n_1639), .B(n_1644), .C(n_1641), .Y(n_1665) );
AND4x1_ASAP7_75t_L g1666 ( .A(n_1653), .B(n_1659), .C(n_1660), .D(n_1652), .Y(n_1666) );
A2O1A1Ixp33_ASAP7_75t_L g1667 ( .A1(n_1648), .A2(n_1662), .B(n_1658), .C(n_1656), .Y(n_1667) );
OAI211xp5_ASAP7_75t_L g1668 ( .A1(n_1655), .A2(n_1640), .B(n_1647), .C(n_1660), .Y(n_1668) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1643), .Y(n_1669) );
NOR3xp33_ASAP7_75t_L g1670 ( .A(n_1663), .B(n_1654), .C(n_1651), .Y(n_1670) );
NAND4xp25_ASAP7_75t_L g1671 ( .A(n_1650), .B(n_1441), .C(n_1657), .D(n_1414), .Y(n_1671) );
AND2x2_ASAP7_75t_L g1672 ( .A(n_1665), .B(n_1661), .Y(n_1672) );
NAND3xp33_ASAP7_75t_SL g1673 ( .A(n_1666), .B(n_1667), .C(n_1668), .Y(n_1673) );
NOR3xp33_ASAP7_75t_L g1674 ( .A(n_1664), .B(n_1412), .C(n_1628), .Y(n_1674) );
OAI211xp5_ASAP7_75t_SL g1675 ( .A1(n_1669), .A2(n_1629), .B(n_1628), .C(n_1627), .Y(n_1675) );
CKINVDCx12_ASAP7_75t_R g1676 ( .A(n_1671), .Y(n_1676) );
NOR2xp33_ASAP7_75t_L g1677 ( .A(n_1673), .B(n_1670), .Y(n_1677) );
AND3x1_ASAP7_75t_L g1678 ( .A(n_1674), .B(n_1398), .C(n_1627), .Y(n_1678) );
NAND2xp5_ASAP7_75t_L g1679 ( .A(n_1672), .B(n_1622), .Y(n_1679) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1676), .Y(n_1680) );
INVx2_ASAP7_75t_L g1681 ( .A(n_1680), .Y(n_1681) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1679), .Y(n_1682) );
NAND2x1p5_ASAP7_75t_L g1683 ( .A(n_1678), .B(n_1486), .Y(n_1683) );
NAND2xp5_ASAP7_75t_SL g1684 ( .A(n_1677), .B(n_1675), .Y(n_1684) );
INVx2_ASAP7_75t_L g1685 ( .A(n_1681), .Y(n_1685) );
INVx2_ASAP7_75t_L g1686 ( .A(n_1682), .Y(n_1686) );
NAND2xp5_ASAP7_75t_L g1687 ( .A(n_1682), .B(n_1587), .Y(n_1687) );
HB1xp67_ASAP7_75t_L g1688 ( .A(n_1685), .Y(n_1688) );
AOI21xp5_ASAP7_75t_L g1689 ( .A1(n_1686), .A2(n_1684), .B(n_1683), .Y(n_1689) );
NAND2xp5_ASAP7_75t_L g1690 ( .A(n_1687), .B(n_1612), .Y(n_1690) );
OAI21xp5_ASAP7_75t_L g1691 ( .A1(n_1689), .A2(n_1479), .B(n_1485), .Y(n_1691) );
AOI22xp5_ASAP7_75t_L g1692 ( .A1(n_1688), .A2(n_1478), .B1(n_1472), .B2(n_1474), .Y(n_1692) );
AOI21xp5_ASAP7_75t_L g1693 ( .A1(n_1690), .A2(n_1485), .B(n_1478), .Y(n_1693) );
OAI21xp5_ASAP7_75t_L g1694 ( .A1(n_1691), .A2(n_1485), .B(n_1421), .Y(n_1694) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1692), .Y(n_1695) );
OAI21xp5_ASAP7_75t_L g1696 ( .A1(n_1693), .A2(n_1421), .B(n_1422), .Y(n_1696) );
AO21x2_ASAP7_75t_L g1697 ( .A1(n_1695), .A2(n_1696), .B(n_1694), .Y(n_1697) );
AOI21xp33_ASAP7_75t_SL g1698 ( .A1(n_1697), .A2(n_1449), .B(n_1467), .Y(n_1698) );
endmodule