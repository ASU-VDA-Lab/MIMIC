module real_aes_9150_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1016;
wire n_908;
wire n_376;
wire n_571;
wire n_1034;
wire n_694;
wire n_491;
wire n_549;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_551;
wire n_666;
wire n_537;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_932;
wire n_399;
wire n_1021;
wire n_700;
wire n_948;
wire n_958;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_1040;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_994;
wire n_578;
wire n_495;
wire n_892;
wire n_370;
wire n_744;
wire n_384;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_875;
wire n_467;
wire n_951;
wire n_992;
wire n_774;
wire n_813;
wire n_791;
wire n_981;
wire n_976;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_726;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_656;
wire n_532;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_973;
wire n_504;
wire n_960;
wire n_671;
wire n_725;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1017;
wire n_1013;
wire n_936;
wire n_610;
wire n_581;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_1006;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_1041;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1000;
wire n_1003;
wire n_366;
wire n_727;
wire n_1014;
wire n_397;
wire n_749;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_354;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_831;
wire n_487;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_968;
wire n_650;
wire n_710;
wire n_743;
wire n_393;
wire n_652;
wire n_703;
wire n_823;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1024;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_0), .A2(n_144), .B1(n_516), .B2(n_518), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_1), .A2(n_149), .B1(n_453), .B2(n_457), .Y(n_452) );
INVx1_ASAP7_75t_L g505 ( .A(n_2), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_3), .A2(n_313), .B1(n_447), .B2(n_654), .Y(n_692) );
AOI22xp33_ASAP7_75t_SL g827 ( .A1(n_4), .A2(n_114), .B1(n_518), .B2(n_711), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_5), .Y(n_593) );
AOI211xp5_ASAP7_75t_L g350 ( .A1(n_6), .A2(n_351), .B(n_359), .C(n_986), .Y(n_350) );
AOI222xp33_ASAP7_75t_L g644 ( .A1(n_7), .A2(n_169), .B1(n_268), .B2(n_479), .C1(n_554), .C2(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_8), .A2(n_85), .B1(n_668), .B2(n_682), .Y(n_1000) );
CKINVDCx20_ASAP7_75t_R g1033 ( .A(n_9), .Y(n_1033) );
AO22x2_ASAP7_75t_L g374 ( .A1(n_10), .A2(n_194), .B1(n_375), .B2(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g984 ( .A(n_10), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_11), .A2(n_133), .B1(n_600), .B2(n_629), .Y(n_705) );
AOI222xp33_ASAP7_75t_L g832 ( .A1(n_12), .A2(n_293), .B1(n_304), .B2(n_551), .C1(n_587), .C2(n_588), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_13), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_14), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_15), .A2(n_43), .B1(n_528), .B2(n_530), .Y(n_527) );
AOI22xp33_ASAP7_75t_SL g923 ( .A1(n_16), .A2(n_103), .B1(n_605), .B2(n_637), .Y(n_923) );
AOI22xp33_ASAP7_75t_SL g914 ( .A1(n_17), .A2(n_254), .B1(n_587), .B2(n_588), .Y(n_914) );
INVx1_ASAP7_75t_L g500 ( .A(n_18), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_19), .A2(n_286), .B1(n_627), .B2(n_763), .Y(n_881) );
AOI22xp5_ASAP7_75t_SL g655 ( .A1(n_20), .A2(n_172), .B1(n_457), .B2(n_656), .Y(n_655) );
AOI22xp33_ASAP7_75t_SL g921 ( .A1(n_21), .A2(n_234), .B1(n_599), .B2(n_876), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_22), .A2(n_77), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp33_ASAP7_75t_SL g1003 ( .A1(n_23), .A2(n_181), .B1(n_875), .B2(n_876), .Y(n_1003) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_24), .A2(n_173), .B1(n_399), .B2(n_480), .Y(n_506) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_25), .A2(n_94), .B1(n_618), .B2(n_619), .C(n_621), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_26), .A2(n_136), .B1(n_742), .B2(n_831), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_27), .A2(n_96), .B1(n_488), .B2(n_489), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_28), .A2(n_289), .B1(n_530), .B2(n_768), .Y(n_767) );
AOI22xp33_ASAP7_75t_SL g1002 ( .A1(n_29), .A2(n_118), .B1(n_561), .B2(n_740), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_30), .A2(n_221), .B1(n_518), .B2(n_544), .Y(n_543) );
AO22x2_ASAP7_75t_L g378 ( .A1(n_31), .A2(n_102), .B1(n_375), .B2(n_379), .Y(n_378) );
AOI22xp33_ASAP7_75t_SL g689 ( .A1(n_32), .A2(n_240), .B1(n_526), .B2(n_600), .Y(n_689) );
AOI222xp33_ASAP7_75t_L g715 ( .A1(n_33), .A2(n_170), .B1(n_267), .B2(n_477), .C1(n_480), .C2(n_716), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_34), .A2(n_281), .B1(n_432), .B2(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_35), .B(n_999), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_36), .A2(n_232), .B1(n_604), .B2(n_742), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_37), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_38), .A2(n_179), .B1(n_512), .B2(n_639), .C(n_641), .Y(n_638) );
AOI22xp33_ASAP7_75t_SL g920 ( .A1(n_39), .A2(n_104), .B1(n_597), .B2(n_619), .Y(n_920) );
AOI22xp33_ASAP7_75t_SL g731 ( .A1(n_40), .A2(n_109), .B1(n_716), .B2(n_732), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_41), .A2(n_81), .B1(n_526), .B2(n_694), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g880 ( .A(n_42), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_44), .A2(n_124), .B1(n_488), .B2(n_748), .Y(n_843) );
INVx1_ASAP7_75t_L g855 ( .A(n_45), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_46), .A2(n_90), .B1(n_426), .B2(n_432), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_47), .A2(n_249), .B1(n_748), .B2(n_749), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_48), .A2(n_200), .B1(n_496), .B2(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_49), .A2(n_79), .B1(n_564), .B2(n_601), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_50), .A2(n_280), .B1(n_494), .B2(n_496), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_51), .B(n_477), .Y(n_1031) );
INVx1_ASAP7_75t_L g635 ( .A(n_52), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_53), .A2(n_165), .B1(n_544), .B2(n_682), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_54), .A2(n_69), .B1(n_709), .B2(n_773), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_55), .A2(n_336), .B1(n_564), .B2(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_56), .B(n_709), .Y(n_826) );
INVx1_ASAP7_75t_L g695 ( .A(n_57), .Y(n_695) );
AOI22xp33_ASAP7_75t_SL g1005 ( .A1(n_58), .A2(n_348), .B1(n_618), .B2(n_1006), .Y(n_1005) );
AOI22xp33_ASAP7_75t_SL g737 ( .A1(n_59), .A2(n_145), .B1(n_738), .B2(n_740), .Y(n_737) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_60), .A2(n_198), .B1(n_432), .B2(n_694), .Y(n_693) );
AOI22xp33_ASAP7_75t_SL g746 ( .A1(n_61), .A2(n_266), .B1(n_569), .B2(n_694), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_62), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_63), .A2(n_301), .B1(n_441), .B2(n_446), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_64), .A2(n_343), .B1(n_544), .B2(n_716), .Y(n_849) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_65), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_66), .Y(n_885) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_67), .A2(n_229), .B1(n_523), .B2(n_619), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_68), .A2(n_247), .B1(n_518), .B2(n_732), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_70), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_71), .A2(n_224), .B1(n_526), .B2(n_831), .Y(n_962) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_72), .A2(n_92), .B1(n_494), .B2(n_627), .C(n_630), .Y(n_626) );
AO22x2_ASAP7_75t_L g382 ( .A1(n_73), .A2(n_231), .B1(n_375), .B2(n_376), .Y(n_382) );
INVx1_ASAP7_75t_L g981 ( .A(n_73), .Y(n_981) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_74), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_75), .A2(n_88), .B1(n_627), .B2(n_765), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_76), .A2(n_128), .B1(n_548), .B2(n_668), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_78), .A2(n_189), .B1(n_668), .B2(n_669), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_80), .A2(n_250), .B1(n_439), .B2(n_496), .Y(n_607) );
AOI22xp33_ASAP7_75t_SL g686 ( .A1(n_82), .A2(n_242), .B1(n_399), .B2(n_516), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_83), .A2(n_166), .B1(n_666), .B2(n_734), .Y(n_931) );
CKINVDCx20_ASAP7_75t_R g953 ( .A(n_84), .Y(n_953) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_86), .A2(n_339), .B1(n_479), .B2(n_711), .Y(n_710) );
AOI222xp33_ASAP7_75t_L g816 ( .A1(n_87), .A2(n_98), .B1(n_159), .B2(n_588), .C1(n_645), .C2(n_817), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_89), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_91), .A2(n_536), .B1(n_570), .B2(n_571), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_91), .Y(n_570) );
INVx1_ASAP7_75t_L g642 ( .A(n_93), .Y(n_642) );
XOR2x2_ASAP7_75t_L g778 ( .A(n_95), .B(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g671 ( .A(n_97), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_99), .A2(n_246), .B1(n_498), .B2(n_597), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_100), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_101), .A2(n_238), .B1(n_443), .B2(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g985 ( .A(n_102), .Y(n_985) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_105), .A2(n_272), .B1(n_618), .B2(n_660), .Y(n_659) );
XOR2x2_ASAP7_75t_L g909 ( .A(n_106), .B(n_910), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_107), .B(n_791), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_108), .A2(n_244), .B1(n_604), .B2(n_606), .Y(n_603) );
AO22x1_ASAP7_75t_L g758 ( .A1(n_110), .A2(n_759), .B1(n_760), .B2(n_776), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_110), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_111), .A2(n_130), .B1(n_458), .B2(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_112), .B(n_789), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_113), .A2(n_132), .B1(n_480), .B2(n_726), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_115), .A2(n_314), .B1(n_439), .B2(n_447), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_116), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_117), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_119), .A2(n_121), .B1(n_498), .B2(n_597), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_120), .A2(n_616), .B1(n_646), .B2(n_647), .Y(n_615) );
INVx1_ASAP7_75t_L g646 ( .A(n_120), .Y(n_646) );
INVx1_ASAP7_75t_L g631 ( .A(n_122), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_123), .A2(n_143), .B1(n_446), .B2(n_449), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_125), .A2(n_197), .B1(n_437), .B2(n_441), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_126), .A2(n_311), .B1(n_599), .B2(n_802), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_127), .A2(n_140), .B1(n_457), .B2(n_564), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_129), .A2(n_324), .B1(n_749), .B2(n_797), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g889 ( .A(n_131), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_134), .A2(n_274), .B1(n_489), .B2(n_765), .Y(n_822) );
AOI22xp33_ASAP7_75t_SL g598 ( .A1(n_135), .A2(n_220), .B1(n_599), .B2(n_601), .Y(n_598) );
AND2x6_ASAP7_75t_L g353 ( .A(n_137), .B(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g978 ( .A(n_137), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_138), .A2(n_253), .B1(n_453), .B2(n_802), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_139), .A2(n_300), .B1(n_479), .B2(n_480), .Y(n_478) );
AOI22xp33_ASAP7_75t_SL g993 ( .A1(n_141), .A2(n_235), .B1(n_863), .B2(n_994), .Y(n_993) );
CKINVDCx20_ASAP7_75t_R g898 ( .A(n_142), .Y(n_898) );
AOI22xp33_ASAP7_75t_SL g1039 ( .A1(n_146), .A2(n_341), .B1(n_428), .B2(n_749), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_147), .A2(n_294), .B1(n_453), .B2(n_565), .Y(n_960) );
AOI222xp33_ASAP7_75t_L g862 ( .A1(n_148), .A2(n_209), .B1(n_230), .B2(n_393), .C1(n_479), .C2(n_863), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_150), .Y(n_833) );
INVx1_ASAP7_75t_L g864 ( .A(n_151), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_152), .A2(n_279), .B1(n_488), .B2(n_662), .Y(n_928) );
AOI22xp33_ASAP7_75t_SL g1008 ( .A1(n_153), .A2(n_308), .B1(n_606), .B2(n_1009), .Y(n_1008) );
AOI22xp33_ASAP7_75t_SL g1040 ( .A1(n_154), .A2(n_323), .B1(n_831), .B2(n_1041), .Y(n_1040) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_155), .A2(n_326), .B1(n_491), .B2(n_523), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_156), .A2(n_284), .B1(n_606), .B2(n_662), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g943 ( .A(n_157), .Y(n_943) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_158), .A2(n_216), .B1(n_453), .B2(n_800), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_160), .A2(n_312), .B1(n_498), .B2(n_499), .Y(n_497) );
AO22x2_ASAP7_75t_L g384 ( .A1(n_161), .A2(n_217), .B1(n_375), .B2(n_379), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g982 ( .A(n_161), .B(n_983), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_162), .A2(n_186), .B1(n_450), .B2(n_802), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_163), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g958 ( .A(n_164), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_167), .A2(n_338), .B1(n_800), .B2(n_936), .Y(n_935) );
INVx1_ASAP7_75t_L g992 ( .A(n_168), .Y(n_992) );
CKINVDCx20_ASAP7_75t_R g913 ( .A(n_171), .Y(n_913) );
AOI222xp33_ASAP7_75t_L g775 ( .A1(n_174), .A2(n_299), .B1(n_307), .B2(n_399), .C1(n_554), .C2(n_645), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_175), .B(n_407), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_176), .A2(n_223), .B1(n_428), .B2(n_765), .Y(n_934) );
XOR2x2_ASAP7_75t_L g803 ( .A(n_177), .B(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_178), .A2(n_277), .B1(n_665), .B2(n_666), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_180), .Y(n_717) );
INVx1_ASAP7_75t_L g857 ( .A(n_182), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_183), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_184), .A2(n_273), .B1(n_509), .B2(n_665), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_185), .B(n_665), .Y(n_684) );
AOI22xp33_ASAP7_75t_SL g1036 ( .A1(n_187), .A2(n_210), .B1(n_450), .B2(n_797), .Y(n_1036) );
AOI22xp33_ASAP7_75t_SL g1037 ( .A1(n_188), .A2(n_206), .B1(n_600), .B2(n_802), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_190), .A2(n_237), .B1(n_447), .B2(n_491), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_191), .B(n_666), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_192), .A2(n_262), .B1(n_619), .B2(n_811), .Y(n_810) );
AOI22xp33_ASAP7_75t_SL g681 ( .A1(n_193), .A2(n_214), .B1(n_407), .B2(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_195), .A2(n_252), .B1(n_523), .B2(n_561), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_196), .A2(n_264), .B1(n_544), .B2(n_817), .Y(n_918) );
CKINVDCx20_ASAP7_75t_R g942 ( .A(n_199), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_201), .A2(n_337), .B1(n_458), .B2(n_654), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_202), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_203), .Y(n_727) );
INVx1_ASAP7_75t_L g1021 ( .A(n_204), .Y(n_1021) );
OA22x2_ASAP7_75t_L g1022 ( .A1(n_204), .A2(n_1021), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
INVx1_ASAP7_75t_L g852 ( .A(n_205), .Y(n_852) );
INVx1_ASAP7_75t_L g643 ( .A(n_207), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_208), .A2(n_303), .B1(n_479), .B2(n_711), .Y(n_807) );
AOI222xp33_ASAP7_75t_L g937 ( .A1(n_211), .A2(n_315), .B1(n_328), .B2(n_393), .C1(n_399), .C2(n_554), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_212), .A2(n_347), .B1(n_639), .B2(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g358 ( .A(n_213), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_215), .A2(n_248), .B1(n_407), .B2(n_785), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_218), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_219), .Y(n_873) );
XNOR2xp5_ASAP7_75t_L g719 ( .A(n_222), .B(n_720), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_225), .A2(n_575), .B1(n_576), .B2(n_608), .Y(n_574) );
CKINVDCx14_ASAP7_75t_R g608 ( .A(n_225), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g1028 ( .A(n_226), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_227), .A2(n_269), .B1(n_480), .B2(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_228), .A2(n_333), .B1(n_426), .B2(n_763), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g1027 ( .A(n_233), .Y(n_1027) );
INVx1_ASAP7_75t_L g484 ( .A(n_236), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_239), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_241), .Y(n_581) );
AOI22xp33_ASAP7_75t_SL g924 ( .A1(n_243), .A2(n_346), .B1(n_437), .B2(n_629), .Y(n_924) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_245), .Y(n_951) );
INVx1_ASAP7_75t_L g375 ( .A(n_251), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_251), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_255), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_256), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_257), .A2(n_335), .B1(n_875), .B2(n_876), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_258), .B(n_709), .Y(n_917) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_259), .Y(n_385) );
INVx1_ASAP7_75t_L g625 ( .A(n_260), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_261), .B(n_509), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_263), .A2(n_868), .B1(n_901), .B2(n_902), .Y(n_867) );
INVx1_ASAP7_75t_L g901 ( .A(n_263), .Y(n_901) );
CKINVDCx20_ASAP7_75t_R g949 ( .A(n_265), .Y(n_949) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_270), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g987 ( .A1(n_271), .A2(n_988), .B1(n_989), .B2(n_1010), .Y(n_987) );
CKINVDCx20_ASAP7_75t_R g1010 ( .A(n_271), .Y(n_1010) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_275), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_276), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_278), .B(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_282), .A2(n_345), .B1(n_510), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_283), .A2(n_316), .B1(n_964), .B2(n_966), .Y(n_963) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_285), .Y(n_959) );
AND2x2_ASAP7_75t_L g357 ( .A(n_287), .B(n_358), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g878 ( .A(n_288), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_290), .Y(n_397) );
INVx1_ASAP7_75t_L g354 ( .A(n_291), .Y(n_354) );
INVx1_ASAP7_75t_L g674 ( .A(n_292), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_295), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_296), .A2(n_302), .B1(n_432), .B2(n_654), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_297), .Y(n_475) );
INVx1_ASAP7_75t_L g860 ( .A(n_298), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_305), .Y(n_416) );
INVx1_ASAP7_75t_L g622 ( .A(n_306), .Y(n_622) );
AOI22xp33_ASAP7_75t_SL g743 ( .A1(n_309), .A2(n_327), .B1(n_453), .B2(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_310), .Y(n_555) );
INVx1_ASAP7_75t_L g846 ( .A(n_317), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g896 ( .A(n_318), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_319), .B(n_509), .Y(n_685) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_320), .A2(n_342), .B1(n_428), .B2(n_499), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_321), .B(n_666), .Y(n_916) );
XOR2x2_ASAP7_75t_L g925 ( .A(n_322), .B(n_926), .Y(n_925) );
AOI22xp5_ASAP7_75t_L g938 ( .A1(n_325), .A2(n_939), .B1(n_967), .B2(n_968), .Y(n_938) );
CKINVDCx20_ASAP7_75t_R g967 ( .A(n_325), .Y(n_967) );
CKINVDCx20_ASAP7_75t_R g891 ( .A(n_329), .Y(n_891) );
CKINVDCx20_ASAP7_75t_R g1034 ( .A(n_330), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_331), .B(n_848), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g954 ( .A(n_332), .Y(n_954) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_334), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g948 ( .A(n_340), .Y(n_948) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_344), .A2(n_366), .B1(n_461), .B2(n_462), .Y(n_365) );
INVx1_ASAP7_75t_L g461 ( .A(n_344), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_349), .Y(n_472) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
HB1xp67_ASAP7_75t_L g977 ( .A(n_354), .Y(n_977) );
OAI21xp5_ASAP7_75t_L g1019 ( .A1(n_355), .A2(n_976), .B(n_1020), .Y(n_1019) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_836), .B1(n_971), .B2(n_972), .C(n_973), .Y(n_359) );
INVx1_ASAP7_75t_L g971 ( .A(n_360), .Y(n_971) );
XNOR2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_613), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_533), .B1(n_611), .B2(n_612), .Y(n_361) );
INVx1_ASAP7_75t_L g611 ( .A(n_362), .Y(n_611) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B1(n_463), .B2(n_464), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g462 ( .A(n_366), .Y(n_462) );
AND2x2_ASAP7_75t_SL g366 ( .A(n_367), .B(n_423), .Y(n_366) );
NOR3xp33_ASAP7_75t_L g367 ( .A(n_368), .B(n_390), .C(n_410), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B1(n_385), .B2(n_386), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g941 ( .A1(n_370), .A2(n_942), .B1(n_943), .B2(n_944), .Y(n_941) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx3_ASAP7_75t_L g471 ( .A(n_371), .Y(n_471) );
INVx2_ASAP7_75t_L g540 ( .A(n_371), .Y(n_540) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_380), .Y(n_371) );
INVx2_ASAP7_75t_L g440 ( .A(n_372), .Y(n_440) );
OR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_378), .Y(n_372) );
AND2x2_ASAP7_75t_L g389 ( .A(n_373), .B(n_378), .Y(n_389) );
AND2x2_ASAP7_75t_L g431 ( .A(n_373), .B(n_403), .Y(n_431) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g394 ( .A(n_374), .B(n_378), .Y(n_394) );
AND2x2_ASAP7_75t_L g404 ( .A(n_374), .B(n_384), .Y(n_404) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_377), .Y(n_379) );
INVx2_ASAP7_75t_L g403 ( .A(n_378), .Y(n_403) );
INVx1_ASAP7_75t_L g460 ( .A(n_378), .Y(n_460) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2x1p5_ASAP7_75t_L g388 ( .A(n_381), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g451 ( .A(n_381), .B(n_431), .Y(n_451) );
AND2x6_ASAP7_75t_L g510 ( .A(n_381), .B(n_389), .Y(n_510) );
AND2x4_ASAP7_75t_L g514 ( .A(n_381), .B(n_440), .Y(n_514) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_L g396 ( .A(n_382), .Y(n_396) );
INVx1_ASAP7_75t_L g402 ( .A(n_382), .Y(n_402) );
INVx1_ASAP7_75t_L g422 ( .A(n_382), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_382), .B(n_384), .Y(n_435) );
AND2x2_ASAP7_75t_L g395 ( .A(n_383), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g430 ( .A(n_384), .B(n_422), .Y(n_430) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g473 ( .A(n_387), .Y(n_473) );
INVx2_ASAP7_75t_L g886 ( .A(n_387), .Y(n_886) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx3_ASAP7_75t_L g583 ( .A(n_388), .Y(n_583) );
AND2x4_ASAP7_75t_L g443 ( .A(n_389), .B(n_395), .Y(n_443) );
AND2x2_ASAP7_75t_L g456 ( .A(n_389), .B(n_430), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_389), .B(n_430), .Y(n_624) );
OAI221xp5_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_397), .B1(n_398), .B2(n_405), .C(n_406), .Y(n_390) );
OAI21xp5_ASAP7_75t_SL g584 ( .A1(n_391), .A2(n_585), .B(n_586), .Y(n_584) );
OAI21xp5_ASAP7_75t_SL g670 ( .A1(n_391), .A2(n_671), .B(n_672), .Y(n_670) );
BUFx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx4_ASAP7_75t_L g551 ( .A(n_392), .Y(n_551) );
INVx4_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx3_ASAP7_75t_L g477 ( .A(n_393), .Y(n_477) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_393), .Y(n_645) );
INVx2_ASAP7_75t_L g679 ( .A(n_393), .Y(n_679) );
INVx2_ASAP7_75t_SL g782 ( .A(n_393), .Y(n_782) );
AND2x6_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g419 ( .A(n_394), .Y(n_419) );
AND2x4_ASAP7_75t_L g518 ( .A(n_394), .B(n_421), .Y(n_518) );
AND2x6_ASAP7_75t_L g439 ( .A(n_395), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g448 ( .A(n_395), .B(n_431), .Y(n_448) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g947 ( .A(n_399), .Y(n_947) );
BUFx4f_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_400), .Y(n_479) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_400), .Y(n_548) );
BUFx2_ASAP7_75t_L g673 ( .A(n_400), .Y(n_673) );
BUFx6f_ASAP7_75t_L g726 ( .A(n_400), .Y(n_726) );
AND2x4_ASAP7_75t_L g400 ( .A(n_401), .B(n_404), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g409 ( .A(n_402), .Y(n_409) );
INVx1_ASAP7_75t_L g415 ( .A(n_403), .Y(n_415) );
AND2x4_ASAP7_75t_L g408 ( .A(n_404), .B(n_409), .Y(n_408) );
NAND2x1p5_ASAP7_75t_L g414 ( .A(n_404), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g516 ( .A(n_404), .B(n_517), .Y(n_516) );
BUFx3_ASAP7_75t_L g893 ( .A(n_407), .Y(n_893) );
INVx2_ASAP7_75t_L g950 ( .A(n_407), .Y(n_950) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx12f_ASAP7_75t_L g480 ( .A(n_408), .Y(n_480) );
INVx1_ASAP7_75t_L g728 ( .A(n_408), .Y(n_728) );
BUFx6f_ASAP7_75t_L g863 ( .A(n_408), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B1(n_416), .B2(n_417), .Y(n_410) );
INVx3_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g897 ( .A(n_413), .Y(n_897) );
INVx4_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx3_ASAP7_75t_L g483 ( .A(n_414), .Y(n_483) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_414), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_414), .A2(n_418), .B1(n_1033), .B2(n_1034), .Y(n_1032) );
AND2x2_ASAP7_75t_L g523 ( .A(n_415), .B(n_434), .Y(n_523) );
BUFx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_418), .A2(n_482), .B1(n_483), .B2(n_484), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_418), .A2(n_591), .B1(n_592), .B2(n_593), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_418), .A2(n_483), .B1(n_642), .B2(n_643), .Y(n_641) );
CKINVDCx16_ASAP7_75t_R g900 ( .A(n_418), .Y(n_900) );
OR2x6_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_444), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_436), .Y(n_424) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g569 ( .A(n_428), .Y(n_569) );
BUFx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx3_ASAP7_75t_L g489 ( .A(n_429), .Y(n_489) );
BUFx3_ASAP7_75t_L g605 ( .A(n_429), .Y(n_605) );
BUFx3_ASAP7_75t_L g654 ( .A(n_429), .Y(n_654) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_430), .B(n_431), .Y(n_634) );
AND2x4_ASAP7_75t_L g433 ( .A(n_431), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g872 ( .A(n_432), .Y(n_872) );
BUFx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g499 ( .A(n_433), .Y(n_499) );
BUFx2_ASAP7_75t_SL g606 ( .A(n_433), .Y(n_606) );
BUFx2_ASAP7_75t_SL g637 ( .A(n_433), .Y(n_637) );
BUFx3_ASAP7_75t_L g749 ( .A(n_433), .Y(n_749) );
BUFx3_ASAP7_75t_L g765 ( .A(n_433), .Y(n_765) );
INVx1_ASAP7_75t_L g812 ( .A(n_433), .Y(n_812) );
BUFx3_ASAP7_75t_L g966 ( .A(n_433), .Y(n_966) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OR2x6_ASAP7_75t_L g459 ( .A(n_435), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx4_ASAP7_75t_L g526 ( .A(n_438), .Y(n_526) );
INVx3_ASAP7_75t_L g859 ( .A(n_438), .Y(n_859) );
INVx4_ASAP7_75t_L g1041 ( .A(n_438), .Y(n_1041) );
INVx11_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx11_ASAP7_75t_L g495 ( .A(n_439), .Y(n_495) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx3_ASAP7_75t_L g496 ( .A(n_442), .Y(n_496) );
INVx2_ASAP7_75t_L g800 ( .A(n_442), .Y(n_800) );
INVx2_ASAP7_75t_L g1009 ( .A(n_442), .Y(n_1009) );
INVx6_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx3_ASAP7_75t_L g629 ( .A(n_443), .Y(n_629) );
BUFx3_ASAP7_75t_L g694 ( .A(n_443), .Y(n_694) );
BUFx3_ASAP7_75t_L g831 ( .A(n_443), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_452), .Y(n_444) );
BUFx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_447), .Y(n_618) );
INVx3_ASAP7_75t_L g739 ( .A(n_447), .Y(n_739) );
BUFx3_ASAP7_75t_L g763 ( .A(n_447), .Y(n_763) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_SL g488 ( .A(n_448), .Y(n_488) );
INVx2_ASAP7_75t_L g529 ( .A(n_448), .Y(n_529) );
BUFx2_ASAP7_75t_SL g597 ( .A(n_448), .Y(n_597) );
INVx1_ASAP7_75t_L g879 ( .A(n_449), .Y(n_879) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx3_ASAP7_75t_L g498 ( .A(n_451), .Y(n_498) );
BUFx3_ASAP7_75t_L g530 ( .A(n_451), .Y(n_530) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_451), .Y(n_561) );
INVx2_ASAP7_75t_L g620 ( .A(n_451), .Y(n_620) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g491 ( .A(n_455), .Y(n_491) );
INVx3_ASAP7_75t_L g564 ( .A(n_455), .Y(n_564) );
INVx5_ASAP7_75t_L g600 ( .A(n_455), .Y(n_600) );
INVx4_ASAP7_75t_L g657 ( .A(n_455), .Y(n_657) );
INVx8_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g601 ( .A(n_458), .Y(n_601) );
BUFx2_ASAP7_75t_L g802 ( .A(n_458), .Y(n_802) );
BUFx2_ASAP7_75t_L g876 ( .A(n_458), .Y(n_876) );
INVx6_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g565 ( .A(n_459), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_459), .A2(n_622), .B1(n_623), .B2(n_625), .Y(n_621) );
INVx1_ASAP7_75t_SL g744 ( .A(n_459), .Y(n_744) );
INVx1_ASAP7_75t_L g517 ( .A(n_460), .Y(n_517) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AO22x1_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B1(n_501), .B2(n_532), .Y(n_464) );
INVx2_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
XOR2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_500), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_485), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_474), .C(n_481), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B1(n_472), .B2(n_473), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_471), .A2(n_583), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
OAI221xp5_ASAP7_75t_SL g538 ( .A1(n_473), .A2(n_539), .B1(n_541), .B2(n_542), .C(n_543), .Y(n_538) );
OAI21xp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_478), .Y(n_474) );
OAI21xp5_ASAP7_75t_SL g504 ( .A1(n_476), .A2(n_505), .B(n_506), .Y(n_504) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_479), .Y(n_587) );
BUFx4f_ASAP7_75t_SL g554 ( .A(n_480), .Y(n_554) );
INVx2_ASAP7_75t_L g589 ( .A(n_480), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_492), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_490), .Y(n_486) );
INVx1_ASAP7_75t_L g957 ( .A(n_488), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_497), .Y(n_492) );
INVx1_ASAP7_75t_SL g558 ( .A(n_494), .Y(n_558) );
INVx4_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g660 ( .A(n_495), .Y(n_660) );
INVx2_ASAP7_75t_SL g742 ( .A(n_495), .Y(n_742) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_495), .Y(n_769) );
INVx1_ASAP7_75t_L g936 ( .A(n_495), .Y(n_936) );
INVx1_ASAP7_75t_L g861 ( .A(n_496), .Y(n_861) );
INVx3_ASAP7_75t_SL g532 ( .A(n_501), .Y(n_532) );
AO22x1_ASAP7_75t_L g573 ( .A1(n_501), .A2(n_532), .B1(n_574), .B2(n_609), .Y(n_573) );
XOR2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_531), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_503), .B(n_519), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_507), .Y(n_503) );
NAND3xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_511), .C(n_515), .Y(n_507) );
BUFx4f_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_SL g640 ( .A(n_510), .Y(n_640) );
BUFx2_ASAP7_75t_L g773 ( .A(n_510), .Y(n_773) );
BUFx2_ASAP7_75t_L g791 ( .A(n_510), .Y(n_791) );
BUFx2_ASAP7_75t_L g848 ( .A(n_512), .Y(n_848) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g665 ( .A(n_513), .Y(n_665) );
INVx5_ASAP7_75t_L g709 ( .A(n_513), .Y(n_709) );
INVx2_ASAP7_75t_L g999 ( .A(n_513), .Y(n_999) );
INVx4_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g545 ( .A(n_516), .Y(n_545) );
BUFx2_ASAP7_75t_L g668 ( .A(n_516), .Y(n_668) );
BUFx3_ASAP7_75t_L g711 ( .A(n_516), .Y(n_711) );
BUFx2_ASAP7_75t_L g732 ( .A(n_516), .Y(n_732) );
BUFx6f_ASAP7_75t_L g669 ( .A(n_518), .Y(n_669) );
BUFx2_ASAP7_75t_SL g682 ( .A(n_518), .Y(n_682) );
BUFx3_ASAP7_75t_L g716 ( .A(n_518), .Y(n_716) );
BUFx2_ASAP7_75t_SL g817 ( .A(n_518), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_520), .B(n_524), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_527), .Y(n_524) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx3_ASAP7_75t_L g797 ( .A(n_529), .Y(n_797) );
INVx1_ASAP7_75t_L g612 ( .A(n_533), .Y(n_612) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_572), .B1(n_573), .B2(n_610), .Y(n_534) );
INVx1_ASAP7_75t_SL g610 ( .A(n_535), .Y(n_610) );
INVx1_ASAP7_75t_L g571 ( .A(n_536), .Y(n_571) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_556), .Y(n_536) );
NOR2xp33_ASAP7_75t_SL g537 ( .A(n_538), .B(n_546), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_539), .A2(n_884), .B1(n_885), .B2(n_886), .Y(n_883) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g580 ( .A(n_540), .Y(n_580) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OAI222xp33_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_549), .B1(n_550), .B2(n_552), .C1(n_553), .C2(n_555), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_548), .Y(n_547) );
OAI21xp5_ASAP7_75t_SL g991 ( .A1(n_550), .A2(n_992), .B(n_993), .Y(n_991) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_566), .Y(n_556) );
OAI221xp5_ASAP7_75t_SL g557 ( .A1(n_558), .A2(n_559), .B1(n_560), .B2(n_562), .C(n_563), .Y(n_557) );
OAI221xp5_ASAP7_75t_SL g877 ( .A1(n_558), .A2(n_878), .B1(n_879), .B2(n_880), .C(n_881), .Y(n_877) );
INVx4_ASAP7_75t_L g662 ( .A(n_560), .Y(n_662) );
INVx3_ASAP7_75t_L g748 ( .A(n_560), .Y(n_748) );
OAI221xp5_ASAP7_75t_SL g956 ( .A1(n_560), .A2(n_957), .B1(n_958), .B2(n_959), .C(n_960), .Y(n_956) );
INVx4_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp33_ASAP7_75t_SL g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx2_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g609 ( .A(n_574), .Y(n_609) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_594), .Y(n_576) );
NOR3xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_584), .C(n_590), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_580), .B1(n_581), .B2(n_582), .Y(n_578) );
OA211x2_ASAP7_75t_L g824 ( .A1(n_582), .A2(n_825), .B(n_826), .C(n_827), .Y(n_824) );
OA211x2_ASAP7_75t_L g845 ( .A1(n_582), .A2(n_846), .B(n_847), .C(n_849), .Y(n_845) );
BUFx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g945 ( .A(n_583), .Y(n_945) );
INVx2_ASAP7_75t_SL g888 ( .A(n_587), .Y(n_888) );
INVx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_602), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx2_ASAP7_75t_L g875 ( .A(n_600), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_607), .Y(n_602) );
BUFx4f_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g965 ( .A(n_605), .Y(n_965) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_699), .B1(n_834), .B2(n_835), .Y(n_613) );
INVx2_ASAP7_75t_SL g834 ( .A(n_614), .Y(n_834) );
OA22x2_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_648), .B1(n_649), .B2(n_698), .Y(n_614) );
INVx1_ASAP7_75t_L g698 ( .A(n_615), .Y(n_698) );
INVx1_ASAP7_75t_L g647 ( .A(n_616), .Y(n_647) );
AND4x1_ASAP7_75t_L g616 ( .A(n_617), .B(n_626), .C(n_638), .D(n_644), .Y(n_616) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
BUFx2_ASAP7_75t_R g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_635), .B2(n_636), .Y(n_630) );
OAI221xp5_ASAP7_75t_SL g870 ( .A1(n_632), .A2(n_871), .B1(n_872), .B2(n_873), .C(n_874), .Y(n_870) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g853 ( .A(n_633), .Y(n_853) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_SL g666 ( .A(n_640), .Y(n_666) );
INVx2_ASAP7_75t_SL g723 ( .A(n_645), .Y(n_723) );
INVx2_ASAP7_75t_L g890 ( .A(n_645), .Y(n_890) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_675), .B1(n_696), .B2(n_697), .Y(n_649) );
INVx2_ASAP7_75t_SL g696 ( .A(n_650), .Y(n_696) );
XOR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_674), .Y(n_650) );
NOR4xp75_ASAP7_75t_L g651 ( .A(n_652), .B(n_658), .C(n_663), .D(n_670), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVx1_ASAP7_75t_L g1007 ( .A(n_654), .Y(n_1007) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2x1_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_664), .B(n_667), .Y(n_663) );
INVx1_ASAP7_75t_SL g786 ( .A(n_669), .Y(n_786) );
INVx1_ASAP7_75t_L g697 ( .A(n_675), .Y(n_697) );
OA22x2_ASAP7_75t_SL g718 ( .A1(n_675), .A2(n_697), .B1(n_719), .B2(n_750), .Y(n_718) );
XOR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_695), .Y(n_675) );
NAND2x1_ASAP7_75t_L g676 ( .A(n_677), .B(n_687), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_683), .Y(n_677) );
OAI21xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_680), .B(n_681), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .C(n_686), .Y(n_683) );
NOR2x1_ASAP7_75t_L g687 ( .A(n_688), .B(n_691), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_L g835 ( .A(n_699), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_753), .B2(n_754), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_718), .B1(n_751), .B2(n_752), .Y(n_701) );
INVx2_ASAP7_75t_SL g751 ( .A(n_702), .Y(n_751) );
XOR2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_717), .Y(n_702) );
NAND4xp75_ASAP7_75t_L g703 ( .A(n_704), .B(n_707), .C(n_712), .D(n_715), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
AND2x2_ASAP7_75t_SL g707 ( .A(n_708), .B(n_710), .Y(n_707) );
BUFx6f_ASAP7_75t_L g734 ( .A(n_709), .Y(n_734) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_709), .Y(n_789) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx2_ASAP7_75t_L g752 ( .A(n_718), .Y(n_752) );
INVx1_ASAP7_75t_L g750 ( .A(n_719), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_735), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_730), .Y(n_721) );
OAI222xp33_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B1(n_725), .B2(n_727), .C1(n_728), .C2(n_729), .Y(n_722) );
OAI21xp5_ASAP7_75t_SL g912 ( .A1(n_723), .A2(n_913), .B(n_914), .Y(n_912) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx4_ASAP7_75t_L g995 ( .A(n_726), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_745), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_737), .B(n_743), .Y(n_736) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
OAI22x1_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B1(n_818), .B2(n_819), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
XNOR2x1_ASAP7_75t_L g756 ( .A(n_757), .B(n_777), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
NAND4xp75_ASAP7_75t_SL g760 ( .A(n_761), .B(n_766), .C(n_771), .D(n_775), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_764), .Y(n_761) );
INVxp67_ASAP7_75t_L g854 ( .A(n_765), .Y(n_854) );
AND2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_770), .Y(n_766) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
AND2x2_ASAP7_75t_SL g771 ( .A(n_772), .B(n_774), .Y(n_771) );
XOR2x2_ASAP7_75t_L g777 ( .A(n_778), .B(n_803), .Y(n_777) );
NAND2xp5_ASAP7_75t_SL g779 ( .A(n_780), .B(n_793), .Y(n_779) );
NOR2xp33_ASAP7_75t_SL g780 ( .A(n_781), .B(n_787), .Y(n_780) );
OAI21xp5_ASAP7_75t_SL g781 ( .A1(n_782), .A2(n_783), .B(n_784), .Y(n_781) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NAND3xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_790), .C(n_792), .Y(n_787) );
NOR2x1_ASAP7_75t_L g793 ( .A(n_794), .B(n_798), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_801), .Y(n_798) );
NAND4xp75_ASAP7_75t_L g804 ( .A(n_805), .B(n_808), .C(n_813), .D(n_816), .Y(n_804) );
AND2x2_ASAP7_75t_SL g805 ( .A(n_806), .B(n_807), .Y(n_805) );
AND2x2_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
AND2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
INVx3_ASAP7_75t_SL g818 ( .A(n_819), .Y(n_818) );
XOR2x2_ASAP7_75t_L g819 ( .A(n_820), .B(n_833), .Y(n_819) );
NAND4xp75_ASAP7_75t_L g820 ( .A(n_821), .B(n_824), .C(n_828), .D(n_832), .Y(n_820) );
AND2x2_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
AND2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
INVx1_ASAP7_75t_L g972 ( .A(n_836), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_838), .B1(n_904), .B2(n_970), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_839), .A2(n_865), .B1(n_866), .B2(n_903), .Y(n_838) );
INVx1_ASAP7_75t_SL g903 ( .A(n_839), .Y(n_903) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
XOR2x2_ASAP7_75t_L g840 ( .A(n_841), .B(n_864), .Y(n_840) );
NAND4xp75_ASAP7_75t_L g841 ( .A(n_842), .B(n_845), .C(n_850), .D(n_862), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_856), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_852), .A2(n_853), .B1(n_854), .B2(n_855), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_858), .B1(n_860), .B2(n_861), .Y(n_856) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g902 ( .A(n_868), .Y(n_902) );
AND2x2_ASAP7_75t_L g868 ( .A(n_869), .B(n_882), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_870), .B(n_877), .Y(n_869) );
NOR3xp33_ASAP7_75t_L g882 ( .A(n_883), .B(n_887), .C(n_895), .Y(n_882) );
OAI222xp33_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .B1(n_890), .B2(n_891), .C1(n_892), .C2(n_894), .Y(n_887) );
OAI222xp33_ASAP7_75t_L g946 ( .A1(n_890), .A2(n_947), .B1(n_948), .B2(n_949), .C1(n_950), .C2(n_951), .Y(n_946) );
INVx2_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_896), .A2(n_897), .B1(n_898), .B2(n_899), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_897), .A2(n_899), .B1(n_953), .B2(n_954), .Y(n_952) );
INVx2_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g970 ( .A(n_904), .Y(n_970) );
INVx2_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_SL g905 ( .A(n_906), .Y(n_905) );
AOI22xp5_ASAP7_75t_L g906 ( .A1(n_907), .A2(n_908), .B1(n_938), .B2(n_969), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
XNOR2xp5_ASAP7_75t_L g908 ( .A(n_909), .B(n_925), .Y(n_908) );
NAND3xp33_ASAP7_75t_L g910 ( .A(n_911), .B(n_919), .C(n_922), .Y(n_910) );
NOR2xp33_ASAP7_75t_L g911 ( .A(n_912), .B(n_915), .Y(n_911) );
NAND3xp33_ASAP7_75t_L g915 ( .A(n_916), .B(n_917), .C(n_918), .Y(n_915) );
AND2x2_ASAP7_75t_L g919 ( .A(n_920), .B(n_921), .Y(n_919) );
AND2x2_ASAP7_75t_L g922 ( .A(n_923), .B(n_924), .Y(n_922) );
NAND4xp75_ASAP7_75t_L g926 ( .A(n_927), .B(n_930), .C(n_933), .D(n_937), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .Y(n_927) );
AND2x2_ASAP7_75t_SL g930 ( .A(n_931), .B(n_932), .Y(n_930) );
AND2x2_ASAP7_75t_L g933 ( .A(n_934), .B(n_935), .Y(n_933) );
INVx1_ASAP7_75t_L g969 ( .A(n_938), .Y(n_969) );
INVx1_ASAP7_75t_L g968 ( .A(n_939), .Y(n_968) );
AND2x2_ASAP7_75t_L g939 ( .A(n_940), .B(n_955), .Y(n_939) );
NOR3xp33_ASAP7_75t_L g940 ( .A(n_941), .B(n_946), .C(n_952), .Y(n_940) );
INVx2_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
NOR2xp33_ASAP7_75t_L g955 ( .A(n_956), .B(n_961), .Y(n_955) );
NAND2xp5_ASAP7_75t_SL g961 ( .A(n_962), .B(n_963), .Y(n_961) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx2_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
NOR2x1_ASAP7_75t_L g974 ( .A(n_975), .B(n_979), .Y(n_974) );
OR2x2_ASAP7_75t_SL g1044 ( .A(n_975), .B(n_980), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_976), .B(n_978), .Y(n_975) );
CKINVDCx20_ASAP7_75t_R g1013 ( .A(n_976), .Y(n_1013) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_977), .B(n_1017), .Y(n_1020) );
CKINVDCx16_ASAP7_75t_R g1017 ( .A(n_978), .Y(n_1017) );
CKINVDCx20_ASAP7_75t_R g979 ( .A(n_980), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_981), .B(n_982), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_984), .B(n_985), .Y(n_983) );
OAI322xp33_ASAP7_75t_L g986 ( .A1(n_987), .A2(n_1011), .A3(n_1014), .B1(n_1018), .B2(n_1021), .C1(n_1022), .C2(n_1042), .Y(n_986) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
NAND3x2_ASAP7_75t_L g989 ( .A(n_990), .B(n_1001), .C(n_1004), .Y(n_989) );
NOR2x1_ASAP7_75t_SL g990 ( .A(n_991), .B(n_996), .Y(n_990) );
INVx3_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
NAND3xp33_ASAP7_75t_L g996 ( .A(n_997), .B(n_998), .C(n_1000), .Y(n_996) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1003), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1008), .Y(n_1004) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
HB1xp67_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
BUFx2_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
HB1xp67_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
CKINVDCx16_ASAP7_75t_R g1018 ( .A(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
AND3x1_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1035), .C(n_1038), .Y(n_1024) );
NOR3xp33_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1029), .C(n_1032), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1031), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1037), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1040), .Y(n_1038) );
CKINVDCx20_ASAP7_75t_R g1042 ( .A(n_1043), .Y(n_1042) );
CKINVDCx20_ASAP7_75t_R g1043 ( .A(n_1044), .Y(n_1043) );
endmodule