module fake_jpeg_25323_n_230 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_33),
.B(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_17),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_20),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_19),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_24),
.B1(n_15),
.B2(n_27),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_41),
.B1(n_40),
.B2(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_49),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_24),
.B1(n_28),
.B2(n_27),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_54),
.B1(n_41),
.B2(n_39),
.Y(n_68)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_55),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_24),
.B1(n_25),
.B2(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_23),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_25),
.B(n_19),
.C(n_20),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_38),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_24),
.B1(n_40),
.B2(n_41),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_64),
.A2(n_67),
.B1(n_70),
.B2(n_75),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_48),
.B1(n_18),
.B2(n_27),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_73),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_31),
.B1(n_30),
.B2(n_36),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_18),
.B1(n_28),
.B2(n_26),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_71),
.Y(n_82)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_60),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_18),
.B1(n_28),
.B2(n_26),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_33),
.Y(n_76)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_1),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_26),
.B1(n_29),
.B2(n_22),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_77),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_52),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_21),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_59),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_86),
.B(n_72),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_51),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_52),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_47),
.B(n_29),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_100),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_74),
.B(n_21),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_93),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_94),
.A2(n_101),
.B1(n_73),
.B2(n_63),
.Y(n_102)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_71),
.B1(n_66),
.B2(n_46),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_58),
.Y(n_100)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_102),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_65),
.B1(n_64),
.B2(n_80),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_108),
.B1(n_89),
.B2(n_85),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_114),
.B(n_119),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_72),
.B1(n_42),
.B2(n_69),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_111),
.B1(n_121),
.B2(n_89),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_106),
.B(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_107),
.B(n_21),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_77),
.B1(n_66),
.B2(n_42),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_100),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_69),
.B1(n_62),
.B2(n_73),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_81),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_62),
.C(n_56),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_89),
.C(n_95),
.Y(n_123)
);

NOR2xp67_ASAP7_75t_SL g114 ( 
.A(n_84),
.B(n_36),
.Y(n_114)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_101),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_29),
.B1(n_22),
.B2(n_16),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_83),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_134),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_129),
.C(n_119),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_97),
.B(n_86),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_133),
.B(n_105),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_128),
.B1(n_131),
.B2(n_108),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_93),
.C(n_90),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_85),
.B1(n_88),
.B2(n_82),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_82),
.B(n_91),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_90),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_120),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_137),
.B(n_138),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_94),
.B(n_2),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_94),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_139),
.B(n_141),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_142),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_1),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_148),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_146),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_147),
.A2(n_142),
.B(n_107),
.Y(n_169)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_153),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_157),
.Y(n_165)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_159),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_161),
.Y(n_167)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_130),
.C(n_133),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_109),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_160),
.B(n_118),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_129),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_128),
.B1(n_132),
.B2(n_127),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_164),
.B1(n_168),
.B2(n_16),
.Y(n_188)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_150),
.A2(n_152),
.B1(n_157),
.B2(n_141),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_170),
.C(n_174),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_155),
.A2(n_136),
.B1(n_111),
.B2(n_130),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_162),
.B(n_165),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_122),
.C(n_121),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_47),
.C(n_22),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_155),
.B(n_14),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_160),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_180),
.Y(n_195)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_171),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_183),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_173),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_176),
.A2(n_149),
.B1(n_147),
.B2(n_144),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

AOI322xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_156),
.A3(n_145),
.B1(n_159),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_191),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_187),
.B(n_9),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_188),
.A2(n_190),
.B1(n_4),
.B2(n_5),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_167),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_199),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_167),
.C(n_174),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_198),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_5),
.B(n_8),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_202),
.B(n_184),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_197),
.A2(n_189),
.B1(n_187),
.B2(n_179),
.Y(n_204)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_10),
.Y(n_215)
);

INVx11_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_210),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_209),
.B(n_13),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_195),
.A2(n_194),
.B1(n_181),
.B2(n_198),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_196),
.B(n_192),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_214),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_210),
.A2(n_201),
.B(n_193),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_217),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_216),
.B(n_205),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_11),
.Y(n_217)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

NAND2xp33_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_204),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_222),
.B(n_216),
.C(n_207),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_208),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_12),
.C(n_223),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_220),
.A2(n_206),
.B(n_11),
.Y(n_225)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_225),
.B(n_218),
.CI(n_12),
.CON(n_226),
.SN(n_226)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_227),
.B(n_12),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_226),
.B(n_227),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_226),
.Y(n_230)
);


endmodule