module fake_netlist_1_10659_n_802 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_92, n_11, n_223, n_25, n_30, n_59, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_96, n_39, n_802);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_96;
input n_39;
output n_802;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_580;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_230;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_565;
wire n_224;
wire n_788;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_774;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g224 ( .A(n_79), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_89), .Y(n_225) );
INVx1_ASAP7_75t_SL g226 ( .A(n_193), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_98), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_156), .Y(n_228) );
INVx1_ASAP7_75t_SL g229 ( .A(n_101), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_37), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_167), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_155), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_40), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_151), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_219), .Y(n_235) );
NOR2xp67_ASAP7_75t_L g236 ( .A(n_5), .B(n_78), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_138), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_108), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_77), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_73), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_129), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_187), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_36), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_123), .Y(n_244) );
CKINVDCx14_ASAP7_75t_R g245 ( .A(n_64), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_38), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_91), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_179), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_60), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_199), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_51), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_109), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_92), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_131), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_130), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_119), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_136), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_139), .Y(n_258) );
BUFx2_ASAP7_75t_L g259 ( .A(n_70), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_102), .Y(n_260) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_110), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_57), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_46), .B(n_124), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_173), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_195), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_125), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_200), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_87), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_180), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_24), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_134), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_29), .Y(n_272) );
CKINVDCx16_ASAP7_75t_R g273 ( .A(n_39), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_161), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_223), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_3), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_117), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_217), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_22), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_215), .B(n_182), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_164), .Y(n_281) );
CKINVDCx16_ASAP7_75t_R g282 ( .A(n_159), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_75), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_47), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_145), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_211), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_18), .Y(n_287) );
BUFx2_ASAP7_75t_L g288 ( .A(n_146), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_53), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_137), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_48), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_220), .Y(n_292) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_175), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_68), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_186), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_196), .Y(n_296) );
NOR2xp67_ASAP7_75t_L g297 ( .A(n_86), .B(n_35), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_132), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_170), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_172), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_162), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_113), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_184), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_114), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_191), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_212), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_222), .Y(n_307) );
BUFx10_ASAP7_75t_L g308 ( .A(n_177), .Y(n_308) );
CKINVDCx14_ASAP7_75t_R g309 ( .A(n_154), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_153), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_190), .Y(n_311) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_208), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_1), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_127), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_8), .Y(n_315) );
BUFx5_ASAP7_75t_L g316 ( .A(n_62), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_183), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_202), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_116), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_66), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_96), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_142), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_7), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_197), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_45), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_112), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_56), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_140), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_178), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_99), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_76), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_23), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_88), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_80), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_69), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_19), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_160), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g338 ( .A(n_16), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_194), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_152), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_165), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_188), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_248), .Y(n_343) );
INVx4_ASAP7_75t_L g344 ( .A(n_259), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_232), .B(n_0), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_232), .B(n_0), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_256), .B(n_1), .Y(n_347) );
OA21x2_ASAP7_75t_L g348 ( .A1(n_225), .A2(n_26), .B(n_25), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_256), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_278), .B(n_2), .Y(n_350) );
BUFx12f_ASAP7_75t_L g351 ( .A(n_308), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_288), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_327), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_327), .Y(n_354) );
BUFx12f_ASAP7_75t_L g355 ( .A(n_308), .Y(n_355) );
CKINVDCx6p67_ASAP7_75t_R g356 ( .A(n_273), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_334), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_327), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_282), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_276), .B(n_4), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_279), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_245), .B(n_6), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_313), .B(n_8), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_316), .Y(n_364) );
INVx2_ASAP7_75t_SL g365 ( .A(n_287), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_327), .Y(n_366) );
BUFx12f_ASAP7_75t_L g367 ( .A(n_227), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_224), .B(n_9), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_364), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_364), .B(n_316), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_343), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_353), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_353), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_349), .B(n_309), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_360), .B(n_316), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_360), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_343), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_360), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_362), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_363), .Y(n_380) );
INVx3_ASAP7_75t_L g381 ( .A(n_363), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_344), .B(n_309), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_346), .Y(n_383) );
AND3x2_ASAP7_75t_L g384 ( .A(n_346), .B(n_347), .C(n_352), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_346), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_365), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_347), .B(n_316), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_361), .B(n_316), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_359), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_356), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_353), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_353), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_354), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_357), .B(n_323), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_371), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_374), .B(n_345), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_382), .B(n_350), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_369), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_381), .B(n_351), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_383), .B(n_228), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_369), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_372), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_381), .B(n_359), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_377), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_385), .A2(n_315), .B1(n_368), .B2(n_238), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_379), .B(n_355), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_384), .B(n_355), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_386), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_384), .B(n_367), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_394), .A2(n_367), .B1(n_237), .B2(n_293), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_380), .B(n_230), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_376), .B(n_261), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_389), .Y(n_413) );
NOR3xp33_ASAP7_75t_L g414 ( .A(n_390), .B(n_336), .C(n_240), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_378), .B(n_231), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_387), .B(n_233), .Y(n_416) );
INVxp67_ASAP7_75t_L g417 ( .A(n_387), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_375), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_372), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_373), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_375), .B(n_226), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_388), .B(n_234), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_388), .B(n_246), .Y(n_423) );
O2A1O1Ixp33_ASAP7_75t_L g424 ( .A1(n_370), .A2(n_241), .B(n_242), .C(n_235), .Y(n_424) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_370), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_373), .B(n_247), .Y(n_426) );
NOR3xp33_ASAP7_75t_L g427 ( .A(n_391), .B(n_244), .C(n_243), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_391), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_392), .B(n_251), .Y(n_429) );
OAI21xp33_ASAP7_75t_L g430 ( .A1(n_396), .A2(n_338), .B(n_229), .Y(n_430) );
O2A1O1Ixp33_ASAP7_75t_SL g431 ( .A1(n_400), .A2(n_280), .B(n_263), .C(n_252), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_397), .B(n_300), .Y(n_432) );
AND2x4_ASAP7_75t_L g433 ( .A(n_407), .B(n_310), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_418), .B(n_253), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_405), .B(n_312), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_400), .A2(n_348), .B(n_257), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_415), .A2(n_348), .B(n_264), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g438 ( .A1(n_417), .A2(n_265), .B(n_254), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_399), .B(n_330), .Y(n_439) );
BUFx3_ASAP7_75t_L g440 ( .A(n_413), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_413), .Y(n_441) );
OAI21xp5_ASAP7_75t_L g442 ( .A1(n_398), .A2(n_270), .B(n_269), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_399), .B(n_229), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_421), .B(n_255), .Y(n_444) );
INVx4_ASAP7_75t_L g445 ( .A(n_412), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_421), .B(n_258), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_401), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_408), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_411), .A2(n_275), .B(n_274), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_416), .A2(n_283), .B(n_281), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_409), .B(n_236), .Y(n_451) );
NAND2xp33_ASAP7_75t_L g452 ( .A(n_425), .B(n_316), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_401), .A2(n_286), .B(n_284), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_403), .B(n_260), .Y(n_454) );
OAI21xp33_ASAP7_75t_SL g455 ( .A1(n_395), .A2(n_295), .B(n_290), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_422), .A2(n_306), .B(n_305), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_406), .B(n_266), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_423), .A2(n_317), .B(n_311), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_404), .B(n_267), .Y(n_459) );
BUFx2_ASAP7_75t_L g460 ( .A(n_412), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_404), .B(n_268), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_426), .A2(n_319), .B(n_318), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_410), .Y(n_463) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_425), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_425), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_425), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_437), .A2(n_429), .B(n_424), .Y(n_467) );
INVx2_ASAP7_75t_SL g468 ( .A(n_440), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_447), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_436), .A2(n_419), .B(n_402), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_441), .B(n_414), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_465), .A2(n_420), .B(n_428), .Y(n_472) );
OAI21x1_ASAP7_75t_L g473 ( .A1(n_466), .A2(n_420), .B(n_324), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_432), .B(n_427), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g475 ( .A1(n_456), .A2(n_325), .B(n_322), .Y(n_475) );
OR2x6_ASAP7_75t_L g476 ( .A(n_445), .B(n_297), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_444), .A2(n_328), .B(n_326), .Y(n_477) );
OAI21x1_ASAP7_75t_L g478 ( .A1(n_453), .A2(n_337), .B(n_331), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_446), .A2(n_342), .B(n_271), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_442), .A2(n_272), .B(n_239), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_447), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_439), .B(n_285), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_431), .A2(n_294), .B(n_289), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_458), .A2(n_329), .B(n_302), .Y(n_484) );
BUFx8_ASAP7_75t_SL g485 ( .A(n_460), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_450), .A2(n_339), .B(n_332), .Y(n_486) );
OAI21x1_ASAP7_75t_L g487 ( .A1(n_462), .A2(n_341), .B(n_392), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_430), .B(n_291), .Y(n_488) );
AO31x2_ASAP7_75t_L g489 ( .A1(n_449), .A2(n_438), .A3(n_443), .B(n_448), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_454), .B(n_451), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_455), .A2(n_249), .B(n_277), .C(n_320), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_447), .Y(n_492) );
NAND2x1p5_ASAP7_75t_L g493 ( .A(n_433), .B(n_250), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_435), .B(n_292), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_452), .A2(n_393), .B(n_298), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_459), .A2(n_299), .B(n_296), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_463), .A2(n_451), .B1(n_457), .B2(n_434), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_461), .Y(n_498) );
OAI21x1_ASAP7_75t_L g499 ( .A1(n_464), .A2(n_262), .B(n_250), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_464), .A2(n_303), .B(n_301), .Y(n_500) );
INVx2_ASAP7_75t_SL g501 ( .A(n_464), .Y(n_501) );
OAI21x1_ASAP7_75t_L g502 ( .A1(n_437), .A2(n_262), .B(n_250), .Y(n_502) );
AOI21x1_ASAP7_75t_L g503 ( .A1(n_437), .A2(n_262), .B(n_354), .Y(n_503) );
OAI21x1_ASAP7_75t_L g504 ( .A1(n_437), .A2(n_28), .B(n_27), .Y(n_504) );
OAI21x1_ASAP7_75t_L g505 ( .A1(n_502), .A2(n_358), .B(n_354), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_468), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_493), .Y(n_507) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_503), .A2(n_307), .B(n_304), .Y(n_508) );
INVxp67_ASAP7_75t_SL g509 ( .A(n_469), .Y(n_509) );
NOR2xp67_ASAP7_75t_L g510 ( .A(n_471), .B(n_10), .Y(n_510) );
BUFx2_ASAP7_75t_R g511 ( .A(n_485), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_498), .Y(n_512) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_467), .A2(n_366), .B(n_358), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_474), .B(n_11), .Y(n_514) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_504), .A2(n_366), .B(n_358), .Y(n_515) );
BUFx3_ASAP7_75t_L g516 ( .A(n_490), .Y(n_516) );
INVx3_ASAP7_75t_L g517 ( .A(n_469), .Y(n_517) );
OAI21x1_ASAP7_75t_L g518 ( .A1(n_499), .A2(n_366), .B(n_31), .Y(n_518) );
AO31x2_ASAP7_75t_L g519 ( .A1(n_470), .A2(n_366), .A3(n_12), .B(n_13), .Y(n_519) );
INVx2_ASAP7_75t_SL g520 ( .A(n_476), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_469), .Y(n_521) );
NOR2xp33_ASAP7_75t_SL g522 ( .A(n_480), .B(n_314), .Y(n_522) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_481), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_478), .Y(n_524) );
OAI21x1_ASAP7_75t_L g525 ( .A1(n_473), .A2(n_32), .B(n_30), .Y(n_525) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_487), .A2(n_333), .B(n_321), .Y(n_526) );
OR2x6_ASAP7_75t_L g527 ( .A(n_476), .B(n_11), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_489), .B(n_12), .Y(n_528) );
OAI21x1_ASAP7_75t_L g529 ( .A1(n_472), .A2(n_34), .B(n_33), .Y(n_529) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_483), .A2(n_340), .B(n_335), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_489), .Y(n_531) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_480), .A2(n_118), .B(n_218), .Y(n_532) );
NAND2x1p5_ASAP7_75t_L g533 ( .A(n_501), .B(n_13), .Y(n_533) );
OAI21x1_ASAP7_75t_L g534 ( .A1(n_492), .A2(n_120), .B(n_216), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_497), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_535) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_491), .A2(n_121), .B(n_214), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_484), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_494), .Y(n_538) );
OAI21x1_ASAP7_75t_L g539 ( .A1(n_486), .A2(n_115), .B(n_213), .Y(n_539) );
INVx3_ASAP7_75t_L g540 ( .A(n_482), .Y(n_540) );
BUFx3_ASAP7_75t_L g541 ( .A(n_488), .Y(n_541) );
OAI21x1_ASAP7_75t_L g542 ( .A1(n_479), .A2(n_111), .B(n_210), .Y(n_542) );
OAI21x1_ASAP7_75t_L g543 ( .A1(n_495), .A2(n_107), .B(n_209), .Y(n_543) );
BUFx2_ASAP7_75t_SL g544 ( .A(n_500), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_475), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_477), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_496), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_485), .Y(n_548) );
OAI21x1_ASAP7_75t_L g549 ( .A1(n_502), .A2(n_106), .B(n_207), .Y(n_549) );
AOI21x1_ASAP7_75t_L g550 ( .A1(n_503), .A2(n_105), .B(n_206), .Y(n_550) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_469), .Y(n_551) );
OAI21x1_ASAP7_75t_L g552 ( .A1(n_502), .A2(n_104), .B(n_205), .Y(n_552) );
OAI21x1_ASAP7_75t_L g553 ( .A1(n_502), .A2(n_103), .B(n_204), .Y(n_553) );
AOI21x1_ASAP7_75t_L g554 ( .A1(n_503), .A2(n_100), .B(n_203), .Y(n_554) );
OR2x6_ASAP7_75t_L g555 ( .A(n_468), .B(n_17), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_485), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_533), .Y(n_557) );
OAI21x1_ASAP7_75t_L g558 ( .A1(n_505), .A2(n_122), .B(n_201), .Y(n_558) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_545), .A2(n_20), .B(n_21), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_531), .Y(n_560) );
OAI221xp5_ASAP7_75t_L g561 ( .A1(n_535), .A2(n_22), .B1(n_41), .B2(n_42), .C(n_43), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_519), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_519), .Y(n_563) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_551), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_533), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_555), .B(n_44), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_535), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_513), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_513), .Y(n_569) );
AO21x1_ASAP7_75t_SL g570 ( .A1(n_507), .A2(n_49), .B(n_50), .Y(n_570) );
CKINVDCx11_ASAP7_75t_R g571 ( .A(n_512), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_519), .Y(n_572) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_521), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_514), .Y(n_574) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_551), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_528), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_506), .B(n_52), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_524), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_514), .Y(n_579) );
AO21x2_ASAP7_75t_L g580 ( .A1(n_515), .A2(n_54), .B(n_55), .Y(n_580) );
INVx2_ASAP7_75t_SL g581 ( .A(n_548), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_510), .Y(n_582) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_521), .Y(n_583) );
CKINVDCx11_ASAP7_75t_R g584 ( .A(n_527), .Y(n_584) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_511), .Y(n_585) );
OAI21x1_ASAP7_75t_L g586 ( .A1(n_549), .A2(n_58), .B(n_59), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_522), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_522), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_546), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_517), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_517), .Y(n_591) );
INVx3_ASAP7_75t_L g592 ( .A(n_540), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_537), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_509), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_516), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_547), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_523), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_538), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_541), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_520), .A2(n_61), .B1(n_63), .B2(n_65), .C(n_67), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_526), .Y(n_601) );
BUFx3_ASAP7_75t_L g602 ( .A(n_556), .Y(n_602) );
INVx2_ASAP7_75t_SL g603 ( .A(n_511), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_542), .Y(n_604) );
CKINVDCx11_ASAP7_75t_R g605 ( .A(n_544), .Y(n_605) );
BUFx2_ASAP7_75t_L g606 ( .A(n_509), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_530), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_525), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_539), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_536), .Y(n_610) );
OA21x2_ASAP7_75t_L g611 ( .A1(n_552), .A2(n_71), .B(n_72), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_529), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_534), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_543), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_532), .Y(n_615) );
NAND2x1p5_ASAP7_75t_L g616 ( .A(n_553), .B(n_74), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_550), .Y(n_617) );
INVx3_ASAP7_75t_L g618 ( .A(n_518), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_554), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_508), .Y(n_620) );
OAI21x1_ASAP7_75t_L g621 ( .A1(n_508), .A2(n_81), .B(n_82), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_515), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_545), .A2(n_221), .B1(n_84), .B2(n_85), .Y(n_623) );
BUFx5_ASAP7_75t_L g624 ( .A(n_557), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_574), .B(n_83), .Y(n_625) );
INVxp67_ASAP7_75t_L g626 ( .A(n_594), .Y(n_626) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_559), .A2(n_90), .B1(n_93), .B2(n_94), .Y(n_627) );
BUFx2_ASAP7_75t_L g628 ( .A(n_606), .Y(n_628) );
AND2x4_ASAP7_75t_L g629 ( .A(n_594), .B(n_95), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_597), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_598), .B(n_97), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_579), .B(n_126), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_589), .Y(n_633) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_560), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_599), .B(n_128), .Y(n_635) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_560), .Y(n_636) );
AND2x4_ASAP7_75t_SL g637 ( .A(n_566), .B(n_133), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_567), .B(n_135), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_593), .Y(n_639) );
INVx3_ASAP7_75t_L g640 ( .A(n_564), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_576), .B(n_141), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_584), .A2(n_143), .B1(n_144), .B2(n_147), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_587), .A2(n_148), .B1(n_149), .B2(n_150), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_592), .Y(n_644) );
INVx4_ASAP7_75t_L g645 ( .A(n_605), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_573), .B(n_157), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_583), .B(n_158), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_596), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_571), .Y(n_649) );
INVx2_ASAP7_75t_SL g650 ( .A(n_602), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_595), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_565), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_578), .Y(n_653) );
BUFx4f_ASAP7_75t_L g654 ( .A(n_603), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_583), .Y(n_655) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_568), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_582), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_559), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_590), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_591), .Y(n_660) );
INVx2_ASAP7_75t_SL g661 ( .A(n_581), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_561), .A2(n_163), .B1(n_166), .B2(n_168), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_577), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_607), .B(n_169), .Y(n_664) );
OAI21xp5_ASAP7_75t_SL g665 ( .A1(n_587), .A2(n_171), .B(n_174), .Y(n_665) );
OR2x2_ASAP7_75t_L g666 ( .A(n_588), .B(n_176), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_564), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_564), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_575), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_585), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_570), .B(n_181), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_562), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_601), .B(n_185), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_563), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_572), .Y(n_675) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_623), .A2(n_189), .B1(n_192), .B2(n_198), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_620), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_569), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_610), .B(n_614), .Y(n_679) );
AO31x2_ASAP7_75t_L g680 ( .A1(n_608), .A2(n_604), .A3(n_619), .B(n_617), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_600), .B(n_621), .Y(n_681) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_622), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_616), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_616), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_586), .Y(n_685) );
BUFx4f_ASAP7_75t_SL g686 ( .A(n_618), .Y(n_686) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_634), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_628), .B(n_609), .Y(n_688) );
BUFx2_ASAP7_75t_L g689 ( .A(n_645), .Y(n_689) );
INVx2_ASAP7_75t_SL g690 ( .A(n_645), .Y(n_690) );
INVx5_ASAP7_75t_L g691 ( .A(n_629), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_651), .B(n_612), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_657), .B(n_613), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_652), .B(n_580), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_665), .A2(n_611), .B1(n_615), .B2(n_618), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_678), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_663), .B(n_558), .Y(n_697) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_634), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_655), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_677), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_653), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_626), .B(n_659), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_660), .B(n_636), .Y(n_703) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_636), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_633), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_639), .Y(n_706) );
BUFx2_ASAP7_75t_SL g707 ( .A(n_649), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_650), .B(n_630), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_648), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_658), .B(n_644), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_646), .B(n_647), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_672), .Y(n_712) );
OR2x2_ASAP7_75t_L g713 ( .A(n_661), .B(n_656), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_674), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_675), .Y(n_715) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_682), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_679), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_624), .Y(n_718) );
INVx3_ASAP7_75t_L g719 ( .A(n_686), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_631), .B(n_668), .Y(n_720) );
AND2x4_ASAP7_75t_L g721 ( .A(n_684), .B(n_683), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_667), .B(n_669), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_624), .Y(n_723) );
AOI22xp33_ASAP7_75t_SL g724 ( .A1(n_681), .A2(n_654), .B1(n_624), .B2(n_637), .Y(n_724) );
BUFx3_ASAP7_75t_L g725 ( .A(n_640), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_654), .A2(n_662), .B1(n_676), .B2(n_627), .Y(n_726) );
AND2x4_ASAP7_75t_L g727 ( .A(n_680), .B(n_640), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_680), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g729 ( .A(n_624), .B(n_686), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_635), .B(n_638), .Y(n_730) );
INVx2_ASAP7_75t_SL g731 ( .A(n_671), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_664), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_664), .Y(n_733) );
OR2x2_ASAP7_75t_L g734 ( .A(n_713), .B(n_666), .Y(n_734) );
OR2x2_ASAP7_75t_L g735 ( .A(n_687), .B(n_673), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_692), .B(n_685), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_693), .B(n_694), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_699), .B(n_625), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_705), .B(n_632), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_698), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_706), .B(n_632), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_708), .B(n_641), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_702), .B(n_641), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_700), .B(n_662), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_704), .Y(n_745) );
INVx1_ASAP7_75t_SL g746 ( .A(n_707), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_688), .B(n_643), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_717), .B(n_643), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_703), .B(n_642), .Y(n_749) );
BUFx2_ASAP7_75t_L g750 ( .A(n_689), .Y(n_750) );
OR2x2_ASAP7_75t_L g751 ( .A(n_716), .B(n_670), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_709), .Y(n_752) );
AND2x4_ASAP7_75t_L g753 ( .A(n_727), .B(n_691), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_696), .B(n_712), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_701), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_712), .B(n_714), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_714), .B(n_715), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_732), .B(n_733), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_737), .B(n_710), .Y(n_759) );
OAI22xp33_ASAP7_75t_SL g760 ( .A1(n_750), .A2(n_751), .B1(n_731), .B2(n_746), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_736), .B(n_697), .Y(n_761) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_757), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_736), .B(n_727), .Y(n_763) );
INVx2_ASAP7_75t_SL g764 ( .A(n_756), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_742), .B(n_731), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_756), .B(n_727), .Y(n_766) );
INVxp67_ASAP7_75t_SL g767 ( .A(n_755), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_754), .B(n_728), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_753), .B(n_728), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_752), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_740), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g772 ( .A(n_760), .B(n_691), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_762), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_762), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_761), .B(n_745), .Y(n_775) );
INVx1_ASAP7_75t_SL g776 ( .A(n_765), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_766), .B(n_753), .Y(n_777) );
AOI322xp5_ASAP7_75t_L g778 ( .A1(n_763), .A2(n_690), .A3(n_726), .B1(n_747), .B2(n_748), .C1(n_724), .C2(n_749), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_759), .B(n_748), .Y(n_779) );
A2O1A1Ixp33_ASAP7_75t_L g780 ( .A1(n_778), .A2(n_719), .B(n_763), .C(n_764), .Y(n_780) );
OR4x1_ASAP7_75t_L g781 ( .A(n_773), .B(n_771), .C(n_770), .D(n_718), .Y(n_781) );
INVx3_ASAP7_75t_L g782 ( .A(n_777), .Y(n_782) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_772), .A2(n_729), .B(n_767), .Y(n_783) );
O2A1O1Ixp33_ASAP7_75t_SL g784 ( .A1(n_780), .A2(n_729), .B(n_776), .C(n_774), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_783), .A2(n_775), .B(n_779), .Y(n_785) );
NOR2x1p5_ASAP7_75t_SL g786 ( .A(n_784), .B(n_781), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_785), .B(n_782), .Y(n_787) );
NOR3x1_ASAP7_75t_L g788 ( .A(n_787), .B(n_758), .C(n_730), .Y(n_788) );
NOR3xp33_ASAP7_75t_L g789 ( .A(n_786), .B(n_782), .C(n_738), .Y(n_789) );
INVxp67_ASAP7_75t_L g790 ( .A(n_789), .Y(n_790) );
AND2x4_ASAP7_75t_L g791 ( .A(n_788), .B(n_769), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_791), .Y(n_792) );
INVxp33_ASAP7_75t_L g793 ( .A(n_790), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_792), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_794), .Y(n_795) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_795), .A2(n_793), .B(n_741), .Y(n_796) );
AOI221x1_ASAP7_75t_L g797 ( .A1(n_796), .A2(n_739), .B1(n_721), .B2(n_695), .C(n_743), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_797), .A2(n_734), .B1(n_725), .B2(n_721), .Y(n_798) );
OAI21xp5_ASAP7_75t_L g799 ( .A1(n_798), .A2(n_744), .B(n_711), .Y(n_799) );
OAI21xp5_ASAP7_75t_L g800 ( .A1(n_799), .A2(n_768), .B(n_735), .Y(n_800) );
OR2x6_ASAP7_75t_L g801 ( .A(n_800), .B(n_722), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_801), .A2(n_768), .B1(n_723), .B2(n_720), .Y(n_802) );
endmodule