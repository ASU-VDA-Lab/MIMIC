module fake_jpeg_3320_n_152 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_12),
.B(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_34),
.B(n_33),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_60),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_58),
.Y(n_66)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

CKINVDCx12_ASAP7_75t_R g67 ( 
.A(n_61),
.Y(n_67)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_62),
.B(n_46),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_43),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_47),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_48),
.B1(n_45),
.B2(n_41),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_72),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_69),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_48),
.B1(n_54),
.B2(n_40),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_77),
.A2(n_82),
.B1(n_53),
.B2(n_1),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_40),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_1),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_61),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_80),
.B(n_0),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_49),
.B1(n_44),
.B2(n_53),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_61),
.B1(n_38),
.B2(n_59),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_84),
.A2(n_79),
.B1(n_73),
.B2(n_80),
.Y(n_89)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_72),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_61),
.B1(n_53),
.B2(n_38),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_103),
.B1(n_9),
.B2(n_10),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_2),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_7),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_76),
.B(n_0),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_98),
.B(n_100),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_99),
.A2(n_75),
.B(n_3),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_79),
.A2(n_76),
.B1(n_3),
.B2(n_4),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_91),
.B1(n_102),
.B2(n_15),
.Y(n_123)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_117),
.Y(n_122)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_112),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_120),
.B1(n_121),
.B2(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_30),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_29),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_116),
.B(n_13),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_8),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_119),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_28),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_132),
.B1(n_116),
.B2(n_109),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_19),
.B(n_24),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_128),
.C(n_104),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_129),
.B(n_120),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_115),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_14),
.B1(n_27),
.B2(n_26),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_134),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_130),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_138),
.A2(n_130),
.B(n_122),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_140),
.B1(n_137),
.B2(n_124),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_143),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_125),
.C(n_114),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_131),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_146),
.B(n_128),
.Y(n_147)
);

AO21x1_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_125),
.B(n_145),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_133),
.C(n_137),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

OAI21x1_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_133),
.B(n_119),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_108),
.Y(n_152)
);


endmodule