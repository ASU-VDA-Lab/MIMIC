module real_aes_14258_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_725;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_102;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_397;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
OA21x2_ASAP7_75t_L g111 ( .A1(n_0), .A2(n_44), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g146 ( .A(n_0), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_1), .B(n_140), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_2), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_3), .B(n_196), .Y(n_231) );
BUFx3_ASAP7_75t_L g499 ( .A(n_4), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_5), .A2(n_491), .B1(n_658), .B2(n_659), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_5), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_6), .B(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g678 ( .A(n_6), .Y(n_678) );
INVx3_ASAP7_75t_L g546 ( .A(n_7), .Y(n_546) );
INVx2_ASAP7_75t_L g503 ( .A(n_8), .Y(n_503) );
INVx1_ASAP7_75t_L g533 ( .A(n_8), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_9), .B(n_142), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_10), .B(n_165), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_11), .B(n_254), .Y(n_253) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_11), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_12), .Y(n_175) );
INVx1_ASAP7_75t_L g97 ( .A(n_13), .Y(n_97) );
BUFx3_ASAP7_75t_L g121 ( .A(n_13), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_14), .B(n_128), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_15), .Y(n_225) );
INVxp33_ASAP7_75t_SL g565 ( .A(n_16), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_16), .A2(n_43), .B1(n_622), .B2(n_623), .Y(n_621) );
BUFx10_ASAP7_75t_L g701 ( .A(n_17), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_18), .A2(n_678), .B1(n_679), .B2(n_680), .Y(n_677) );
CKINVDCx5p33_ASAP7_75t_R g679 ( .A(n_18), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g115 ( .A(n_19), .B(n_116), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_20), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_21), .B(n_140), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_22), .B(n_116), .Y(n_126) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_23), .A2(n_58), .B1(n_606), .B2(n_608), .Y(n_605) );
INVx1_ASAP7_75t_L g638 ( .A(n_23), .Y(n_638) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_24), .Y(n_594) );
INVxp33_ASAP7_75t_L g634 ( .A(n_24), .Y(n_634) );
INVx1_ASAP7_75t_L g649 ( .A(n_24), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_25), .B(n_128), .Y(n_266) );
NAND2xp33_ASAP7_75t_L g258 ( .A(n_26), .B(n_120), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g162 ( .A1(n_27), .A2(n_163), .B(n_166), .C(n_168), .Y(n_162) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_27), .Y(n_714) );
INVx1_ASAP7_75t_L g88 ( .A(n_28), .Y(n_88) );
INVx2_ASAP7_75t_L g554 ( .A(n_29), .Y(n_554) );
INVxp33_ASAP7_75t_SL g511 ( .A(n_30), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_30), .A2(n_76), .B1(n_643), .B2(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g516 ( .A(n_31), .Y(n_516) );
OAI211xp5_ASAP7_75t_L g572 ( .A1(n_31), .A2(n_573), .B(n_574), .C(n_589), .Y(n_572) );
OAI222xp33_ASAP7_75t_L g527 ( .A1(n_32), .A2(n_53), .B1(n_68), .B2(n_528), .C1(n_530), .C2(n_534), .Y(n_527) );
INVx1_ASAP7_75t_L g585 ( .A(n_32), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_33), .B(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_34), .B(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g575 ( .A(n_35), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_36), .B(n_194), .Y(n_193) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_37), .Y(n_556) );
INVx2_ASAP7_75t_L g562 ( .A(n_37), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_37), .B(n_649), .Y(n_648) );
AO221x1_ASAP7_75t_L g133 ( .A1(n_38), .A2(n_65), .B1(n_116), .B2(n_123), .C(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_39), .B(n_190), .Y(n_227) );
AND2x4_ASAP7_75t_L g87 ( .A(n_40), .B(n_88), .Y(n_87) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_40), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g270 ( .A(n_41), .B(n_168), .C(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g504 ( .A(n_42), .Y(n_504) );
INVx1_ASAP7_75t_L g521 ( .A(n_42), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_43), .A2(n_51), .B1(n_643), .B2(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g147 ( .A(n_44), .Y(n_147) );
INVx1_ASAP7_75t_L g112 ( .A(n_45), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_46), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_47), .A2(n_202), .B(n_203), .C(n_205), .Y(n_201) );
INVx2_ASAP7_75t_L g204 ( .A(n_48), .Y(n_204) );
INVx1_ASAP7_75t_L g494 ( .A(n_49), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_50), .B(n_110), .Y(n_233) );
INVxp67_ASAP7_75t_SL g618 ( .A(n_51), .Y(n_618) );
OAI21xp33_ASAP7_75t_L g549 ( .A1(n_52), .A2(n_550), .B(n_557), .Y(n_549) );
INVx1_ASAP7_75t_L g602 ( .A(n_52), .Y(n_602) );
INVx1_ASAP7_75t_L g652 ( .A(n_53), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_54), .B(n_189), .Y(n_188) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_55), .Y(n_685) );
AND2x2_ASAP7_75t_L g199 ( .A(n_56), .B(n_110), .Y(n_199) );
INVx1_ASAP7_75t_L g150 ( .A(n_57), .Y(n_150) );
INVxp67_ASAP7_75t_SL g641 ( .A(n_58), .Y(n_641) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_59), .Y(n_690) );
OAI22xp33_ASAP7_75t_L g139 ( .A1(n_60), .A2(n_62), .B1(n_140), .B2(n_142), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_61), .B(n_168), .Y(n_268) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_63), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_64), .A2(n_673), .B1(n_674), .B2(n_675), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_64), .Y(n_673) );
AND2x2_ASAP7_75t_L g213 ( .A(n_66), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g92 ( .A(n_67), .Y(n_92) );
BUFx3_ASAP7_75t_L g124 ( .A(n_67), .Y(n_124) );
INVx1_ASAP7_75t_L g138 ( .A(n_67), .Y(n_138) );
INVx1_ASAP7_75t_L g582 ( .A(n_68), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g107 ( .A(n_69), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g558 ( .A(n_70), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_71), .B(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g553 ( .A(n_72), .Y(n_553) );
AND2x2_ASAP7_75t_L g564 ( .A(n_72), .B(n_554), .Y(n_564) );
INVxp67_ASAP7_75t_SL g588 ( .A(n_72), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_73), .B(n_190), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_74), .B(n_110), .Y(n_259) );
INVx2_ASAP7_75t_L g543 ( .A(n_75), .Y(n_543) );
INVxp67_ASAP7_75t_SL g505 ( .A(n_76), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_77), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_98), .B(n_489), .Y(n_78) );
CKINVDCx6p67_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
CKINVDCx11_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
BUFx6f_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_89), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
BUFx2_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx3_ASAP7_75t_L g131 ( .A(n_87), .Y(n_131) );
INVx2_ASAP7_75t_L g160 ( .A(n_87), .Y(n_160) );
BUFx6f_ASAP7_75t_SL g232 ( .A(n_87), .Y(n_232) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_88), .Y(n_666) );
AO21x2_ASAP7_75t_L g726 ( .A1(n_89), .A2(n_665), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g89 ( .A(n_90), .B(n_93), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
AOI21xp5_ASAP7_75t_SL g186 ( .A1(n_91), .A2(n_187), .B(n_188), .Y(n_186) );
BUFx3_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g198 ( .A(n_92), .Y(n_198) );
HB1xp67_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx1_ASAP7_75t_L g173 ( .A(n_96), .Y(n_173) );
INVx2_ASAP7_75t_L g210 ( .A(n_96), .Y(n_210) );
INVx2_ASAP7_75t_L g230 ( .A(n_96), .Y(n_230) );
INVx2_ASAP7_75t_L g271 ( .A(n_96), .Y(n_271) );
BUFx6f_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx2_ASAP7_75t_L g117 ( .A(n_97), .Y(n_117) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x4_ASAP7_75t_L g99 ( .A(n_100), .B(n_390), .Y(n_99) );
NOR3xp33_ASAP7_75t_SL g100 ( .A(n_101), .B(n_292), .C(n_329), .Y(n_100) );
OAI211xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_152), .B(n_234), .C(n_282), .Y(n_101) );
AOI321xp33_ASAP7_75t_L g468 ( .A1(n_102), .A2(n_382), .A3(n_436), .B1(n_469), .B2(n_471), .C(n_473), .Y(n_468) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_103), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_103), .B(n_410), .Y(n_417) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_132), .Y(n_103) );
INVx1_ASAP7_75t_L g333 ( .A(n_104), .Y(n_333) );
INVx1_ASAP7_75t_L g357 ( .A(n_104), .Y(n_357) );
AND2x2_ASAP7_75t_L g373 ( .A(n_104), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_105), .B(n_261), .Y(n_281) );
AND2x2_ASAP7_75t_L g302 ( .A(n_105), .B(n_132), .Y(n_302) );
INVx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g246 ( .A(n_106), .B(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g287 ( .A(n_106), .B(n_132), .Y(n_287) );
AND2x2_ASAP7_75t_L g344 ( .A(n_106), .B(n_248), .Y(n_344) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_113), .Y(n_106) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_110), .B(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g185 ( .A(n_110), .Y(n_185) );
INVx1_ASAP7_75t_L g250 ( .A(n_110), .Y(n_250) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g215 ( .A(n_111), .Y(n_215) );
BUFx2_ASAP7_75t_L g218 ( .A(n_111), .Y(n_218) );
INVx1_ASAP7_75t_L g148 ( .A(n_112), .Y(n_148) );
OAI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_125), .B(n_130), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_118), .B(n_122), .Y(n_114) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx3_ASAP7_75t_L g165 ( .A(n_117), .Y(n_165) );
INVx2_ASAP7_75t_L g269 ( .A(n_119), .Y(n_269) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx3_ASAP7_75t_L g128 ( .A(n_120), .Y(n_128) );
INVx3_ASAP7_75t_L g134 ( .A(n_120), .Y(n_134) );
INVx2_ASAP7_75t_L g196 ( .A(n_120), .Y(n_196) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g141 ( .A(n_121), .Y(n_141) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_121), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g170 ( .A1(n_122), .A2(n_171), .B(n_174), .Y(n_170) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g129 ( .A(n_124), .Y(n_129) );
INVx2_ASAP7_75t_L g168 ( .A(n_124), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B(n_129), .Y(n_125) );
O2A1O1Ixp5_ASAP7_75t_L g224 ( .A1(n_129), .A2(n_225), .B(n_226), .C(n_227), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_129), .A2(n_265), .B(n_266), .Y(n_264) );
NOR2xp33_ASAP7_75t_R g144 ( .A(n_131), .B(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g184 ( .A(n_131), .Y(n_184) );
AND2x2_ASAP7_75t_L g260 ( .A(n_132), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g280 ( .A(n_132), .B(n_247), .Y(n_280) );
BUFx3_ASAP7_75t_L g336 ( .A(n_132), .Y(n_336) );
INVx2_ASAP7_75t_SL g374 ( .A(n_132), .Y(n_374) );
AND2x2_ASAP7_75t_L g470 ( .A(n_132), .B(n_425), .Y(n_470) );
AO31x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_135), .A3(n_144), .B(n_149), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_139), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_137), .A2(n_253), .B(n_255), .Y(n_252) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx3_ASAP7_75t_L g206 ( .A(n_138), .Y(n_206) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g190 ( .A(n_141), .Y(n_190) );
INVx2_ASAP7_75t_L g194 ( .A(n_141), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_142), .B(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g254 ( .A(n_143), .Y(n_254) );
INVx2_ASAP7_75t_L g151 ( .A(n_145), .Y(n_151) );
AOI21x1_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_148), .Y(n_145) );
AO21x2_ASAP7_75t_L g158 ( .A1(n_146), .A2(n_147), .B(n_148), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_178), .Y(n_153) );
OR2x2_ASAP7_75t_L g306 ( .A(n_154), .B(n_275), .Y(n_306) );
AND2x2_ASAP7_75t_L g308 ( .A(n_154), .B(n_309), .Y(n_308) );
INVx5_ASAP7_75t_L g313 ( .A(n_154), .Y(n_313) );
AND2x4_ASAP7_75t_L g341 ( .A(n_154), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g351 ( .A(n_154), .B(n_328), .Y(n_351) );
AND2x2_ASAP7_75t_L g378 ( .A(n_154), .B(n_336), .Y(n_378) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVxp67_ASAP7_75t_L g323 ( .A(n_155), .Y(n_323) );
AO21x1_ASAP7_75t_SL g155 ( .A1(n_156), .A2(n_161), .B(n_169), .Y(n_155) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_156), .A2(n_161), .B(n_169), .Y(n_242) );
INVxp67_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
OAI21x1_ASAP7_75t_SL g169 ( .A1(n_157), .A2(n_170), .B(n_176), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
INVx2_ASAP7_75t_L g177 ( .A(n_158), .Y(n_177) );
INVx2_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_165), .B(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
INVx1_ASAP7_75t_L g725 ( .A(n_172), .Y(n_725) );
INVx1_ASAP7_75t_L g202 ( .A(n_173), .Y(n_202) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
OR2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_219), .Y(n_179) );
INVx1_ASAP7_75t_L g237 ( .A(n_180), .Y(n_237) );
INVx2_ASAP7_75t_L g338 ( .A(n_180), .Y(n_338) );
OR2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_200), .Y(n_180) );
INVx2_ASAP7_75t_L g244 ( .A(n_181), .Y(n_244) );
INVx1_ASAP7_75t_L g298 ( .A(n_181), .Y(n_298) );
AND2x2_ASAP7_75t_L g311 ( .A(n_181), .B(n_221), .Y(n_311) );
AND2x2_ASAP7_75t_L g324 ( .A(n_181), .B(n_220), .Y(n_324) );
NAND2x1p5_ASAP7_75t_L g181 ( .A(n_182), .B(n_191), .Y(n_181) );
NAND2x1_ASAP7_75t_L g182 ( .A(n_183), .B(n_186), .Y(n_182) );
AOI21x1_ASAP7_75t_L g191 ( .A1(n_183), .A2(n_192), .B(n_199), .Y(n_191) );
O2A1O1Ixp5_ASAP7_75t_L g263 ( .A1(n_183), .A2(n_264), .B(n_267), .C(n_272), .Y(n_263) );
AND2x4_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
AOI21xp33_ASAP7_75t_L g216 ( .A1(n_184), .A2(n_213), .B(n_217), .Y(n_216) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_184), .A2(n_252), .B(n_256), .Y(n_251) );
INVx2_ASAP7_75t_SL g189 ( .A(n_190), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_195), .B(n_197), .Y(n_192) );
INVx1_ASAP7_75t_L g212 ( .A(n_197), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_197), .A2(n_229), .B(n_231), .Y(n_228) );
BUFx10_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g276 ( .A(n_200), .Y(n_276) );
AND2x2_ASAP7_75t_L g328 ( .A(n_200), .B(n_244), .Y(n_328) );
AND2x2_ASAP7_75t_L g342 ( .A(n_200), .B(n_243), .Y(n_342) );
INVx1_ASAP7_75t_L g349 ( .A(n_200), .Y(n_349) );
AND2x2_ASAP7_75t_L g384 ( .A(n_200), .B(n_241), .Y(n_384) );
INVx1_ASAP7_75t_L g404 ( .A(n_200), .Y(n_404) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_207), .B(n_216), .Y(n_200) );
NOR2xp67_ASAP7_75t_L g203 ( .A(n_202), .B(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_206), .A2(n_257), .B(n_258), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_212), .B(n_213), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_211), .Y(n_208) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_217), .B(n_273), .Y(n_272) );
INVxp67_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
BUFx3_ASAP7_75t_L g222 ( .A(n_218), .Y(n_222) );
AND2x2_ASAP7_75t_L g297 ( .A(n_219), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g370 ( .A(n_219), .Y(n_370) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g277 ( .A(n_220), .Y(n_277) );
INVx1_ASAP7_75t_L g350 ( .A(n_220), .Y(n_350) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVxp33_ASAP7_75t_L g315 ( .A(n_221), .Y(n_315) );
OAI21x1_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_233), .Y(n_221) );
OAI21x1_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_228), .B(n_232), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_245), .B1(n_274), .B2(n_278), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_238), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x4_ASAP7_75t_SL g366 ( .A(n_237), .B(n_350), .Y(n_366) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_243), .Y(n_239) );
INVx2_ASAP7_75t_L g327 ( .A(n_240), .Y(n_327) );
BUFx2_ASAP7_75t_SL g483 ( .A(n_240), .Y(n_483) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g290 ( .A(n_241), .B(n_276), .Y(n_290) );
AND2x2_ASAP7_75t_L g438 ( .A(n_241), .B(n_276), .Y(n_438) );
AND2x2_ASAP7_75t_L g445 ( .A(n_241), .B(n_315), .Y(n_445) );
INVx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g296 ( .A(n_242), .B(n_277), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_242), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g291 ( .A(n_243), .B(n_277), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_243), .B(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x4_ASAP7_75t_L g245 ( .A(n_246), .B(n_260), .Y(n_245) );
AND2x4_ASAP7_75t_L g469 ( .A(n_246), .B(n_470), .Y(n_469) );
NAND2x1_ASAP7_75t_L g488 ( .A(n_246), .B(n_424), .Y(n_488) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g286 ( .A(n_248), .Y(n_286) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_248), .Y(n_358) );
INVx1_ASAP7_75t_L g363 ( .A(n_248), .Y(n_363) );
AND2x2_ASAP7_75t_L g389 ( .A(n_248), .B(n_262), .Y(n_389) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_251), .B(n_259), .Y(n_248) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g385 ( .A(n_260), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g425 ( .A(n_261), .Y(n_425) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_262), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g319 ( .A(n_262), .Y(n_319) );
BUFx2_ASAP7_75t_SL g376 ( .A(n_262), .Y(n_376) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_269), .B(n_270), .Y(n_267) );
INVxp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_L g295 ( .A(n_276), .Y(n_295) );
AND2x2_ASAP7_75t_L g314 ( .A(n_276), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g430 ( .A(n_277), .B(n_349), .Y(n_430) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_279), .A2(n_321), .B(n_325), .Y(n_320) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx2_ASAP7_75t_L g364 ( .A(n_281), .Y(n_364) );
OR2x2_ASAP7_75t_L g405 ( .A(n_281), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_288), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_283), .A2(n_421), .B1(n_422), .B2(n_427), .Y(n_420) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx2_ASAP7_75t_L g303 ( .A(n_285), .Y(n_303) );
BUFx2_ASAP7_75t_L g383 ( .A(n_285), .Y(n_383) );
INVx1_ASAP7_75t_L g412 ( .A(n_287), .Y(n_412) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
OR2x2_ASAP7_75t_L g418 ( .A(n_290), .B(n_419), .Y(n_418) );
NAND3xp33_ASAP7_75t_L g292 ( .A(n_293), .B(n_304), .C(n_307), .Y(n_292) );
OAI21xp33_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_297), .B(n_299), .Y(n_293) );
INVx1_ASAP7_75t_L g450 ( .A(n_294), .Y(n_450) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NAND2x1_ASAP7_75t_L g480 ( .A(n_295), .B(n_309), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_297), .B(n_313), .Y(n_416) );
INVx3_ASAP7_75t_L g399 ( .A(n_298), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_299), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AND2x4_ASAP7_75t_L g388 ( .A(n_302), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g426 ( .A(n_302), .Y(n_426) );
AND2x2_ASAP7_75t_L g477 ( .A(n_302), .B(n_319), .Y(n_477) );
AND2x2_ASAP7_75t_L g372 ( .A(n_303), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g454 ( .A(n_303), .B(n_374), .Y(n_454) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AOI21xp33_ASAP7_75t_L g484 ( .A1(n_306), .A2(n_485), .B(n_488), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_312), .B(n_316), .C(n_320), .Y(n_307) );
INVx6_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND4xp25_ASAP7_75t_L g427 ( .A(n_310), .B(n_428), .C(n_431), .D(n_433), .Y(n_427) );
AOI211xp5_ASAP7_75t_L g473 ( .A1(n_310), .A2(n_384), .B(n_474), .C(n_476), .Y(n_473) );
INVx4_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g387 ( .A(n_311), .B(n_384), .Y(n_387) );
INVx2_ASAP7_75t_L g465 ( .A(n_312), .Y(n_465) );
AND2x4_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AND2x2_ASAP7_75t_L g337 ( .A(n_313), .B(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g421 ( .A(n_313), .B(n_366), .Y(n_421) );
AND2x2_ASAP7_75t_L g432 ( .A(n_313), .B(n_342), .Y(n_432) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g461 ( .A(n_318), .Y(n_461) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_319), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g343 ( .A(n_319), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_322), .Y(n_456) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
NAND2x1p5_ASAP7_75t_L g459 ( .A(n_323), .B(n_399), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_324), .B(n_384), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_324), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
OR2x2_ASAP7_75t_L g440 ( .A(n_327), .B(n_348), .Y(n_440) );
INVx1_ASAP7_75t_L g371 ( .A(n_328), .Y(n_371) );
NAND4xp25_ASAP7_75t_SL g329 ( .A(n_330), .B(n_345), .C(n_367), .D(n_377), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_337), .B(n_339), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g359 ( .A1(n_332), .A2(n_360), .B(n_365), .Y(n_359) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g354 ( .A(n_336), .Y(n_354) );
INVx1_ASAP7_75t_L g396 ( .A(n_336), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_336), .B(n_344), .Y(n_415) );
OAI322xp33_ASAP7_75t_L g457 ( .A1(n_336), .A2(n_458), .A3(n_461), .B1(n_462), .B2(n_464), .C1(n_465), .C2(n_466), .Y(n_457) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_336), .Y(n_482) );
INVx1_ASAP7_75t_L g433 ( .A(n_337), .Y(n_433) );
INVx1_ASAP7_75t_L g381 ( .A(n_338), .Y(n_381) );
AND2x2_ASAP7_75t_L g444 ( .A(n_338), .B(n_445), .Y(n_444) );
INVxp67_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_342), .B(n_463), .Y(n_462) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_343), .A2(n_479), .B1(n_481), .B2(n_483), .C(n_484), .Y(n_478) );
AND2x2_ASAP7_75t_L g375 ( .A(n_344), .B(n_376), .Y(n_375) );
BUFx2_ASAP7_75t_L g386 ( .A(n_344), .Y(n_386) );
AND2x4_ASAP7_75t_SL g467 ( .A(n_344), .B(n_374), .Y(n_467) );
O2A1O1Ixp5_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_351), .B(n_352), .C(n_359), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_346), .A2(n_368), .B1(n_372), .B2(n_375), .Y(n_367) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_350), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g463 ( .A(n_350), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_350), .B(n_384), .Y(n_472) );
INVxp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVxp67_ASAP7_75t_L g449 ( .A(n_354), .Y(n_449) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_356), .B(n_396), .Y(n_464) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
OR2x2_ASAP7_75t_L g447 ( .A(n_358), .B(n_425), .Y(n_447) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g481 ( .A(n_361), .B(n_482), .Y(n_481) );
AND2x4_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .Y(n_361) );
INVx2_ASAP7_75t_SL g410 ( .A(n_362), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_362), .B(n_411), .Y(n_441) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_363), .B(n_374), .Y(n_406) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI321xp33_ASAP7_75t_L g407 ( .A1(n_368), .A2(n_408), .A3(n_410), .B1(n_411), .B2(n_413), .C(n_414), .Y(n_407) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
AND2x2_ASAP7_75t_L g401 ( .A(n_370), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g419 ( .A(n_370), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_375), .B(n_395), .Y(n_394) );
AOI322xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .A3(n_382), .B1(n_384), .B2(n_385), .C1(n_387), .C2(n_388), .Y(n_377) );
AOI21xp33_ASAP7_75t_L g392 ( .A1(n_379), .A2(n_393), .B(n_397), .Y(n_392) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
O2A1O1Ixp33_ASAP7_75t_L g397 ( .A1(n_384), .A2(n_398), .B(n_400), .C(n_405), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_385), .A2(n_452), .B1(n_455), .B2(n_456), .C(n_457), .Y(n_451) );
NOR2xp67_ASAP7_75t_L g390 ( .A(n_391), .B(n_434), .Y(n_390) );
NAND3xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_407), .C(n_420), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g446 ( .A(n_396), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x4_ASAP7_75t_L g455 ( .A(n_399), .B(n_430), .Y(n_455) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g475 ( .A(n_402), .Y(n_475) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_403), .Y(n_487) );
INVx1_ASAP7_75t_L g413 ( .A(n_405), .Y(n_413) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI22xp33_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_416), .B1(n_417), .B2(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_426), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g460 ( .A(n_430), .Y(n_460) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND4xp25_ASAP7_75t_L g434 ( .A(n_435), .B(n_451), .C(n_468), .D(n_478), .Y(n_434) );
O2A1O1Ixp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_439), .B(n_441), .C(n_442), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_446), .B1(n_448), .B2(n_450), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g448 ( .A(n_447), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
OR2x2_ASAP7_75t_L g474 ( .A(n_463), .B(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OAI221xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B1(n_660), .B2(n_669), .C(n_721), .Y(n_489) );
INVx2_ASAP7_75t_L g659 ( .A(n_491), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_491), .A2(n_722), .B1(n_725), .B2(n_726), .Y(n_721) );
NOR2x1_ASAP7_75t_L g491 ( .A(n_492), .B(n_547), .Y(n_491) );
AOI31xp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_510), .A3(n_523), .B(n_538), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_505), .B2(n_506), .Y(n_493) );
OAI221xp5_ASAP7_75t_SL g650 ( .A1(n_494), .A2(n_651), .B1(n_652), .B2(n_653), .C(n_656), .Y(n_650) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_500), .Y(n_495) );
AND2x4_ASAP7_75t_L g512 ( .A(n_496), .B(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_SL g517 ( .A(n_496), .B(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g524 ( .A(n_497), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g614 ( .A(n_498), .B(n_542), .Y(n_614) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g507 ( .A(n_499), .Y(n_507) );
AND2x4_ASAP7_75t_L g628 ( .A(n_499), .B(n_542), .Y(n_628) );
OR2x2_ASAP7_75t_L g703 ( .A(n_499), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g713 ( .A(n_499), .B(n_704), .Y(n_713) );
INVx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g509 ( .A(n_502), .Y(n_509) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_502), .Y(n_607) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
AND2x2_ASAP7_75t_L g514 ( .A(n_503), .B(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g522 ( .A(n_503), .Y(n_522) );
INVx2_ASAP7_75t_L g515 ( .A(n_504), .Y(n_515) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
AND2x4_ASAP7_75t_L g531 ( .A(n_507), .B(n_532), .Y(n_531) );
AND2x4_ASAP7_75t_L g535 ( .A(n_507), .B(n_536), .Y(n_535) );
INVx5_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_516), .B2(n_517), .Y(n_510) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g610 ( .A(n_514), .Y(n_610) );
AND2x4_ASAP7_75t_L g526 ( .A(n_515), .B(n_522), .Y(n_526) );
INVx1_ASAP7_75t_L g537 ( .A(n_515), .Y(n_537) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx4_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_520), .Y(n_601) );
AND2x4_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
AND2x4_ASAP7_75t_L g617 ( .A(n_521), .B(n_533), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_524), .B(n_527), .Y(n_523) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_525), .Y(n_604) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_526), .Y(n_529) );
INVx1_ASAP7_75t_L g620 ( .A(n_528), .Y(n_620) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
CKINVDCx14_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
NAND3xp33_ASAP7_75t_L g699 ( .A(n_532), .B(n_700), .C(n_702), .Y(n_699) );
AND2x4_ASAP7_75t_L g710 ( .A(n_532), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
CKINVDCx8_ASAP7_75t_R g534 ( .A(n_535), .Y(n_534) );
INVx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_540), .B(n_544), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g704 ( .A(n_543), .Y(n_704) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g595 ( .A(n_545), .Y(n_595) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g613 ( .A(n_546), .Y(n_613) );
INVx1_ASAP7_75t_L g627 ( .A(n_546), .Y(n_627) );
AND3x1_ASAP7_75t_L g632 ( .A(n_546), .B(n_633), .C(n_634), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_596), .Y(n_547) );
OAI21xp5_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_572), .B(n_591), .Y(n_548) );
OR2x2_ASAP7_75t_SL g550 ( .A(n_551), .B(n_555), .Y(n_550) );
OR2x6_ASAP7_75t_L g573 ( .A(n_551), .B(n_560), .Y(n_573) );
INVx1_ASAP7_75t_L g637 ( .A(n_551), .Y(n_637) );
BUFx3_ASAP7_75t_L g651 ( .A(n_551), .Y(n_651) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
AND2x4_ASAP7_75t_L g570 ( .A(n_553), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g581 ( .A(n_553), .Y(n_581) );
INVx2_ASAP7_75t_L g571 ( .A(n_554), .Y(n_571) );
INVx2_ASAP7_75t_L g580 ( .A(n_554), .Y(n_580) );
INVx3_ASAP7_75t_R g567 ( .A(n_555), .Y(n_567) );
AND2x4_ASAP7_75t_L g590 ( .A(n_555), .B(n_579), .Y(n_590) );
BUFx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B1(n_565), .B2(n_566), .Y(n_557) );
OAI221xp5_ASAP7_75t_L g598 ( .A1(n_558), .A2(n_599), .B1(n_602), .B2(n_603), .C(n_605), .Y(n_598) );
AND2x2_ASAP7_75t_SL g559 ( .A(n_560), .B(n_563), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x4_ASAP7_75t_L g583 ( .A(n_561), .B(n_584), .Y(n_583) );
AND2x4_ASAP7_75t_SL g586 ( .A(n_561), .B(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g633 ( .A(n_561), .Y(n_633) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx12f_ASAP7_75t_SL g640 ( .A(n_563), .Y(n_640) );
BUFx3_ASAP7_75t_L g657 ( .A(n_563), .Y(n_657) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x4_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx4_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx5_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_570), .Y(n_644) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_571), .Y(n_584) );
AOI222xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B1(n_582), .B2(n_583), .C1(n_585), .C2(n_586), .Y(n_574) );
OAI221xp5_ASAP7_75t_SL g615 ( .A1(n_575), .A2(n_616), .B1(n_618), .B2(n_619), .C(n_621), .Y(n_615) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
BUFx4f_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx2_ASAP7_75t_L g645 ( .A(n_579), .Y(n_645) );
AND2x4_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2x1p5_ASAP7_75t_L g655 ( .A(n_580), .B(n_581), .Y(n_655) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
CKINVDCx8_ASAP7_75t_R g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_629), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_611), .B1(n_615), .B2(n_625), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g624 ( .A(n_601), .Y(n_624) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
BUFx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx5_ASAP7_75t_L g622 ( .A(n_610), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_612), .Y(n_611) );
AND2x6_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
OR2x6_ASAP7_75t_L g647 ( .A(n_613), .B(n_648), .Y(n_647) );
INVx8_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x6_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_635), .B1(n_646), .B2(n_650), .Y(n_629) );
BUFx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI221xp5_ASAP7_75t_SL g635 ( .A1(n_636), .A2(n_638), .B1(n_639), .B2(n_641), .C(n_642), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
BUFx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
BUFx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_661), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_662), .Y(n_661) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_667), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
BUFx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g697 ( .A(n_666), .Y(n_697) );
AND2x2_ASAP7_75t_L g727 ( .A(n_667), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_668), .B(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_693), .B1(n_714), .B2(n_715), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_670), .A2(n_714), .B1(n_723), .B2(n_724), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_682), .B1(n_683), .B2(n_692), .Y(n_670) );
INVx1_ASAP7_75t_L g692 ( .A(n_671), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_676), .B1(n_677), .B2(n_681), .Y(n_671) );
INVx1_ASAP7_75t_L g681 ( .A(n_672), .Y(n_681) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g680 ( .A(n_678), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_685), .B1(n_686), .B2(n_687), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B1(n_690), .B2(n_691), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_690), .Y(n_691) );
BUFx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
CKINVDCx16_ASAP7_75t_R g723 ( .A(n_694), .Y(n_723) );
AND2x6_ASAP7_75t_L g694 ( .A(n_695), .B(n_705), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_698), .Y(n_695) );
INVxp67_ASAP7_75t_L g719 ( .A(n_696), .Y(n_719) );
INVx1_ASAP7_75t_L g728 ( .A(n_697), .Y(n_728) );
INVxp67_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_699), .B(n_709), .Y(n_720) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
CKINVDCx11_ASAP7_75t_R g707 ( .A(n_701), .Y(n_707) );
BUFx6f_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .Y(n_705) );
CKINVDCx5p33_ASAP7_75t_R g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
BUFx4f_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_717), .Y(n_724) );
INVx4_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
endmodule