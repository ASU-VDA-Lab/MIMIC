module fake_netlist_6_3644_n_1870 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1870);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1870;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1866;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_171;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_70),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_61),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_22),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_28),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_94),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_3),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_22),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_157),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_149),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_136),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_88),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_113),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_106),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_14),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_144),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_134),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_112),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_1),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_12),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_102),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_57),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_53),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_96),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_42),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_35),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_14),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_76),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_109),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_108),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_8),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_48),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_99),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_74),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_7),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_38),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_130),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_11),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_13),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_35),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_37),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_41),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_151),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_154),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_80),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_85),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_166),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_81),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_128),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_84),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_64),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_83),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_118),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_103),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_47),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_153),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_141),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_68),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_18),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_57),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_115),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_122),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_164),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_23),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_66),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_116),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_124),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_49),
.Y(n_242)
);

BUFx8_ASAP7_75t_SL g243 ( 
.A(n_125),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_77),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_47),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_10),
.Y(n_246)
);

BUFx2_ASAP7_75t_SL g247 ( 
.A(n_63),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_158),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_120),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_7),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_55),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_33),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_92),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_169),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_72),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_69),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_37),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_159),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_21),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_63),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_58),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_82),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_10),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_45),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_20),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_27),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_9),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_52),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_139),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_28),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_101),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_42),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_2),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_38),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_17),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_43),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_90),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_93),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_170),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_104),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_19),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_16),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_21),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_32),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_133),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_167),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_129),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_39),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_146),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_100),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_39),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_59),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_49),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_156),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_132),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_9),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_95),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_123),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_110),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_12),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_143),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_24),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_117),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_23),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_3),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_44),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_48),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_40),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_111),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_31),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_25),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_16),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_43),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_67),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_79),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_114),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_54),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_131),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_71),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_44),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_45),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_17),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_161),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_91),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_73),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_0),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_32),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_40),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_147),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_155),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_51),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_65),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_1),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_30),
.Y(n_334)
);

BUFx2_ASAP7_75t_SL g335 ( 
.A(n_168),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_56),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_86),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_15),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_165),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_145),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_197),
.B(n_0),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_207),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_207),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_192),
.B(n_2),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_195),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_207),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_207),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_243),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_201),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_171),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_173),
.B(n_4),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_207),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_177),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_210),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_180),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_210),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_195),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_277),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_181),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_183),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_299),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_210),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_210),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_173),
.B(n_4),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_210),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_185),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_212),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_186),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_189),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_193),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_212),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_212),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_212),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_196),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_200),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_202),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_228),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_287),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_205),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_221),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_212),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_208),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_215),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_216),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_208),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_220),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_224),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_225),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_197),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_211),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_211),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_226),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_227),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_175),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_231),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_232),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_235),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_229),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_229),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_237),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_239),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_311),
.B(n_5),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_242),
.Y(n_403)
);

INVxp33_ASAP7_75t_SL g404 ( 
.A(n_172),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_241),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_242),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_249),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_246),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_253),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_255),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_256),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_246),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_251),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_258),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_260),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_251),
.B(n_5),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_278),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_289),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_260),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_221),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_295),
.Y(n_421)
);

INVxp33_ASAP7_75t_SL g422 ( 
.A(n_174),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_297),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_380),
.B(n_340),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_342),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_230),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_230),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_343),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_343),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_346),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_346),
.Y(n_432)
);

BUFx8_ASAP7_75t_L g433 ( 
.A(n_413),
.Y(n_433)
);

BUFx8_ASAP7_75t_L g434 ( 
.A(n_413),
.Y(n_434)
);

BUFx8_ASAP7_75t_L g435 ( 
.A(n_341),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_347),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_347),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_352),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_339),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_352),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_354),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_377),
.B(n_378),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_361),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_354),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_356),
.B(n_362),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_357),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_356),
.B(n_298),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_362),
.Y(n_448)
);

AND2x6_ASAP7_75t_L g449 ( 
.A(n_363),
.B(n_279),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_363),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_365),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_365),
.B(n_244),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_367),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_367),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_371),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_371),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_372),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_372),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_394),
.B(n_175),
.Y(n_459)
);

AND2x6_ASAP7_75t_L g460 ( 
.A(n_373),
.B(n_279),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_373),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_350),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_381),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_381),
.B(n_309),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_389),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_389),
.Y(n_466)
);

AND2x2_ASAP7_75t_SL g467 ( 
.A(n_351),
.B(n_244),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_382),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_364),
.B(n_279),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_382),
.B(n_385),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_353),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_390),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_385),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_390),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_391),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_391),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_398),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_344),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_398),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_399),
.B(n_314),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_399),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_403),
.B(n_248),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_403),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_406),
.B(n_323),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_406),
.B(n_182),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_408),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_408),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_402),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_404),
.B(n_316),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_422),
.B(n_348),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_412),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_412),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_415),
.B(n_330),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_415),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_419),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_349),
.A2(n_199),
.B1(n_300),
.B2(n_288),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_419),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_341),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_355),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_454),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_489),
.B(n_359),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_445),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_489),
.B(n_360),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_454),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_499),
.B(n_366),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_454),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_368),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_459),
.B(n_345),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_445),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_474),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_445),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_445),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_445),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_432),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_426),
.B(n_182),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_426),
.Y(n_516)
);

BUFx4f_ASAP7_75t_L g517 ( 
.A(n_469),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_424),
.B(n_369),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_437),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_437),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_424),
.B(n_370),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_439),
.B(n_374),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_459),
.B(n_375),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_446),
.B(n_376),
.Y(n_524)
);

INVxp67_ASAP7_75t_R g525 ( 
.A(n_446),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_425),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_467),
.A2(n_245),
.B1(n_322),
.B2(n_282),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_437),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_467),
.A2(n_423),
.B1(n_386),
.B2(n_388),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_437),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_425),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_432),
.Y(n_532)
);

AND3x2_ASAP7_75t_L g533 ( 
.A(n_462),
.B(n_269),
.C(n_248),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_427),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_432),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_427),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_467),
.A2(n_469),
.B1(n_426),
.B2(n_498),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_428),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_L g539 ( 
.A(n_469),
.B(n_379),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_499),
.B(n_383),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_447),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_439),
.B(n_384),
.Y(n_542)
);

BUFx10_ASAP7_75t_L g543 ( 
.A(n_426),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_438),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_433),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_428),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_438),
.Y(n_547)
);

OAI21xp33_ASAP7_75t_SL g548 ( 
.A1(n_498),
.A2(n_485),
.B(n_428),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_429),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_429),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_430),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_426),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_435),
.A2(n_320),
.B1(n_331),
.B2(n_317),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_447),
.B(n_387),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_438),
.Y(n_555)
);

NAND3xp33_ASAP7_75t_L g556 ( 
.A(n_480),
.B(n_396),
.C(n_395),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_464),
.B(n_401),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_435),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_469),
.A2(n_245),
.B1(n_322),
.B2(n_291),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_440),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_440),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_430),
.Y(n_562)
);

CKINVDCx6p67_ASAP7_75t_R g563 ( 
.A(n_442),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_431),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_431),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_436),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_440),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_436),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_437),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_435),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_464),
.B(n_407),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_469),
.A2(n_275),
.B1(n_336),
.B2(n_291),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_448),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_448),
.Y(n_574)
);

BUFx6f_ASAP7_75t_SL g575 ( 
.A(n_469),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_437),
.Y(n_576)
);

INVx6_ASAP7_75t_L g577 ( 
.A(n_437),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_480),
.B(n_409),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_478),
.A2(n_392),
.B1(n_393),
.B2(n_397),
.Y(n_579)
);

INVx6_ASAP7_75t_L g580 ( 
.A(n_444),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_435),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_450),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_443),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_469),
.B(n_410),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_459),
.B(n_414),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_448),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_444),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_469),
.B(n_417),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_478),
.B(n_418),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_451),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_451),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_488),
.B(n_421),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_469),
.B(n_188),
.Y(n_593)
);

OAI22xp33_ASAP7_75t_L g594 ( 
.A1(n_488),
.A2(n_274),
.B1(n_261),
.B2(n_259),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_444),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_451),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_450),
.Y(n_597)
);

OR2x6_ASAP7_75t_L g598 ( 
.A(n_462),
.B(n_247),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_474),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_453),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_453),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_455),
.Y(n_602)
);

AND2x6_ASAP7_75t_L g603 ( 
.A(n_485),
.B(n_269),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_455),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_474),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_471),
.B(n_400),
.Y(n_606)
);

AO22x2_ASAP7_75t_L g607 ( 
.A1(n_485),
.A2(n_247),
.B1(n_336),
.B2(n_276),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_457),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_435),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_457),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_452),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_484),
.B(n_405),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_474),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_433),
.Y(n_614)
);

AO22x2_ASAP7_75t_L g615 ( 
.A1(n_482),
.A2(n_276),
.B1(n_270),
.B2(n_272),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_484),
.B(n_411),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_474),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_458),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_458),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_493),
.B(n_358),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_461),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_471),
.B(n_280),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_493),
.B(n_332),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_474),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_474),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_482),
.A2(n_282),
.B1(n_296),
.B2(n_293),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_444),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_461),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_463),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_490),
.B(n_338),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_463),
.Y(n_631)
);

INVxp33_ASAP7_75t_L g632 ( 
.A(n_496),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_452),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_477),
.B(n_337),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_444),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_433),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_477),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_476),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_477),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_476),
.Y(n_640)
);

INVxp33_ASAP7_75t_SL g641 ( 
.A(n_496),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_476),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_433),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_444),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_476),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_477),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_433),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_434),
.B(n_280),
.Y(n_648)
);

BUFx4f_ASAP7_75t_L g649 ( 
.A(n_476),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_476),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_476),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_441),
.B(n_219),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_517),
.B(n_434),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_541),
.B(n_479),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_526),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_SL g656 ( 
.A(n_553),
.B(n_529),
.C(n_630),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_578),
.B(n_479),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_517),
.B(n_434),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_518),
.B(n_434),
.Y(n_659)
);

NAND3xp33_ASAP7_75t_L g660 ( 
.A(n_527),
.B(n_434),
.C(n_178),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_538),
.B(n_479),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_538),
.B(n_479),
.Y(n_662)
);

NAND2xp33_ASAP7_75t_L g663 ( 
.A(n_603),
.B(n_537),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_509),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_526),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_524),
.B(n_443),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_517),
.B(n_279),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_546),
.B(n_479),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_516),
.B(n_470),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_546),
.B(n_479),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_521),
.B(n_176),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_508),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_508),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_531),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_505),
.B(n_479),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_509),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_507),
.B(n_491),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_522),
.B(n_542),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_552),
.B(n_279),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_511),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_612),
.B(n_179),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_554),
.B(n_491),
.Y(n_682)
);

NOR2x1p5_ASAP7_75t_L g683 ( 
.A(n_614),
.B(n_187),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_557),
.B(n_491),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_511),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_598),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_571),
.B(n_552),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_548),
.B(n_491),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_500),
.B(n_491),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_500),
.B(n_491),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_516),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_515),
.A2(n_482),
.B1(n_452),
.B2(n_325),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_616),
.B(n_191),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_512),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_548),
.B(n_491),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_512),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_L g697 ( 
.A(n_603),
.B(n_286),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_515),
.A2(n_482),
.B1(n_452),
.B2(n_325),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_504),
.B(n_494),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_501),
.B(n_194),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_636),
.B(n_335),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_524),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_504),
.B(n_494),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_523),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_531),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_523),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_502),
.B(n_494),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_534),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_513),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_579),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_502),
.B(n_494),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_620),
.A2(n_335),
.B1(n_217),
.B2(n_482),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_614),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_513),
.B(n_494),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_623),
.B(n_494),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_515),
.B(n_494),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_611),
.Y(n_717)
);

NAND3xp33_ASAP7_75t_L g718 ( 
.A(n_585),
.B(n_203),
.C(n_198),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_611),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_506),
.B(n_470),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_503),
.B(n_204),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_515),
.B(n_452),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_534),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_585),
.B(n_470),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_633),
.Y(n_725)
);

XOR2xp5_ASAP7_75t_L g726 ( 
.A(n_545),
.B(n_75),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_536),
.B(n_473),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_536),
.B(n_473),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_633),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_543),
.B(n_286),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_549),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_549),
.B(n_473),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_525),
.B(n_465),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_550),
.Y(n_734)
);

A2O1A1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_632),
.A2(n_626),
.B(n_270),
.C(n_273),
.Y(n_735)
);

OAI22xp33_ASAP7_75t_L g736 ( 
.A1(n_598),
.A2(n_285),
.B1(n_240),
.B2(n_294),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_550),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_551),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_551),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_562),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_562),
.B(n_473),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_556),
.B(n_213),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_543),
.B(n_286),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_R g744 ( 
.A(n_643),
.B(n_214),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_543),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_593),
.B(n_286),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_540),
.B(n_233),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_564),
.B(n_441),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_603),
.A2(n_254),
.B1(n_329),
.B2(n_324),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_564),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_525),
.B(n_465),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_565),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_565),
.B(n_441),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_R g754 ( 
.A(n_643),
.B(n_234),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_589),
.B(n_250),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_566),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_566),
.B(n_441),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_568),
.B(n_468),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_598),
.Y(n_759)
);

NAND3xp33_ASAP7_75t_L g760 ( 
.A(n_592),
.B(n_252),
.C(n_334),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_568),
.B(n_468),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_582),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_622),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_582),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_506),
.B(n_466),
.Y(n_765)
);

INVx6_ASAP7_75t_L g766 ( 
.A(n_598),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_603),
.A2(n_303),
.B1(n_285),
.B2(n_184),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_597),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_597),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_600),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_583),
.B(n_466),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_584),
.B(n_286),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_588),
.B(n_286),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_600),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_L g775 ( 
.A1(n_637),
.A2(n_240),
.B(n_329),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_634),
.A2(n_481),
.B(n_483),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_601),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_606),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_603),
.A2(n_223),
.B1(n_222),
.B2(n_218),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_601),
.B(n_468),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_602),
.B(n_468),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_572),
.A2(n_273),
.B(n_272),
.C(n_275),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_602),
.B(n_468),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_604),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_637),
.B(n_639),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_604),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_608),
.B(n_468),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_563),
.B(n_472),
.Y(n_788)
);

NAND2xp33_ASAP7_75t_L g789 ( 
.A(n_603),
.B(n_286),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_533),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_639),
.B(n_286),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_553),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_603),
.A2(n_223),
.B1(n_324),
.B2(n_319),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_608),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_558),
.A2(n_303),
.B1(n_319),
.B2(n_318),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_646),
.B(n_184),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_539),
.A2(n_497),
.B(n_495),
.C(n_492),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_610),
.B(n_468),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_610),
.B(n_481),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_510),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_559),
.A2(n_218),
.B1(n_190),
.B2(n_206),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_618),
.B(n_481),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_618),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_619),
.B(n_483),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_594),
.B(n_257),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_619),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_621),
.B(n_483),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_621),
.B(n_487),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_628),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_628),
.B(n_487),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_629),
.B(n_487),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_629),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_646),
.B(n_190),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_648),
.B(n_263),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_631),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_652),
.B(n_206),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_631),
.B(n_444),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_563),
.B(n_264),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_607),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_514),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_514),
.Y(n_821)
);

NAND2xp33_ASAP7_75t_L g822 ( 
.A(n_599),
.B(n_209),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_650),
.B(n_456),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_636),
.B(n_472),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_650),
.B(n_599),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_678),
.A2(n_581),
.B1(n_558),
.B2(n_570),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_745),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_654),
.A2(n_649),
.B(n_520),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_720),
.B(n_647),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_663),
.A2(n_607),
.B1(n_615),
.B2(n_641),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_671),
.B(n_607),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_687),
.A2(n_649),
.B(n_520),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_745),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_681),
.B(n_607),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_693),
.B(n_615),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_731),
.B(n_615),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_739),
.B(n_615),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_675),
.A2(n_649),
.B(n_520),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_669),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_655),
.Y(n_840)
);

AOI21x1_ASAP7_75t_L g841 ( 
.A1(n_772),
.A2(n_613),
.B(n_605),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_664),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_740),
.B(n_570),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_SL g844 ( 
.A(n_713),
.B(n_641),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_663),
.A2(n_647),
.B(n_581),
.C(n_284),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_750),
.B(n_605),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_756),
.B(n_613),
.Y(n_847)
);

NAND2xp33_ASAP7_75t_L g848 ( 
.A(n_745),
.B(n_510),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_677),
.A2(n_528),
.B(n_519),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_657),
.A2(n_528),
.B(n_519),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_682),
.A2(n_684),
.B(n_715),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_688),
.A2(n_625),
.B(n_617),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_704),
.B(n_702),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_769),
.B(n_617),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_688),
.A2(n_638),
.B(n_625),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_695),
.A2(n_640),
.B(n_638),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_666),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_706),
.B(n_609),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_745),
.B(n_609),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_656),
.A2(n_575),
.B1(n_645),
.B2(n_651),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_735),
.A2(n_209),
.B(n_222),
.C(n_236),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_655),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_771),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_672),
.B(n_640),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_770),
.B(n_642),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_774),
.B(n_642),
.Y(n_866)
);

INVx4_ASAP7_75t_L g867 ( 
.A(n_669),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_695),
.A2(n_651),
.B(n_645),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_669),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_691),
.Y(n_870)
);

BUFx4f_ASAP7_75t_L g871 ( 
.A(n_766),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_673),
.B(n_265),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_786),
.B(n_803),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_676),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_772),
.A2(n_535),
.B(n_532),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_806),
.B(n_569),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_809),
.B(n_569),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_773),
.A2(n_535),
.B(n_532),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_724),
.B(n_302),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_722),
.A2(n_716),
.B(n_662),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_680),
.B(n_569),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_661),
.A2(n_528),
.B(n_635),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_773),
.A2(n_561),
.B(n_544),
.Y(n_883)
);

BUFx4f_ASAP7_75t_L g884 ( 
.A(n_766),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_668),
.A2(n_519),
.B(n_635),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_685),
.B(n_694),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_696),
.B(n_644),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_709),
.B(n_644),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_665),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_670),
.A2(n_530),
.B(n_635),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_788),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_819),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_825),
.A2(n_595),
.B(n_576),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_691),
.Y(n_894)
);

NOR3xp33_ASAP7_75t_L g895 ( 
.A(n_805),
.B(n_315),
.C(n_318),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_735),
.A2(n_271),
.B(n_254),
.C(n_262),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_665),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_720),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_707),
.A2(n_595),
.B(n_576),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_707),
.A2(n_595),
.B(n_576),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_711),
.A2(n_530),
.B(n_624),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_674),
.B(n_587),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_705),
.B(n_587),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_691),
.B(n_510),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_720),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_765),
.B(n_475),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_765),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_711),
.A2(n_530),
.B(n_624),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_705),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_785),
.A2(n_544),
.B(n_555),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_708),
.B(n_587),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_733),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_708),
.B(n_644),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_723),
.B(n_627),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_730),
.A2(n_743),
.B(n_697),
.Y(n_915)
);

O2A1O1Ixp33_ASAP7_75t_SL g916 ( 
.A1(n_782),
.A2(n_236),
.B(n_294),
.C(n_262),
.Y(n_916)
);

INVx11_ASAP7_75t_L g917 ( 
.A(n_763),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_659),
.A2(n_575),
.B1(n_290),
.B2(n_315),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_751),
.B(n_302),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_734),
.B(n_627),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_734),
.Y(n_921)
);

BUFx4f_ASAP7_75t_L g922 ( 
.A(n_766),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_730),
.A2(n_510),
.B(n_624),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_737),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_824),
.A2(n_575),
.B1(n_271),
.B2(n_290),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_743),
.A2(n_624),
.B(n_510),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_737),
.B(n_627),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_738),
.B(n_547),
.Y(n_928)
);

NOR2x2_ASAP7_75t_L g929 ( 
.A(n_701),
.B(n_302),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_697),
.A2(n_789),
.B(n_714),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_686),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_789),
.A2(n_624),
.B(n_596),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_752),
.B(n_547),
.Y(n_933)
);

NOR2x1p5_ASAP7_75t_SL g934 ( 
.A(n_752),
.B(n_555),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_SL g935 ( 
.A(n_713),
.B(n_280),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_714),
.A2(n_690),
.B(n_689),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_762),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_762),
.B(n_560),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_764),
.B(n_560),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_765),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_744),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_778),
.B(n_792),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_764),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_814),
.A2(n_283),
.B(n_284),
.C(n_293),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_818),
.B(n_266),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_768),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_785),
.A2(n_667),
.B(n_776),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_700),
.A2(n_721),
.B1(n_729),
.B2(n_725),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_768),
.B(n_561),
.Y(n_949)
);

BUFx8_ASAP7_75t_SL g950 ( 
.A(n_710),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_777),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_777),
.B(n_567),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_699),
.A2(n_596),
.B(n_591),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_784),
.B(n_794),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_755),
.B(n_321),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_784),
.B(n_567),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_703),
.A2(n_591),
.B(n_590),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_667),
.A2(n_590),
.B(n_586),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_794),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_823),
.A2(n_586),
.B(n_573),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_812),
.B(n_573),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_812),
.B(n_815),
.Y(n_962)
);

AOI21x1_ASAP7_75t_L g963 ( 
.A1(n_746),
.A2(n_574),
.B(n_486),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_815),
.B(n_717),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_816),
.A2(n_497),
.B(n_475),
.C(n_495),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_746),
.A2(n_574),
.B(n_492),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_719),
.A2(n_580),
.B1(n_577),
.B2(n_486),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_718),
.B(n_267),
.Y(n_968)
);

BUFx4f_ASAP7_75t_L g969 ( 
.A(n_759),
.Y(n_969)
);

NOR2xp67_ASAP7_75t_L g970 ( 
.A(n_760),
.B(n_660),
.Y(n_970)
);

O2A1O1Ixp5_ASAP7_75t_L g971 ( 
.A1(n_816),
.A2(n_283),
.B(n_296),
.C(n_238),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_747),
.B(n_799),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_802),
.B(n_577),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_790),
.B(n_78),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_744),
.Y(n_975)
);

AOI21xp33_ASAP7_75t_L g976 ( 
.A1(n_742),
.A2(n_268),
.B(n_281),
.Y(n_976)
);

INVx11_ASAP7_75t_L g977 ( 
.A(n_683),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_782),
.A2(n_292),
.B(n_333),
.C(n_304),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_692),
.A2(n_456),
.B(n_577),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_804),
.B(n_577),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_807),
.B(n_580),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_712),
.A2(n_580),
.B1(n_460),
.B2(n_449),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_698),
.A2(n_456),
.B(n_580),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_808),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_820),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_810),
.B(n_456),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_811),
.B(n_456),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_727),
.B(n_456),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_728),
.B(n_456),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_701),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_821),
.Y(n_991)
);

NOR2xp67_ASAP7_75t_L g992 ( 
.A(n_795),
.B(n_150),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_817),
.A2(n_460),
.B(n_449),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_800),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_732),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_741),
.A2(n_460),
.B(n_449),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_775),
.B(n_312),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_748),
.B(n_310),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_753),
.B(n_313),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_754),
.B(n_321),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_800),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_758),
.B(n_301),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_754),
.B(n_321),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_796),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_797),
.A2(n_328),
.B(n_327),
.C(n_326),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_800),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_757),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_796),
.B(n_308),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_653),
.A2(n_658),
.B1(n_701),
.B2(n_767),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_701),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_761),
.A2(n_460),
.B(n_449),
.Y(n_1011)
);

BUFx4f_ASAP7_75t_L g1012 ( 
.A(n_726),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_801),
.A2(n_307),
.B(n_306),
.C(n_305),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_813),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_813),
.B(n_460),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_827),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_851),
.A2(n_658),
.B(n_653),
.Y(n_1017)
);

CKINVDCx10_ASAP7_75t_R g1018 ( 
.A(n_950),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_857),
.B(n_736),
.Y(n_1019)
);

AOI21x1_ASAP7_75t_L g1020 ( 
.A1(n_954),
.A2(n_781),
.B(n_798),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_912),
.B(n_780),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_930),
.A2(n_679),
.B(n_787),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_863),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_912),
.B(n_783),
.Y(n_1024)
);

AO32x1_ASAP7_75t_L g1025 ( 
.A1(n_1009),
.A2(n_822),
.A3(n_679),
.B1(n_791),
.B2(n_779),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_940),
.B(n_793),
.Y(n_1026)
);

BUFx4f_ASAP7_75t_SL g1027 ( 
.A(n_941),
.Y(n_1027)
);

CKINVDCx14_ASAP7_75t_R g1028 ( 
.A(n_1012),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_862),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_880),
.A2(n_791),
.B(n_822),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_862),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_919),
.B(n_301),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_827),
.Y(n_1033)
);

NOR2xp67_ASAP7_75t_SL g1034 ( 
.A(n_827),
.B(n_301),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_895),
.A2(n_749),
.B(n_8),
.C(n_11),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_951),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_SL g1037 ( 
.A1(n_845),
.A2(n_162),
.B(n_160),
.C(n_152),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_945),
.A2(n_6),
.B(n_13),
.C(n_15),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_984),
.B(n_6),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_931),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_915),
.A2(n_460),
.B(n_449),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_827),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_848),
.A2(n_460),
.B(n_449),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_972),
.B(n_18),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_849),
.A2(n_460),
.B(n_449),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_945),
.A2(n_19),
.B(n_20),
.C(n_24),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_R g1047 ( 
.A(n_975),
.B(n_148),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_895),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_842),
.B(n_26),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_942),
.B(n_853),
.Y(n_1050)
);

O2A1O1Ixp5_ASAP7_75t_L g1051 ( 
.A1(n_918),
.A2(n_142),
.B(n_140),
.C(n_135),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_940),
.B(n_127),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_850),
.A2(n_460),
.B(n_449),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_951),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_947),
.A2(n_449),
.B(n_121),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_SL g1056 ( 
.A1(n_968),
.A2(n_107),
.B(n_105),
.C(n_98),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_950),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_940),
.B(n_97),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_897),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_940),
.B(n_89),
.Y(n_1060)
);

AOI22x1_ASAP7_75t_SL g1061 ( 
.A1(n_874),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_833),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_831),
.A2(n_968),
.B(n_942),
.C(n_834),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_976),
.A2(n_29),
.B(n_33),
.C(n_34),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_917),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_891),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_909),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_873),
.B(n_34),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_944),
.A2(n_36),
.B(n_41),
.C(n_46),
.Y(n_1069)
);

NAND2x1_ASAP7_75t_L g1070 ( 
.A(n_833),
.B(n_87),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_838),
.A2(n_36),
.B(n_46),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_969),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_995),
.B(n_1007),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_828),
.A2(n_50),
.B(n_51),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_955),
.B(n_50),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_924),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_962),
.A2(n_52),
.B(n_53),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_832),
.A2(n_54),
.B(n_55),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_909),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_835),
.A2(n_56),
.B(n_58),
.C(n_59),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_948),
.A2(n_830),
.B1(n_869),
.B2(n_886),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_959),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_936),
.A2(n_60),
.B(n_61),
.Y(n_1083)
);

NOR2xp67_ASAP7_75t_SL g1084 ( 
.A(n_833),
.B(n_60),
.Y(n_1084)
);

AND2x2_ASAP7_75t_SL g1085 ( 
.A(n_830),
.B(n_62),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_833),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_997),
.A2(n_1004),
.B(n_1014),
.C(n_970),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_867),
.B(n_62),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_840),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_889),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_871),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_853),
.A2(n_858),
.B(n_872),
.C(n_1005),
.Y(n_1092)
);

NOR3xp33_ASAP7_75t_SL g1093 ( 
.A(n_858),
.B(n_944),
.C(n_978),
.Y(n_1093)
);

NAND2x1p5_ASAP7_75t_L g1094 ( 
.A(n_867),
.B(n_871),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_937),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_882),
.A2(n_890),
.B(n_885),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_SL g1097 ( 
.A1(n_935),
.A2(n_844),
.B1(n_1000),
.B2(n_1003),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_893),
.A2(n_904),
.B(n_900),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_884),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_906),
.B(n_892),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_869),
.A2(n_905),
.B1(n_839),
.B2(n_898),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_932),
.A2(n_980),
.B(n_981),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_943),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_905),
.B(n_907),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_974),
.Y(n_1105)
);

OAI21xp33_ASAP7_75t_L g1106 ( 
.A1(n_872),
.A2(n_879),
.B(n_1008),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_839),
.A2(n_898),
.B1(n_894),
.B2(n_884),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_870),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_894),
.A2(n_922),
.B1(n_843),
.B2(n_907),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_906),
.B(n_892),
.Y(n_1110)
);

OAI21xp33_ASAP7_75t_SL g1111 ( 
.A1(n_954),
.A2(n_964),
.B(n_836),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_946),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_SL g1113 ( 
.A(n_974),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1005),
.A2(n_845),
.B(n_864),
.C(n_837),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_921),
.Y(n_1115)
);

NAND2xp33_ASAP7_75t_SL g1116 ( 
.A(n_1010),
.B(n_990),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_998),
.B(n_999),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_978),
.A2(n_1002),
.B(n_1013),
.C(n_896),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_864),
.B(n_921),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_973),
.A2(n_986),
.B(n_987),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_829),
.A2(n_1002),
.B1(n_1010),
.B2(n_991),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_922),
.B(n_1010),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_1010),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_985),
.B(n_829),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_859),
.A2(n_826),
.B1(n_964),
.B2(n_860),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_969),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_985),
.B(n_1013),
.Y(n_1127)
);

BUFx12f_ASAP7_75t_L g1128 ( 
.A(n_870),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_979),
.A2(n_983),
.B(n_989),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_859),
.B(n_994),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_988),
.A2(n_904),
.B(n_952),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_846),
.Y(n_1132)
);

BUFx8_ASAP7_75t_L g1133 ( 
.A(n_977),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_870),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_870),
.B(n_865),
.Y(n_1135)
);

O2A1O1Ixp5_ASAP7_75t_L g1136 ( 
.A1(n_925),
.A2(n_926),
.B(n_923),
.C(n_961),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_1012),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_SL g1138 ( 
.A1(n_929),
.A2(n_1006),
.B1(n_994),
.B2(n_1001),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_1001),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_1001),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_SL g1141 ( 
.A1(n_1001),
.A2(n_847),
.B1(n_854),
.B2(n_866),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_SL g1142 ( 
.A(n_992),
.B(n_965),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_928),
.B(n_939),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_933),
.A2(n_956),
.B(n_938),
.Y(n_1144)
);

OAI22x1_ASAP7_75t_L g1145 ( 
.A1(n_967),
.A2(n_841),
.B1(n_963),
.B2(n_961),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_876),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_877),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_949),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_881),
.B(n_887),
.Y(n_1149)
);

BUFx2_ASAP7_75t_L g1150 ( 
.A(n_852),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_855),
.A2(n_856),
.B(n_868),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_902),
.B(n_920),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_875),
.A2(n_883),
.B(n_878),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_903),
.A2(n_914),
.B(n_927),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_911),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_971),
.B(n_861),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_958),
.A2(n_957),
.B(n_953),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_913),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_SL g1159 ( 
.A1(n_910),
.A2(n_966),
.B(n_901),
.C(n_908),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_888),
.B(n_1015),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_934),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_899),
.A2(n_960),
.B(n_996),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_971),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_916),
.A2(n_993),
.B(n_1011),
.C(n_982),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_916),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_851),
.A2(n_663),
.B(n_930),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_851),
.A2(n_663),
.B(n_930),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_862),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_948),
.A2(n_678),
.B1(n_972),
.B2(n_687),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_948),
.A2(n_678),
.B1(n_972),
.B2(n_687),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_851),
.A2(n_663),
.B(n_930),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_SL g1172 ( 
.A1(n_945),
.A2(n_641),
.B1(n_496),
.B2(n_710),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_862),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_942),
.B(n_678),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1169),
.A2(n_1170),
.B(n_1174),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1050),
.B(n_1117),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1091),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1092),
.A2(n_1106),
.B(n_1118),
.C(n_1063),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1017),
.A2(n_1167),
.B(n_1166),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1017),
.A2(n_1167),
.B(n_1166),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_SL g1181 ( 
.A(n_1097),
.B(n_1075),
.C(n_1064),
.Y(n_1181)
);

AOI221xp5_ASAP7_75t_SL g1182 ( 
.A1(n_1080),
.A2(n_1046),
.B1(n_1038),
.B2(n_1048),
.C(n_1035),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1073),
.B(n_1132),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1040),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1096),
.A2(n_1098),
.B(n_1162),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_SL g1186 ( 
.A(n_1032),
.B(n_1087),
.C(n_1069),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1091),
.B(n_1172),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1021),
.B(n_1024),
.Y(n_1188)
);

AOI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_1044),
.A2(n_1081),
.B1(n_1093),
.B2(n_1083),
.C(n_1077),
.Y(n_1189)
);

INVx3_ASAP7_75t_SL g1190 ( 
.A(n_1057),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1039),
.A2(n_1088),
.B(n_1049),
.C(n_1068),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1171),
.A2(n_1151),
.B(n_1030),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1083),
.A2(n_1019),
.B(n_1056),
.C(n_1074),
.Y(n_1193)
);

NAND2x1p5_ASAP7_75t_L g1194 ( 
.A(n_1099),
.B(n_1091),
.Y(n_1194)
);

AOI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1085),
.A2(n_1138),
.B1(n_1146),
.B2(n_1116),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1162),
.A2(n_1157),
.B(n_1102),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_SL g1197 ( 
.A1(n_1127),
.A2(n_1052),
.B(n_1058),
.C(n_1060),
.Y(n_1197)
);

AOI221x1_ASAP7_75t_L g1198 ( 
.A1(n_1071),
.A2(n_1074),
.B1(n_1078),
.B2(n_1141),
.C(n_1055),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1105),
.B(n_1100),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1148),
.B(n_1147),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1102),
.A2(n_1129),
.B(n_1171),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1030),
.A2(n_1120),
.B(n_1142),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_1133),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1059),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_1120),
.A2(n_1153),
.A3(n_1055),
.B(n_1150),
.Y(n_1205)
);

O2A1O1Ixp5_ASAP7_75t_L g1206 ( 
.A1(n_1051),
.A2(n_1071),
.B(n_1136),
.C(n_1034),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1153),
.A2(n_1144),
.B(n_1159),
.Y(n_1207)
);

AO21x2_ASAP7_75t_L g1208 ( 
.A1(n_1125),
.A2(n_1022),
.B(n_1131),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1111),
.A2(n_1130),
.B(n_1022),
.Y(n_1209)
);

OAI22x1_ASAP7_75t_L g1210 ( 
.A1(n_1122),
.A2(n_1099),
.B1(n_1082),
.B2(n_1076),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1113),
.A2(n_1124),
.B1(n_1101),
.B2(n_1066),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1027),
.B(n_1110),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1072),
.B(n_1126),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1144),
.A2(n_1143),
.B(n_1154),
.Y(n_1214)
);

NAND3xp33_ASAP7_75t_L g1215 ( 
.A(n_1077),
.B(n_1121),
.C(n_1084),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1131),
.A2(n_1154),
.B(n_1160),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1113),
.A2(n_1107),
.B1(n_1067),
.B2(n_1079),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1023),
.Y(n_1218)
);

INVx6_ASAP7_75t_L g1219 ( 
.A(n_1133),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1139),
.A2(n_1119),
.B1(n_1094),
.B2(n_1135),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_SL g1221 ( 
.A(n_1137),
.B(n_1065),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1155),
.B(n_1158),
.Y(n_1222)
);

INVx4_ASAP7_75t_L g1223 ( 
.A(n_1128),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_SL g1224 ( 
.A1(n_1026),
.A2(n_1165),
.B(n_1070),
.C(n_1104),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_SL g1225 ( 
.A1(n_1149),
.A2(n_1109),
.B(n_1163),
.C(n_1054),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1037),
.A2(n_1164),
.B(n_1123),
.C(n_1089),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1152),
.A2(n_1025),
.B(n_1161),
.Y(n_1227)
);

NAND3xp33_ASAP7_75t_SL g1228 ( 
.A(n_1047),
.B(n_1094),
.C(n_1156),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1090),
.B(n_1095),
.Y(n_1229)
);

INVx5_ASAP7_75t_L g1230 ( 
.A(n_1042),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1042),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1103),
.A2(n_1112),
.B(n_1020),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_SL g1233 ( 
.A1(n_1029),
.A2(n_1173),
.B(n_1036),
.C(n_1031),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1115),
.A2(n_1168),
.B(n_1041),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1161),
.A2(n_1045),
.B(n_1053),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1025),
.A2(n_1043),
.B(n_1134),
.Y(n_1236)
);

INVx4_ASAP7_75t_L g1237 ( 
.A(n_1042),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1028),
.A2(n_1134),
.B1(n_1108),
.B2(n_1016),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1025),
.A2(n_1108),
.A3(n_1016),
.B(n_1033),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1033),
.B(n_1062),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1062),
.Y(n_1241)
);

NOR2xp67_ASAP7_75t_L g1242 ( 
.A(n_1062),
.B(n_1086),
.Y(n_1242)
);

NAND3xp33_ASAP7_75t_SL g1243 ( 
.A(n_1061),
.B(n_1018),
.C(n_1086),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1140),
.A2(n_656),
.B1(n_1174),
.B2(n_1172),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1140),
.B(n_1086),
.Y(n_1245)
);

INVxp67_ASAP7_75t_L g1246 ( 
.A(n_1140),
.Y(n_1246)
);

INVx1_ASAP7_75t_SL g1247 ( 
.A(n_1040),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1174),
.B(n_678),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1072),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1169),
.A2(n_1170),
.B(n_1174),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1059),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1168),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1174),
.A2(n_678),
.B(n_693),
.C(n_681),
.Y(n_1253)
);

AO31x2_ASAP7_75t_L g1254 ( 
.A1(n_1017),
.A2(n_1114),
.A3(n_1145),
.B(n_1151),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1059),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1017),
.A2(n_517),
.B(n_848),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1174),
.B(n_1050),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1017),
.A2(n_1114),
.A3(n_1145),
.B(n_1151),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1174),
.B(n_678),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1072),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1017),
.A2(n_517),
.B(n_848),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1174),
.B(n_1050),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1059),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1169),
.A2(n_1170),
.B(n_1174),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1017),
.A2(n_517),
.B(n_848),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1028),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_SL g1267 ( 
.A1(n_1172),
.A2(n_641),
.B1(n_1174),
.B2(n_1085),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1099),
.B(n_1091),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1040),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1017),
.A2(n_517),
.B(n_848),
.Y(n_1270)
);

AO31x2_ASAP7_75t_L g1271 ( 
.A1(n_1017),
.A2(n_1114),
.A3(n_1145),
.B(n_1151),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1059),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1096),
.A2(n_1098),
.B(n_1162),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1133),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1174),
.B(n_1050),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1017),
.A2(n_1114),
.A3(n_1145),
.B(n_1151),
.Y(n_1276)
);

AO31x2_ASAP7_75t_L g1277 ( 
.A1(n_1017),
.A2(n_1114),
.A3(n_1145),
.B(n_1151),
.Y(n_1277)
);

AND2x2_ASAP7_75t_SL g1278 ( 
.A(n_1085),
.B(n_1174),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_SL g1279 ( 
.A1(n_1169),
.A2(n_658),
.B(n_653),
.Y(n_1279)
);

INVx4_ASAP7_75t_L g1280 ( 
.A(n_1091),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_SL g1281 ( 
.A1(n_1127),
.A2(n_1083),
.B(n_1074),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1174),
.A2(n_1050),
.B1(n_1170),
.B2(n_1169),
.Y(n_1282)
);

O2A1O1Ixp33_ASAP7_75t_SL g1283 ( 
.A1(n_1092),
.A2(n_1063),
.B(n_1087),
.C(n_1114),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1017),
.A2(n_517),
.B(n_848),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1017),
.A2(n_517),
.B(n_848),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1096),
.A2(n_1098),
.B(n_1162),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_SL g1287 ( 
.A1(n_1092),
.A2(n_1063),
.B(n_1087),
.C(n_1114),
.Y(n_1287)
);

NOR2xp67_ASAP7_75t_L g1288 ( 
.A(n_1099),
.B(n_948),
.Y(n_1288)
);

AOI221x1_ASAP7_75t_L g1289 ( 
.A1(n_1174),
.A2(n_895),
.B1(n_1083),
.B2(n_1063),
.C(n_1071),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1174),
.B(n_678),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1151),
.A2(n_1120),
.B(n_1153),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1017),
.A2(n_1114),
.A3(n_1145),
.B(n_1151),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1174),
.B(n_678),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1174),
.A2(n_678),
.B(n_693),
.C(n_681),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1096),
.A2(n_1098),
.B(n_1162),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1174),
.B(n_678),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1174),
.A2(n_1172),
.B1(n_656),
.B2(n_1050),
.Y(n_1297)
);

OR2x6_ASAP7_75t_L g1298 ( 
.A(n_1099),
.B(n_1094),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1174),
.B(n_678),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1174),
.A2(n_678),
.B(n_693),
.C(n_681),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1017),
.A2(n_517),
.B(n_848),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1174),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1017),
.A2(n_1114),
.A3(n_1145),
.B(n_1151),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1099),
.B(n_1091),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1017),
.A2(n_517),
.B(n_848),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1059),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1096),
.A2(n_1098),
.B(n_1162),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1040),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1017),
.A2(n_517),
.B(n_848),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1017),
.A2(n_517),
.B(n_848),
.Y(n_1310)
);

AO32x2_ASAP7_75t_L g1311 ( 
.A1(n_1141),
.A2(n_1081),
.A3(n_1170),
.B1(n_1169),
.B2(n_1101),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1096),
.A2(n_1098),
.B(n_1162),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_SL g1313 ( 
.A1(n_1092),
.A2(n_1063),
.B(n_1087),
.C(n_1114),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1174),
.B(n_678),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1017),
.A2(n_517),
.B(n_848),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1059),
.Y(n_1316)
);

AND2x6_ASAP7_75t_L g1317 ( 
.A(n_1042),
.B(n_1062),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_1040),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1174),
.A2(n_678),
.B(n_693),
.C(n_681),
.Y(n_1319)
);

AO22x2_ASAP7_75t_L g1320 ( 
.A1(n_1169),
.A2(n_656),
.B1(n_895),
.B2(n_1170),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1017),
.A2(n_1114),
.A3(n_1145),
.B(n_1151),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1040),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1072),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1059),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1059),
.Y(n_1325)
);

INVx5_ASAP7_75t_L g1326 ( 
.A(n_1042),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1059),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1168),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1096),
.A2(n_1098),
.B(n_1162),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1151),
.A2(n_1120),
.B(n_1153),
.Y(n_1330)
);

AOI21xp33_ASAP7_75t_L g1331 ( 
.A1(n_1174),
.A2(n_693),
.B(n_681),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1239),
.Y(n_1332)
);

OAI22x1_ASAP7_75t_L g1333 ( 
.A1(n_1297),
.A2(n_1262),
.B1(n_1275),
.B2(n_1257),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1298),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1253),
.A2(n_1300),
.B(n_1294),
.Y(n_1335)
);

CKINVDCx11_ASAP7_75t_R g1336 ( 
.A(n_1190),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_1247),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1278),
.A2(n_1331),
.B1(n_1282),
.B2(n_1297),
.Y(n_1338)
);

OAI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1176),
.A2(n_1314),
.B1(n_1248),
.B2(n_1299),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1259),
.B(n_1290),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_1266),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1267),
.A2(n_1175),
.B1(n_1264),
.B2(n_1250),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1298),
.Y(n_1343)
);

INVx3_ASAP7_75t_L g1344 ( 
.A(n_1298),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1293),
.A2(n_1296),
.B1(n_1319),
.B2(n_1302),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1269),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_SL g1347 ( 
.A(n_1203),
.Y(n_1347)
);

CKINVDCx6p67_ASAP7_75t_R g1348 ( 
.A(n_1274),
.Y(n_1348)
);

INVx2_ASAP7_75t_SL g1349 ( 
.A(n_1213),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1267),
.A2(n_1181),
.B1(n_1320),
.B2(n_1189),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1252),
.Y(n_1351)
);

BUFx12f_ASAP7_75t_L g1352 ( 
.A(n_1219),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1320),
.A2(n_1186),
.B1(n_1244),
.B2(n_1215),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1251),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1183),
.B(n_1188),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_SL g1356 ( 
.A1(n_1215),
.A2(n_1221),
.B1(n_1209),
.B2(n_1200),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1255),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1243),
.A2(n_1288),
.B1(n_1195),
.B2(n_1208),
.Y(n_1358)
);

OAI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1195),
.A2(n_1289),
.B1(n_1222),
.B2(n_1221),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1211),
.A2(n_1178),
.B1(n_1288),
.B2(n_1217),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1263),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1208),
.A2(n_1187),
.B1(n_1281),
.B2(n_1228),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1272),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1202),
.A2(n_1324),
.B1(n_1325),
.B2(n_1306),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1316),
.A2(n_1327),
.B1(n_1210),
.B2(n_1247),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1229),
.Y(n_1366)
);

CKINVDCx12_ASAP7_75t_R g1367 ( 
.A(n_1199),
.Y(n_1367)
);

OAI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1318),
.A2(n_1198),
.B1(n_1322),
.B2(n_1308),
.Y(n_1368)
);

INVx6_ASAP7_75t_L g1369 ( 
.A(n_1230),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1213),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1328),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1191),
.A2(n_1212),
.B(n_1193),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1182),
.A2(n_1268),
.B1(n_1304),
.B2(n_1220),
.Y(n_1373)
);

CKINVDCx6p67_ASAP7_75t_R g1374 ( 
.A(n_1177),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1318),
.A2(n_1238),
.B1(n_1184),
.B2(n_1194),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1268),
.B(n_1304),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_1230),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1218),
.A2(n_1279),
.B1(n_1323),
.B2(n_1260),
.Y(n_1378)
);

CKINVDCx6p67_ASAP7_75t_R g1379 ( 
.A(n_1177),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1245),
.Y(n_1380)
);

BUFx4f_ASAP7_75t_SL g1381 ( 
.A(n_1177),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1237),
.Y(n_1382)
);

CKINVDCx6p67_ASAP7_75t_R g1383 ( 
.A(n_1223),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1230),
.Y(n_1384)
);

INVx3_ASAP7_75t_L g1385 ( 
.A(n_1231),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1192),
.A2(n_1330),
.B1(n_1291),
.B2(n_1179),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_1219),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1233),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1291),
.A2(n_1330),
.B1(n_1180),
.B2(n_1216),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1249),
.A2(n_1246),
.B1(n_1223),
.B2(n_1326),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1231),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1232),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1240),
.Y(n_1393)
);

INVx6_ASAP7_75t_L g1394 ( 
.A(n_1326),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1182),
.A2(n_1313),
.B1(n_1287),
.B2(n_1283),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1231),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1326),
.A2(n_1265),
.B1(n_1305),
.B2(n_1315),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1241),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1239),
.Y(n_1399)
);

OAI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1214),
.A2(n_1227),
.B1(n_1311),
.B2(n_1234),
.Y(n_1400)
);

BUFx4f_ASAP7_75t_SL g1401 ( 
.A(n_1241),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1197),
.A2(n_1224),
.B1(n_1225),
.B2(n_1242),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_SL g1403 ( 
.A1(n_1311),
.A2(n_1284),
.B1(n_1285),
.B2(n_1270),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1239),
.Y(n_1404)
);

BUFx8_ASAP7_75t_L g1405 ( 
.A(n_1241),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1226),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1317),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1311),
.A2(n_1301),
.B1(n_1310),
.B2(n_1309),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1207),
.A2(n_1235),
.B1(n_1236),
.B2(n_1201),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1256),
.A2(n_1261),
.B1(n_1329),
.B2(n_1286),
.Y(n_1410)
);

AOI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1242),
.A2(n_1317),
.B1(n_1185),
.B2(n_1312),
.Y(n_1411)
);

CKINVDCx6p67_ASAP7_75t_R g1412 ( 
.A(n_1317),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1317),
.A2(n_1307),
.B1(n_1295),
.B2(n_1273),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_1205),
.Y(n_1414)
);

INVx3_ASAP7_75t_SL g1415 ( 
.A(n_1206),
.Y(n_1415)
);

CKINVDCx11_ASAP7_75t_R g1416 ( 
.A(n_1205),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1196),
.A2(n_1277),
.B1(n_1254),
.B2(n_1258),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1205),
.A2(n_1254),
.B1(n_1258),
.B2(n_1271),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1271),
.A2(n_1276),
.B1(n_1277),
.B2(n_1292),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1271),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1276),
.A2(n_1277),
.B1(n_1292),
.B2(n_1303),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1292),
.A2(n_1174),
.B1(n_1176),
.B2(n_1299),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1303),
.A2(n_1174),
.B1(n_1176),
.B2(n_1314),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_1303),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1321),
.Y(n_1425)
);

OAI21xp33_ASAP7_75t_L g1426 ( 
.A1(n_1257),
.A2(n_1174),
.B(n_1262),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1257),
.A2(n_1275),
.B1(n_1262),
.B2(n_1172),
.Y(n_1427)
);

CKINVDCx11_ASAP7_75t_R g1428 ( 
.A(n_1190),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1190),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1257),
.A2(n_1275),
.B1(n_1262),
.B2(n_1174),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1204),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1266),
.Y(n_1432)
);

CKINVDCx6p67_ASAP7_75t_R g1433 ( 
.A(n_1190),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1176),
.A2(n_1259),
.B1(n_1290),
.B2(n_1248),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1257),
.A2(n_1275),
.B1(n_1262),
.B2(n_1174),
.Y(n_1435)
);

CKINVDCx11_ASAP7_75t_R g1436 ( 
.A(n_1190),
.Y(n_1436)
);

INVxp67_ASAP7_75t_SL g1437 ( 
.A(n_1226),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1278),
.A2(n_1267),
.B1(n_1257),
.B2(n_1262),
.Y(n_1438)
);

CKINVDCx11_ASAP7_75t_R g1439 ( 
.A(n_1190),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1204),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_SL g1441 ( 
.A(n_1203),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1176),
.A2(n_1259),
.B1(n_1290),
.B2(n_1248),
.Y(n_1442)
);

INVx6_ASAP7_75t_L g1443 ( 
.A(n_1280),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1278),
.A2(n_1267),
.B1(n_1257),
.B2(n_1262),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1257),
.A2(n_1275),
.B1(n_1262),
.B2(n_1174),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_1266),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1204),
.Y(n_1447)
);

BUFx8_ASAP7_75t_L g1448 ( 
.A(n_1177),
.Y(n_1448)
);

AOI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1257),
.A2(n_1275),
.B1(n_1262),
.B2(n_1172),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1269),
.Y(n_1450)
);

CKINVDCx11_ASAP7_75t_R g1451 ( 
.A(n_1190),
.Y(n_1451)
);

CKINVDCx11_ASAP7_75t_R g1452 ( 
.A(n_1190),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1230),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1252),
.Y(n_1454)
);

OAI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1176),
.A2(n_1259),
.B1(n_1290),
.B2(n_1248),
.Y(n_1455)
);

OAI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1176),
.A2(n_1259),
.B1(n_1290),
.B2(n_1248),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1213),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1204),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1213),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1257),
.B(n_1262),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1257),
.B(n_1262),
.Y(n_1461)
);

CKINVDCx8_ASAP7_75t_R g1462 ( 
.A(n_1177),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1257),
.B(n_1262),
.Y(n_1463)
);

AO21x2_ASAP7_75t_L g1464 ( 
.A1(n_1400),
.A2(n_1335),
.B(n_1397),
.Y(n_1464)
);

NOR2x1_ASAP7_75t_SL g1465 ( 
.A(n_1406),
.B(n_1388),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1427),
.A2(n_1449),
.B1(n_1430),
.B2(n_1435),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1410),
.A2(n_1386),
.B(n_1409),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_R g1468 ( 
.A(n_1398),
.B(n_1341),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1337),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1334),
.B(n_1343),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1424),
.B(n_1342),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1420),
.Y(n_1472)
);

OA21x2_ASAP7_75t_L g1473 ( 
.A1(n_1409),
.A2(n_1386),
.B(n_1389),
.Y(n_1473)
);

AO21x1_ASAP7_75t_SL g1474 ( 
.A1(n_1350),
.A2(n_1342),
.B(n_1353),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1410),
.A2(n_1389),
.B(n_1411),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1344),
.B(n_1362),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1399),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1360),
.A2(n_1345),
.B1(n_1437),
.B2(n_1461),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1426),
.B(n_1460),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_1369),
.Y(n_1480)
);

AO21x2_ASAP7_75t_L g1481 ( 
.A1(n_1400),
.A2(n_1368),
.B(n_1402),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1404),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1339),
.B(n_1434),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1392),
.Y(n_1484)
);

AO21x2_ASAP7_75t_L g1485 ( 
.A1(n_1368),
.A2(n_1437),
.B(n_1359),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1418),
.A2(n_1362),
.B(n_1421),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1346),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1421),
.B(n_1419),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1332),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1332),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1373),
.B(n_1425),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1418),
.A2(n_1353),
.B(n_1364),
.Y(n_1492)
);

INVxp67_ASAP7_75t_L g1493 ( 
.A(n_1450),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1350),
.B(n_1414),
.Y(n_1494)
);

INVxp33_ASAP7_75t_SL g1495 ( 
.A(n_1429),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1354),
.Y(n_1496)
);

OAI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1372),
.A2(n_1338),
.B(n_1445),
.Y(n_1497)
);

AO31x2_ASAP7_75t_L g1498 ( 
.A1(n_1422),
.A2(n_1423),
.A3(n_1333),
.B(n_1417),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1357),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1361),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1363),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1369),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1367),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1431),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1440),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1447),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1338),
.B(n_1393),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1380),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1339),
.B(n_1434),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1405),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1458),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1416),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1415),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1415),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1364),
.B(n_1356),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1369),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1375),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1365),
.B(n_1359),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1336),
.Y(n_1519)
);

OR2x6_ASAP7_75t_L g1520 ( 
.A(n_1378),
.B(n_1394),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1371),
.B(n_1351),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1366),
.Y(n_1522)
);

BUFx4f_ASAP7_75t_SL g1523 ( 
.A(n_1352),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1412),
.Y(n_1524)
);

AOI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1430),
.A2(n_1445),
.B1(n_1435),
.B2(n_1455),
.C(n_1456),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1463),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1454),
.B(n_1365),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1403),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1355),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1358),
.B(n_1395),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1408),
.Y(n_1531)
);

NOR2x1_ASAP7_75t_R g1532 ( 
.A(n_1428),
.B(n_1452),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1413),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1358),
.B(n_1456),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1442),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1442),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1438),
.A2(n_1444),
.B1(n_1455),
.B2(n_1340),
.Y(n_1537)
);

OR2x6_ASAP7_75t_L g1538 ( 
.A(n_1394),
.B(n_1384),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1377),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1376),
.B(n_1459),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1391),
.B(n_1396),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1453),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1453),
.Y(n_1543)
);

AND2x6_ASAP7_75t_L g1544 ( 
.A(n_1453),
.B(n_1382),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1457),
.B(n_1349),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1385),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1370),
.B(n_1385),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1390),
.B(n_1462),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1407),
.B(n_1387),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1405),
.Y(n_1550)
);

A2O1A1Ixp33_ASAP7_75t_L g1551 ( 
.A1(n_1381),
.A2(n_1401),
.B(n_1448),
.C(n_1443),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1448),
.B(n_1379),
.Y(n_1552)
);

BUFx2_ASAP7_75t_R g1553 ( 
.A(n_1441),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1374),
.B(n_1443),
.Y(n_1554)
);

AOI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1466),
.A2(n_1347),
.B1(n_1432),
.B2(n_1446),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1468),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1529),
.B(n_1433),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1483),
.B(n_1383),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_R g1559 ( 
.A(n_1519),
.B(n_1436),
.Y(n_1559)
);

BUFx8_ASAP7_75t_L g1560 ( 
.A(n_1510),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_SL g1561 ( 
.A1(n_1497),
.A2(n_1347),
.B(n_1439),
.Y(n_1561)
);

OAI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1478),
.A2(n_1451),
.B(n_1381),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1488),
.B(n_1348),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1529),
.B(n_1526),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_SL g1565 ( 
.A1(n_1515),
.A2(n_1509),
.B1(n_1471),
.B2(n_1494),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1499),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1472),
.B(n_1470),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1525),
.A2(n_1537),
.B(n_1479),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1469),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1507),
.B(n_1535),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1534),
.A2(n_1518),
.B1(n_1512),
.B2(n_1471),
.Y(n_1571)
);

OAI211xp5_ASAP7_75t_L g1572 ( 
.A1(n_1534),
.A2(n_1535),
.B(n_1536),
.C(n_1518),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1511),
.B(n_1498),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1520),
.B(n_1476),
.Y(n_1574)
);

NOR2xp67_ASAP7_75t_L g1575 ( 
.A(n_1513),
.B(n_1514),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1498),
.B(n_1496),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1508),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1536),
.B(n_1517),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1541),
.B(n_1512),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1541),
.B(n_1494),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1527),
.B(n_1470),
.Y(n_1581)
);

NOR2x1_ASAP7_75t_SL g1582 ( 
.A(n_1520),
.B(n_1485),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1498),
.B(n_1500),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1498),
.B(n_1500),
.Y(n_1584)
);

NOR2x1_ASAP7_75t_SL g1585 ( 
.A(n_1520),
.B(n_1485),
.Y(n_1585)
);

INVx3_ASAP7_75t_L g1586 ( 
.A(n_1470),
.Y(n_1586)
);

A2O1A1Ixp33_ASAP7_75t_L g1587 ( 
.A1(n_1515),
.A2(n_1530),
.B(n_1531),
.C(n_1528),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1532),
.A2(n_1551),
.B(n_1520),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1498),
.B(n_1501),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1487),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1530),
.A2(n_1548),
.B1(n_1553),
.B2(n_1493),
.Y(n_1591)
);

INVx4_ASAP7_75t_L g1592 ( 
.A(n_1520),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1503),
.A2(n_1485),
.B1(n_1491),
.B2(n_1528),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1522),
.Y(n_1594)
);

A2O1A1Ixp33_ASAP7_75t_L g1595 ( 
.A1(n_1531),
.A2(n_1491),
.B(n_1486),
.C(n_1474),
.Y(n_1595)
);

OAI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1475),
.A2(n_1467),
.B(n_1513),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1498),
.B(n_1504),
.Y(n_1597)
);

AOI21xp33_ASAP7_75t_L g1598 ( 
.A1(n_1481),
.A2(n_1514),
.B(n_1464),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1505),
.B(n_1506),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1524),
.A2(n_1550),
.B1(n_1510),
.B2(n_1552),
.Y(n_1600)
);

NOR2x1_ASAP7_75t_SL g1601 ( 
.A(n_1481),
.B(n_1538),
.Y(n_1601)
);

AO32x2_ASAP7_75t_L g1602 ( 
.A1(n_1480),
.A2(n_1516),
.A3(n_1502),
.B1(n_1489),
.B2(n_1490),
.Y(n_1602)
);

NAND4xp25_ASAP7_75t_L g1603 ( 
.A(n_1484),
.B(n_1506),
.C(n_1540),
.D(n_1521),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1524),
.A2(n_1550),
.B1(n_1510),
.B2(n_1545),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1464),
.A2(n_1465),
.B(n_1481),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1477),
.Y(n_1606)
);

INVxp67_ASAP7_75t_L g1607 ( 
.A(n_1547),
.Y(n_1607)
);

AOI221x1_ASAP7_75t_L g1608 ( 
.A1(n_1533),
.A2(n_1543),
.B1(n_1539),
.B2(n_1542),
.C(n_1546),
.Y(n_1608)
);

NAND2x1_ASAP7_75t_L g1609 ( 
.A(n_1544),
.B(n_1538),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1549),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1594),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1573),
.B(n_1464),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1573),
.B(n_1473),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1566),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1586),
.B(n_1475),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1586),
.B(n_1482),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1576),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1606),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1576),
.B(n_1473),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1564),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1568),
.A2(n_1474),
.B1(n_1492),
.B2(n_1491),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1583),
.B(n_1473),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1567),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1602),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1584),
.B(n_1486),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1558),
.B(n_1587),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1587),
.A2(n_1492),
.B1(n_1491),
.B2(n_1550),
.Y(n_1627)
);

AND2x4_ASAP7_75t_SL g1628 ( 
.A(n_1592),
.B(n_1472),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1599),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1589),
.B(n_1597),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1597),
.B(n_1596),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1555),
.A2(n_1565),
.B1(n_1591),
.B2(n_1558),
.Y(n_1632)
);

NOR2x1p5_ASAP7_75t_L g1633 ( 
.A(n_1609),
.B(n_1550),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1617),
.B(n_1577),
.Y(n_1634)
);

AOI221xp5_ASAP7_75t_L g1635 ( 
.A1(n_1626),
.A2(n_1571),
.B1(n_1572),
.B2(n_1578),
.C(n_1598),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1614),
.Y(n_1636)
);

AOI33xp33_ASAP7_75t_L g1637 ( 
.A1(n_1621),
.A2(n_1593),
.A3(n_1563),
.B1(n_1579),
.B2(n_1580),
.B3(n_1610),
.Y(n_1637)
);

NAND4xp25_ASAP7_75t_L g1638 ( 
.A(n_1632),
.B(n_1562),
.C(n_1578),
.D(n_1595),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1614),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1625),
.B(n_1630),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1625),
.B(n_1582),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1620),
.B(n_1611),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1633),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1629),
.Y(n_1644)
);

BUFx3_ASAP7_75t_L g1645 ( 
.A(n_1628),
.Y(n_1645)
);

NAND4xp25_ASAP7_75t_SL g1646 ( 
.A(n_1632),
.B(n_1588),
.C(n_1595),
.D(n_1563),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1629),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1620),
.B(n_1570),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1633),
.B(n_1601),
.Y(n_1649)
);

OR2x6_ASAP7_75t_L g1650 ( 
.A(n_1633),
.B(n_1574),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_R g1651 ( 
.A(n_1626),
.B(n_1556),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1615),
.B(n_1616),
.Y(n_1652)
);

BUFx2_ASAP7_75t_L g1653 ( 
.A(n_1623),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1611),
.Y(n_1654)
);

AOI221xp5_ASAP7_75t_L g1655 ( 
.A1(n_1627),
.A2(n_1569),
.B1(n_1603),
.B2(n_1605),
.C(n_1590),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1618),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1625),
.B(n_1585),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1630),
.B(n_1613),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1618),
.Y(n_1659)
);

INVxp67_ASAP7_75t_SL g1660 ( 
.A(n_1617),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1629),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1613),
.B(n_1581),
.Y(n_1662)
);

NAND3xp33_ASAP7_75t_L g1663 ( 
.A(n_1621),
.B(n_1607),
.C(n_1608),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1639),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1644),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1644),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1644),
.B(n_1624),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1647),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1640),
.B(n_1624),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1640),
.B(n_1624),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1645),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1647),
.B(n_1619),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1653),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1640),
.B(n_1631),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1658),
.B(n_1631),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1658),
.B(n_1631),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1639),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1656),
.B(n_1659),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1636),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1661),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1663),
.A2(n_1575),
.B(n_1612),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1652),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1661),
.Y(n_1683)
);

INVx4_ASAP7_75t_L g1684 ( 
.A(n_1650),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1636),
.Y(n_1685)
);

INVx4_ASAP7_75t_L g1686 ( 
.A(n_1650),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1641),
.B(n_1622),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1661),
.B(n_1622),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1641),
.B(n_1612),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1646),
.A2(n_1492),
.B1(n_1561),
.B2(n_1612),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1674),
.B(n_1643),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1681),
.A2(n_1646),
.B(n_1655),
.Y(n_1692)
);

INVx2_ASAP7_75t_SL g1693 ( 
.A(n_1671),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1681),
.B(n_1667),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1667),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1671),
.B(n_1643),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_SL g1697 ( 
.A(n_1690),
.B(n_1651),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1674),
.B(n_1643),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1674),
.B(n_1657),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1684),
.B(n_1532),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1673),
.Y(n_1701)
);

O2A1O1Ixp5_ASAP7_75t_SL g1702 ( 
.A1(n_1681),
.A2(n_1664),
.B(n_1677),
.C(n_1679),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1678),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1667),
.B(n_1634),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1675),
.B(n_1637),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1667),
.B(n_1634),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1678),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1672),
.B(n_1642),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1678),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1673),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1671),
.Y(n_1711)
);

OR2x6_ASAP7_75t_L g1712 ( 
.A(n_1684),
.B(n_1650),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1675),
.B(n_1635),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1671),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1675),
.B(n_1635),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1664),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1672),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1664),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1675),
.B(n_1662),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1676),
.B(n_1662),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1676),
.B(n_1662),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1671),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1677),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1677),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1672),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1674),
.B(n_1676),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1673),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1685),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1676),
.B(n_1648),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1685),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1685),
.Y(n_1731)
);

NAND3xp33_ASAP7_75t_L g1732 ( 
.A(n_1690),
.B(n_1655),
.C(n_1663),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1672),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1713),
.B(n_1689),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1705),
.B(n_1688),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1732),
.A2(n_1692),
.B1(n_1638),
.B2(n_1697),
.Y(n_1736)
);

OAI221xp5_ASAP7_75t_SL g1737 ( 
.A1(n_1715),
.A2(n_1690),
.B1(n_1638),
.B2(n_1650),
.C(n_1657),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1722),
.B(n_1689),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1714),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1716),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1716),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1723),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1726),
.B(n_1684),
.Y(n_1743)
);

INVx1_ASAP7_75t_SL g1744 ( 
.A(n_1714),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1693),
.B(n_1689),
.Y(n_1745)
);

INVx2_ASAP7_75t_SL g1746 ( 
.A(n_1696),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1693),
.B(n_1689),
.Y(n_1747)
);

OR2x6_ASAP7_75t_L g1748 ( 
.A(n_1711),
.B(n_1684),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1729),
.B(n_1688),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1723),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1726),
.B(n_1684),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1691),
.B(n_1684),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1695),
.Y(n_1753)
);

NAND2x1_ASAP7_75t_L g1754 ( 
.A(n_1696),
.B(n_1684),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1691),
.B(n_1686),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1698),
.B(n_1686),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1695),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1711),
.B(n_1687),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1718),
.Y(n_1759)
);

OA21x2_ASAP7_75t_L g1760 ( 
.A1(n_1728),
.A2(n_1666),
.B(n_1665),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1700),
.B(n_1495),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1724),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1701),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1717),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1710),
.Y(n_1765)
);

INVx1_ASAP7_75t_SL g1766 ( 
.A(n_1696),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1698),
.B(n_1712),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1727),
.B(n_1687),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1728),
.Y(n_1769)
);

O2A1O1Ixp33_ASAP7_75t_L g1770 ( 
.A1(n_1737),
.A2(n_1694),
.B(n_1702),
.C(n_1712),
.Y(n_1770)
);

INVxp67_ASAP7_75t_L g1771 ( 
.A(n_1765),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_SL g1772 ( 
.A1(n_1736),
.A2(n_1694),
.B(n_1600),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1736),
.A2(n_1712),
.B1(n_1686),
.B2(n_1650),
.Y(n_1773)
);

AOI21xp33_ASAP7_75t_L g1774 ( 
.A1(n_1754),
.A2(n_1712),
.B(n_1686),
.Y(n_1774)
);

NOR3xp33_ASAP7_75t_L g1775 ( 
.A(n_1763),
.B(n_1686),
.C(n_1557),
.Y(n_1775)
);

NAND3xp33_ASAP7_75t_L g1776 ( 
.A(n_1763),
.B(n_1702),
.C(n_1686),
.Y(n_1776)
);

NAND4xp75_ASAP7_75t_SL g1777 ( 
.A(n_1767),
.B(n_1699),
.C(n_1670),
.D(n_1669),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1739),
.B(n_1699),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1734),
.A2(n_1686),
.B1(n_1533),
.B2(n_1709),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1766),
.B(n_1719),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1754),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1767),
.B(n_1687),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1752),
.B(n_1687),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1740),
.Y(n_1784)
);

OAI221xp5_ASAP7_75t_L g1785 ( 
.A1(n_1746),
.A2(n_1706),
.B1(n_1704),
.B2(n_1708),
.C(n_1721),
.Y(n_1785)
);

A2O1A1Ixp33_ASAP7_75t_L g1786 ( 
.A1(n_1761),
.A2(n_1556),
.B(n_1660),
.C(n_1549),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1752),
.A2(n_1649),
.B1(n_1650),
.B2(n_1604),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1740),
.Y(n_1788)
);

OAI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1746),
.A2(n_1707),
.B(n_1703),
.Y(n_1789)
);

AOI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1744),
.A2(n_1709),
.B1(n_1703),
.B2(n_1707),
.C(n_1733),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1741),
.Y(n_1791)
);

OAI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1735),
.A2(n_1660),
.B1(n_1592),
.B2(n_1720),
.Y(n_1792)
);

OAI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1735),
.A2(n_1592),
.B1(n_1645),
.B2(n_1708),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1744),
.B(n_1704),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1741),
.Y(n_1795)
);

OAI21xp33_ASAP7_75t_SL g1796 ( 
.A1(n_1777),
.A2(n_1748),
.B(n_1755),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1782),
.B(n_1755),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1784),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1771),
.B(n_1768),
.Y(n_1799)
);

AOI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1770),
.A2(n_1769),
.B1(n_1756),
.B2(n_1743),
.C(n_1751),
.Y(n_1800)
);

NAND3xp33_ASAP7_75t_SL g1801 ( 
.A(n_1772),
.B(n_1559),
.C(n_1769),
.Y(n_1801)
);

BUFx2_ASAP7_75t_L g1802 ( 
.A(n_1781),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1794),
.B(n_1738),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1788),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1779),
.B(n_1775),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1780),
.B(n_1745),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1778),
.B(n_1747),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1791),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1785),
.B(n_1758),
.Y(n_1809)
);

O2A1O1Ixp33_ASAP7_75t_L g1810 ( 
.A1(n_1776),
.A2(n_1762),
.B(n_1759),
.C(n_1748),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1779),
.B(n_1756),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1790),
.B(n_1743),
.Y(n_1812)
);

INVx1_ASAP7_75t_SL g1813 ( 
.A(n_1774),
.Y(n_1813)
);

NAND2xp33_ASAP7_75t_L g1814 ( 
.A(n_1786),
.B(n_1559),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1795),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1802),
.B(n_1813),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1798),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1804),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1805),
.A2(n_1786),
.B1(n_1789),
.B2(n_1787),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1808),
.Y(n_1820)
);

AOI21xp33_ASAP7_75t_L g1821 ( 
.A1(n_1810),
.A2(n_1773),
.B(n_1792),
.Y(n_1821)
);

AOI211x1_ASAP7_75t_L g1822 ( 
.A1(n_1801),
.A2(n_1792),
.B(n_1793),
.C(n_1751),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1815),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1799),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1800),
.B(n_1783),
.Y(n_1825)
);

XOR2x2_ASAP7_75t_L g1826 ( 
.A(n_1801),
.B(n_1549),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1797),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1827),
.Y(n_1828)
);

O2A1O1Ixp33_ASAP7_75t_SL g1829 ( 
.A1(n_1821),
.A2(n_1810),
.B(n_1812),
.C(n_1811),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1816),
.Y(n_1830)
);

NOR2xp67_ASAP7_75t_L g1831 ( 
.A(n_1817),
.B(n_1796),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1825),
.B(n_1803),
.Y(n_1832)
);

NOR2x1_ASAP7_75t_L g1833 ( 
.A(n_1818),
.B(n_1814),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1824),
.B(n_1809),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1822),
.A2(n_1807),
.B1(n_1806),
.B2(n_1748),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1819),
.B(n_1814),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1819),
.B(n_1793),
.Y(n_1837)
);

NAND3xp33_ASAP7_75t_SL g1838 ( 
.A(n_1820),
.B(n_1757),
.C(n_1753),
.Y(n_1838)
);

AOI222xp33_ASAP7_75t_L g1839 ( 
.A1(n_1832),
.A2(n_1823),
.B1(n_1826),
.B2(n_1821),
.C1(n_1759),
.C2(n_1762),
.Y(n_1839)
);

AOI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1829),
.A2(n_1757),
.B1(n_1753),
.B2(n_1764),
.C(n_1742),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1833),
.B(n_1748),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_L g1842 ( 
.A(n_1836),
.B(n_1748),
.C(n_1753),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1828),
.Y(n_1843)
);

O2A1O1Ixp33_ASAP7_75t_L g1844 ( 
.A1(n_1839),
.A2(n_1837),
.B(n_1834),
.C(n_1830),
.Y(n_1844)
);

AOI221xp5_ASAP7_75t_L g1845 ( 
.A1(n_1842),
.A2(n_1835),
.B1(n_1838),
.B2(n_1757),
.C(n_1831),
.Y(n_1845)
);

OAI222xp33_ASAP7_75t_L g1846 ( 
.A1(n_1841),
.A2(n_1843),
.B1(n_1764),
.B2(n_1750),
.C1(n_1742),
.C2(n_1749),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1840),
.A2(n_1764),
.B1(n_1750),
.B2(n_1730),
.C(n_1731),
.Y(n_1847)
);

AOI211xp5_ASAP7_75t_SL g1848 ( 
.A1(n_1843),
.A2(n_1523),
.B(n_1730),
.C(n_1731),
.Y(n_1848)
);

NOR2x1_ASAP7_75t_L g1849 ( 
.A(n_1842),
.B(n_1760),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1845),
.A2(n_1560),
.B1(n_1549),
.B2(n_1733),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1849),
.Y(n_1851)
);

NAND2xp33_ASAP7_75t_L g1852 ( 
.A(n_1847),
.B(n_1706),
.Y(n_1852)
);

OAI211xp5_ASAP7_75t_L g1853 ( 
.A1(n_1844),
.A2(n_1760),
.B(n_1749),
.C(n_1725),
.Y(n_1853)
);

OAI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1848),
.A2(n_1717),
.B1(n_1725),
.B2(n_1524),
.C(n_1760),
.Y(n_1854)
);

AOI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1853),
.A2(n_1846),
.B1(n_1642),
.B2(n_1654),
.C(n_1682),
.Y(n_1855)
);

OAI211xp5_ASAP7_75t_SL g1856 ( 
.A1(n_1850),
.A2(n_1524),
.B(n_1560),
.C(n_1682),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1851),
.B(n_1682),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1857),
.B(n_1854),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1858),
.A2(n_1856),
.B1(n_1852),
.B2(n_1855),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1859),
.Y(n_1860)
);

NOR3xp33_ASAP7_75t_L g1861 ( 
.A(n_1859),
.B(n_1560),
.C(n_1554),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1860),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1861),
.Y(n_1863)
);

OAI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1862),
.A2(n_1760),
.B1(n_1682),
.B2(n_1683),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1863),
.Y(n_1865)
);

OA21x2_ASAP7_75t_L g1866 ( 
.A1(n_1865),
.A2(n_1666),
.B(n_1665),
.Y(n_1866)
);

OAI21xp5_ASAP7_75t_SL g1867 ( 
.A1(n_1866),
.A2(n_1864),
.B(n_1554),
.Y(n_1867)
);

CKINVDCx20_ASAP7_75t_R g1868 ( 
.A(n_1867),
.Y(n_1868)
);

AOI221xp5_ASAP7_75t_L g1869 ( 
.A1(n_1868),
.A2(n_1683),
.B1(n_1680),
.B2(n_1668),
.C(n_1665),
.Y(n_1869)
);

AOI211xp5_ASAP7_75t_L g1870 ( 
.A1(n_1869),
.A2(n_1480),
.B(n_1516),
.C(n_1502),
.Y(n_1870)
);


endmodule