module fake_ibex_768_n_1353 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_247, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_8, n_118, n_224, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_256, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_14, n_0, n_239, n_94, n_134, n_12, n_42, n_77, n_112, n_257, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_258, n_80, n_172, n_215, n_250, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_259, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1353);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_247;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_8;
input n_118;
input n_224;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_256;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_257;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_258;
input n_80;
input n_172;
input n_215;
input n_250;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_259;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1353;

wire n_1084;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_280;
wire n_375;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_573;
wire n_359;
wire n_262;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_397;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1108;
wire n_382;
wire n_1239;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_1281;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_282;
wire n_870;
wire n_1298;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_737;
wire n_606;
wire n_462;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_657;
wire n_1156;
wire n_1293;
wire n_749;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1015;
wire n_663;
wire n_1152;
wire n_371;
wire n_1036;
wire n_974;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_840;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_413;
wire n_1069;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_998;
wire n_1115;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_291;
wire n_318;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_997;
wire n_891;
wire n_303;
wire n_717;
wire n_668;
wire n_871;
wire n_266;
wire n_1339;
wire n_485;
wire n_1315;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1048;
wire n_774;
wire n_588;
wire n_1251;
wire n_1247;
wire n_528;
wire n_260;
wire n_836;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_423;
wire n_357;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1291;
wire n_317;
wire n_326;
wire n_270;
wire n_1340;
wire n_276;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_1112;
wire n_1267;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_804;
wire n_484;
wire n_480;
wire n_354;
wire n_1057;
wire n_516;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_277;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1221;
wire n_284;
wire n_1047;
wire n_792;
wire n_1314;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_478;
wire n_336;
wire n_861;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1098;
wire n_584;
wire n_1187;
wire n_698;
wire n_1061;
wire n_682;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_265;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1023;
wire n_568;
wire n_813;
wire n_1211;
wire n_1284;
wire n_1116;
wire n_791;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1074;
wire n_759;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_263;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_735;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1033;
wire n_627;
wire n_990;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_264;
wire n_1145;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1277;
wire n_1016;
wire n_680;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_271;
wire n_984;
wire n_394;
wire n_364;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_137),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_34),
.Y(n_261)
);

BUFx2_ASAP7_75t_SL g262 ( 
.A(n_124),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_112),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_L g264 ( 
.A(n_25),
.B(n_252),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_3),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_91),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_175),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_194),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_118),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_30),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_64),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_186),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_188),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_107),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_250),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_218),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_79),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_102),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_162),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_18),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_203),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_7),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_192),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_184),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_145),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_133),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_87),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_73),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_249),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_138),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_254),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_22),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_168),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_245),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_131),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_2),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_216),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_8),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_209),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_211),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_146),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_94),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_38),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_155),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_46),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_244),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_79),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_251),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_7),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_24),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_117),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_191),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_176),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_222),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_182),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_5),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_243),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_253),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_29),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_148),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_10),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_72),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_246),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_60),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_152),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_167),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_129),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_190),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_165),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_157),
.Y(n_330)
);

BUFx2_ASAP7_75t_SL g331 ( 
.A(n_185),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_159),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_220),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_95),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_230),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_196),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_44),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_49),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_67),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_151),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_213),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_147),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_144),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_240),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_227),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_8),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_180),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_241),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_257),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_174),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_31),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_30),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_14),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_46),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_228),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_189),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_67),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_52),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_173),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_116),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_89),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_68),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_74),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_224),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_161),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_120),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g367 ( 
.A(n_166),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_210),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_22),
.B(n_199),
.Y(n_369)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_248),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_135),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_141),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_127),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_92),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_181),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_238),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_223),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_247),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_27),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_206),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_51),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_78),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_150),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_221),
.B(n_164),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_71),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_156),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_76),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_202),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_69),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_12),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_178),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_98),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_1),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_77),
.Y(n_394)
);

BUFx5_ASAP7_75t_L g395 ( 
.A(n_187),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g396 ( 
.A(n_139),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_128),
.B(n_105),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_134),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_16),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_255),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_235),
.Y(n_401)
);

BUFx2_ASAP7_75t_SL g402 ( 
.A(n_4),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_231),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_234),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_83),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_226),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_86),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_236),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_197),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_179),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_59),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_132),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_170),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_36),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_130),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_177),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_61),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_29),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_55),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_102),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_64),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_163),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_110),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_193),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_69),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_15),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_94),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_126),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_72),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_237),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_62),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_225),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_54),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_258),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_12),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_42),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_3),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_229),
.Y(n_438)
);

INVxp33_ASAP7_75t_L g439 ( 
.A(n_172),
.Y(n_439)
);

NOR2xp67_ASAP7_75t_L g440 ( 
.A(n_62),
.B(n_54),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_233),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_198),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_239),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_0),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_160),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_61),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_195),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_53),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_158),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_65),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_11),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_279),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_429),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_429),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_315),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_309),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_265),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_370),
.Y(n_459)
);

OA21x2_ASAP7_75t_L g460 ( 
.A1(n_293),
.A2(n_333),
.B(n_330),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_370),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_411),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_265),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_411),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_286),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_315),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_315),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_358),
.B(n_1),
.Y(n_468)
);

OAI21x1_ASAP7_75t_L g469 ( 
.A1(n_293),
.A2(n_111),
.B(n_109),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_334),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_358),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_263),
.B(n_2),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_274),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_334),
.Y(n_474)
);

OAI22x1_ASAP7_75t_R g475 ( 
.A1(n_302),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_399),
.Y(n_476)
);

AND2x2_ASAP7_75t_SL g477 ( 
.A(n_428),
.B(n_113),
.Y(n_477)
);

BUFx8_ASAP7_75t_L g478 ( 
.A(n_263),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_279),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_370),
.Y(n_480)
);

CKINVDCx6p67_ASAP7_75t_R g481 ( 
.A(n_286),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_421),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_370),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_421),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_298),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_446),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_302),
.A2(n_337),
.B1(n_346),
.B2(n_303),
.Y(n_487)
);

INVx5_ASAP7_75t_L g488 ( 
.A(n_286),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_370),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_399),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_303),
.A2(n_337),
.B1(n_420),
.B2(n_346),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_446),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g493 ( 
.A1(n_330),
.A2(n_115),
.B(n_114),
.Y(n_493)
);

INVx5_ASAP7_75t_L g494 ( 
.A(n_289),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_305),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_495)
);

OAI22x1_ASAP7_75t_R g496 ( 
.A1(n_420),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_289),
.B(n_17),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_360),
.B(n_19),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_273),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_267),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_370),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_304),
.Y(n_502)
);

BUFx8_ASAP7_75t_L g503 ( 
.A(n_367),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_439),
.B(n_19),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_370),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_268),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_395),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_361),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_508)
);

OA21x2_ASAP7_75t_L g509 ( 
.A1(n_333),
.A2(n_121),
.B(n_119),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_269),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_367),
.B(n_20),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_271),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_273),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_304),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_396),
.B(n_21),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_395),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_395),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_313),
.Y(n_518)
);

BUFx8_ASAP7_75t_L g519 ( 
.A(n_396),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_426),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_520)
);

AND2x6_ASAP7_75t_L g521 ( 
.A(n_313),
.B(n_122),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_274),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_522)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_412),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_281),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_395),
.Y(n_525)
);

CKINVDCx11_ASAP7_75t_R g526 ( 
.A(n_426),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_413),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_284),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_413),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_422),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_395),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_422),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_291),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_395),
.Y(n_534)
);

OA21x2_ASAP7_75t_L g535 ( 
.A1(n_345),
.A2(n_125),
.B(n_123),
.Y(n_535)
);

INVx5_ASAP7_75t_L g536 ( 
.A(n_438),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_294),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_438),
.B(n_28),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_261),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_345),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_277),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_297),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_299),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_459),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_465),
.B(n_439),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_465),
.B(n_277),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_540),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_540),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_488),
.B(n_340),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_511),
.Y(n_550)
);

NAND3xp33_ASAP7_75t_L g551 ( 
.A(n_504),
.B(n_282),
.C(n_278),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_468),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_488),
.B(n_260),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_462),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_481),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_462),
.B(n_278),
.Y(n_556)
);

BUFx6f_ASAP7_75t_SL g557 ( 
.A(n_477),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_460),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_460),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_468),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_460),
.Y(n_561)
);

INVxp67_ASAP7_75t_SL g562 ( 
.A(n_464),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_473),
.B(n_357),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_504),
.A2(n_270),
.B1(n_280),
.B2(n_266),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_481),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_477),
.A2(n_448),
.B1(n_451),
.B2(n_357),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_479),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_459),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_541),
.B(n_448),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_490),
.B(n_432),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_461),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_453),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_480),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_491),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_453),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_476),
.Y(n_576)
);

AND2x4_ASAP7_75t_SL g577 ( 
.A(n_485),
.B(n_276),
.Y(n_577)
);

INVxp33_ASAP7_75t_L g578 ( 
.A(n_476),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_453),
.B(n_451),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_502),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_454),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_500),
.B(n_506),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_458),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_458),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_526),
.Y(n_585)
);

AND3x1_ASAP7_75t_L g586 ( 
.A(n_508),
.B(n_450),
.C(n_288),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_478),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_458),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g589 ( 
.A(n_472),
.B(n_296),
.C(n_292),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_502),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_454),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_455),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_478),
.B(n_275),
.Y(n_593)
);

NOR2x1p5_ASAP7_75t_L g594 ( 
.A(n_499),
.B(n_287),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_503),
.B(n_519),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_455),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_503),
.B(n_275),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_503),
.B(n_519),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_518),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_518),
.Y(n_600)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_499),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_519),
.B(n_500),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_513),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_518),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_456),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_527),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_463),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_527),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_527),
.Y(n_609)
);

INVx11_ASAP7_75t_L g610 ( 
.A(n_521),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_521),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_506),
.B(n_301),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_510),
.B(n_283),
.Y(n_613)
);

OAI22xp33_ASAP7_75t_L g614 ( 
.A1(n_522),
.A2(n_444),
.B1(n_400),
.B2(n_416),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_471),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_452),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_452),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_L g618 ( 
.A(n_521),
.B(n_395),
.Y(n_618)
);

BUFx10_ASAP7_75t_L g619 ( 
.A(n_497),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_471),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_487),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_527),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_539),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_530),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_530),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_457),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_524),
.B(n_285),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_513),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_528),
.B(n_285),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_530),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_457),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_470),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_530),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_514),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_529),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_529),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_533),
.B(n_290),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_532),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_474),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_SL g640 ( 
.A(n_498),
.B(n_314),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_532),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_532),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_482),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_482),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_537),
.B(n_542),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_542),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_543),
.B(n_442),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_543),
.B(n_443),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_484),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_494),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_494),
.B(n_523),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_475),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_492),
.B(n_443),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_515),
.A2(n_400),
.B1(n_416),
.B2(n_314),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_532),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_483),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_494),
.B(n_523),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_520),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_532),
.Y(n_659)
);

OR2x6_ASAP7_75t_L g660 ( 
.A(n_495),
.B(n_402),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_489),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_521),
.A2(n_319),
.B1(n_321),
.B2(n_310),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_501),
.Y(n_663)
);

BUFx10_ASAP7_75t_L g664 ( 
.A(n_521),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_501),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_L g666 ( 
.A(n_505),
.B(n_449),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_505),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_507),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_507),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_492),
.B(n_440),
.Y(n_670)
);

AOI21x1_ASAP7_75t_L g671 ( 
.A1(n_516),
.A2(n_410),
.B(n_312),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_492),
.B(n_392),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_646),
.B(n_516),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_653),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_579),
.A2(n_538),
.B1(n_525),
.B2(n_531),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_645),
.B(n_517),
.Y(n_676)
);

INVx8_ASAP7_75t_L g677 ( 
.A(n_555),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_554),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_645),
.B(n_517),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_579),
.B(n_525),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_572),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_572),
.Y(n_682)
);

NOR2x1p5_ASAP7_75t_L g683 ( 
.A(n_555),
.B(n_496),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_582),
.B(n_531),
.Y(n_684)
);

AOI221xp5_ASAP7_75t_L g685 ( 
.A1(n_586),
.A2(n_614),
.B1(n_640),
.B2(n_564),
.C(n_578),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_545),
.B(n_534),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_575),
.Y(n_687)
);

OAI22xp33_ASAP7_75t_L g688 ( 
.A1(n_566),
.A2(n_444),
.B1(n_316),
.B2(n_322),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_623),
.B(n_534),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_583),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_583),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_552),
.A2(n_352),
.B1(n_353),
.B2(n_338),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_584),
.Y(n_693)
);

OAI22xp5_ASAP7_75t_L g694 ( 
.A1(n_658),
.A2(n_384),
.B1(n_390),
.B2(n_389),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_587),
.B(n_536),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_546),
.B(n_578),
.Y(n_696)
);

OAI22xp33_ASAP7_75t_L g697 ( 
.A1(n_660),
.A2(n_339),
.B1(n_351),
.B2(n_307),
.Y(n_697)
);

OR2x6_ASAP7_75t_L g698 ( 
.A(n_660),
.B(n_262),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_584),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_576),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_560),
.A2(n_407),
.B1(n_414),
.B2(n_405),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_588),
.Y(n_702)
);

NAND2x1p5_ASAP7_75t_L g703 ( 
.A(n_595),
.B(n_418),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_607),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_607),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_648),
.B(n_486),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_556),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_565),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_556),
.B(n_272),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_570),
.B(n_300),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_611),
.B(n_306),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_562),
.B(n_388),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_664),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_551),
.B(n_469),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_662),
.B(n_308),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_563),
.B(n_354),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_615),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_613),
.B(n_318),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_602),
.B(n_406),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_589),
.B(n_415),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_598),
.B(n_326),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_672),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_557),
.A2(n_363),
.B1(n_374),
.B2(n_362),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_654),
.A2(n_379),
.B1(n_385),
.B2(n_382),
.Y(n_724)
);

NAND2xp33_ASAP7_75t_L g725 ( 
.A(n_550),
.B(n_327),
.Y(n_725)
);

INVx8_ASAP7_75t_L g726 ( 
.A(n_565),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_619),
.B(n_328),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_581),
.B(n_493),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_635),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_591),
.B(n_295),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_619),
.B(n_332),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_619),
.B(n_336),
.Y(n_732)
);

BUFx6f_ASAP7_75t_SL g733 ( 
.A(n_660),
.Y(n_733)
);

INVx8_ASAP7_75t_L g734 ( 
.A(n_557),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_627),
.B(n_341),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_620),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_592),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_596),
.B(n_403),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_664),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_557),
.A2(n_271),
.B1(n_381),
.B2(n_324),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_636),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_569),
.B(n_434),
.Y(n_742)
);

INVxp33_ASAP7_75t_L g743 ( 
.A(n_569),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_544),
.B(n_509),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_672),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_544),
.B(n_509),
.Y(n_746)
);

A2O1A1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_612),
.A2(n_311),
.B(n_320),
.C(n_317),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_629),
.B(n_348),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_626),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_593),
.B(n_350),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_594),
.B(n_264),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_597),
.B(n_356),
.Y(n_752)
);

OAI22xp33_ASAP7_75t_L g753 ( 
.A1(n_660),
.A2(n_393),
.B1(n_394),
.B2(n_387),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_631),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_637),
.B(n_647),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_666),
.B(n_365),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_616),
.B(n_372),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_616),
.B(n_373),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_617),
.B(n_380),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_634),
.B(n_391),
.Y(n_760)
);

OR2x6_ASAP7_75t_L g761 ( 
.A(n_621),
.B(n_331),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_634),
.B(n_398),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_632),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_640),
.A2(n_419),
.B1(n_425),
.B2(n_417),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_639),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_549),
.B(n_408),
.Y(n_766)
);

NOR3xp33_ASAP7_75t_L g767 ( 
.A(n_603),
.B(n_431),
.C(n_427),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_618),
.A2(n_435),
.B1(n_436),
.B2(n_433),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_643),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_670),
.B(n_437),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_553),
.B(n_409),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_558),
.A2(n_325),
.B(n_329),
.C(n_323),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_644),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_649),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_559),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_568),
.B(n_509),
.Y(n_776)
);

OR2x6_ASAP7_75t_L g777 ( 
.A(n_670),
.B(n_369),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_561),
.Y(n_778)
);

NAND2xp33_ASAP7_75t_SL g779 ( 
.A(n_628),
.B(n_652),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_661),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_661),
.B(n_423),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_671),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_571),
.B(n_335),
.Y(n_783)
);

O2A1O1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_618),
.A2(n_342),
.B(n_344),
.C(n_343),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_665),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_573),
.B(n_347),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_573),
.B(n_349),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_656),
.B(n_355),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_656),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_663),
.B(n_667),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_663),
.B(n_667),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_668),
.B(n_535),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_668),
.B(n_535),
.Y(n_793)
);

NOR3xp33_ASAP7_75t_L g794 ( 
.A(n_585),
.B(n_364),
.C(n_359),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_577),
.B(n_324),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_R g796 ( 
.A(n_610),
.B(n_535),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_669),
.B(n_366),
.Y(n_797)
);

BUFx8_ASAP7_75t_L g798 ( 
.A(n_652),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_650),
.B(n_368),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_669),
.B(n_535),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_650),
.B(n_371),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_567),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_651),
.B(n_375),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_574),
.A2(n_376),
.B1(n_377),
.B2(n_378),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_657),
.B(n_383),
.Y(n_805)
);

NOR3xp33_ASAP7_75t_L g806 ( 
.A(n_574),
.B(n_401),
.C(n_386),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_580),
.A2(n_430),
.B1(n_424),
.B2(n_404),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_778),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_677),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_700),
.B(n_441),
.Y(n_810)
);

AO22x1_ASAP7_75t_L g811 ( 
.A1(n_694),
.A2(n_445),
.B1(n_447),
.B2(n_410),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_745),
.B(n_397),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_707),
.A2(n_512),
.B1(n_655),
.B2(n_659),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_674),
.A2(n_512),
.B(n_655),
.C(n_659),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_800),
.A2(n_548),
.B(n_547),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_737),
.B(n_590),
.Y(n_816)
);

BUFx4f_ASAP7_75t_L g817 ( 
.A(n_734),
.Y(n_817)
);

BUFx12f_ASAP7_75t_L g818 ( 
.A(n_798),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_677),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_680),
.B(n_590),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_789),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_696),
.B(n_32),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_742),
.B(n_33),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_790),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_680),
.B(n_33),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_784),
.A2(n_609),
.B(n_642),
.C(n_641),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_790),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_791),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_709),
.B(n_35),
.Y(n_829)
);

AO21x1_ASAP7_75t_L g830 ( 
.A1(n_714),
.A2(n_600),
.B(n_599),
.Y(n_830)
);

BUFx12f_ASAP7_75t_L g831 ( 
.A(n_798),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_800),
.A2(n_746),
.B(n_744),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_744),
.A2(n_604),
.B(n_600),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_676),
.B(n_36),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_743),
.B(n_37),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_791),
.Y(n_836)
);

AO21x1_ASAP7_75t_L g837 ( 
.A1(n_728),
.A2(n_608),
.B(n_606),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_676),
.B(n_679),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_678),
.B(n_37),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_716),
.B(n_39),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_746),
.A2(n_609),
.B(n_608),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_677),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_685),
.A2(n_622),
.B1(n_638),
.B2(n_633),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_679),
.B(n_39),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_712),
.B(n_40),
.Y(n_845)
);

INVx11_ASAP7_75t_L g846 ( 
.A(n_726),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_673),
.B(n_40),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_698),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_776),
.A2(n_625),
.B(n_624),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_673),
.B(n_41),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_698),
.Y(n_851)
);

NOR3xp33_ASAP7_75t_L g852 ( 
.A(n_694),
.B(n_630),
.C(n_625),
.Y(n_852)
);

BUFx2_ASAP7_75t_SL g853 ( 
.A(n_733),
.Y(n_853)
);

OR2x2_ASAP7_75t_SL g854 ( 
.A(n_683),
.B(n_41),
.Y(n_854)
);

BUFx4f_ASAP7_75t_L g855 ( 
.A(n_734),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_730),
.B(n_42),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_792),
.A2(n_793),
.B(n_782),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_730),
.B(n_43),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_726),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_749),
.B(n_754),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_772),
.A2(n_44),
.B(n_45),
.C(n_47),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_763),
.A2(n_769),
.B(n_773),
.C(n_765),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_774),
.A2(n_467),
.B(n_466),
.C(n_605),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_726),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_706),
.A2(n_684),
.B1(n_701),
.B2(n_692),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_724),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_738),
.B(n_48),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_724),
.A2(n_747),
.B(n_688),
.C(n_697),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_770),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_686),
.B(n_50),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_723),
.B(n_50),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_686),
.B(n_689),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_738),
.B(n_51),
.Y(n_873)
);

INVx3_ASAP7_75t_SL g874 ( 
.A(n_708),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_795),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_806),
.B(n_56),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_717),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_675),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_755),
.B(n_58),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_719),
.B(n_59),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_783),
.A2(n_787),
.B1(n_788),
.B2(n_786),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_753),
.A2(n_63),
.B(n_65),
.C(n_66),
.Y(n_882)
);

O2A1O1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_725),
.A2(n_66),
.B(n_70),
.C(n_71),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_703),
.B(n_70),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_703),
.B(n_73),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_768),
.B(n_75),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_775),
.Y(n_887)
);

OA21x2_ASAP7_75t_L g888 ( 
.A1(n_801),
.A2(n_183),
.B(n_256),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_720),
.B(n_76),
.Y(n_889)
);

AO32x1_ASAP7_75t_L g890 ( 
.A1(n_729),
.A2(n_77),
.A3(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_890)
);

AO21x1_ASAP7_75t_L g891 ( 
.A1(n_803),
.A2(n_80),
.B(n_81),
.Y(n_891)
);

OAI22x1_ASAP7_75t_L g892 ( 
.A1(n_764),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_721),
.B(n_82),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_736),
.B(n_84),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_727),
.B(n_85),
.Y(n_895)
);

AO22x1_ASAP7_75t_L g896 ( 
.A1(n_767),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_731),
.B(n_88),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_804),
.B(n_90),
.Y(n_898)
);

NOR3xp33_ASAP7_75t_L g899 ( 
.A(n_779),
.B(n_90),
.C(n_91),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_732),
.B(n_92),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_710),
.B(n_750),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_799),
.A2(n_691),
.B(n_705),
.C(n_704),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_752),
.B(n_93),
.Y(n_903)
);

OAI321xp33_ASAP7_75t_L g904 ( 
.A1(n_777),
.A2(n_93),
.A3(n_95),
.B1(n_96),
.B2(n_97),
.C(n_98),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_741),
.Y(n_905)
);

BUFx8_ASAP7_75t_SL g906 ( 
.A(n_761),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_713),
.Y(n_907)
);

NAND2x2_ASAP7_75t_L g908 ( 
.A(n_761),
.B(n_97),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_690),
.A2(n_200),
.B(n_242),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_748),
.B(n_99),
.Y(n_910)
);

OAI21xp33_ASAP7_75t_L g911 ( 
.A1(n_807),
.A2(n_756),
.B(n_794),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_681),
.B(n_99),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_L g913 ( 
.A(n_740),
.B(n_100),
.C(n_101),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_682),
.B(n_100),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_715),
.A2(n_101),
.B(n_103),
.C(n_104),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_751),
.B(n_106),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_734),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_718),
.B(n_108),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_693),
.A2(n_136),
.B(n_140),
.C(n_142),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_751),
.B(n_259),
.Y(n_920)
);

AND2x6_ASAP7_75t_L g921 ( 
.A(n_739),
.B(n_143),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_780),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_739),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_699),
.A2(n_149),
.B(n_153),
.Y(n_924)
);

NOR2xp67_ASAP7_75t_L g925 ( 
.A(n_805),
.B(n_154),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_735),
.B(n_687),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_785),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_777),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_702),
.A2(n_169),
.B(n_171),
.Y(n_929)
);

OAI321xp33_ASAP7_75t_L g930 ( 
.A1(n_805),
.A2(n_201),
.A3(n_204),
.B1(n_205),
.B2(n_207),
.C(n_208),
.Y(n_930)
);

AO21x1_ASAP7_75t_L g931 ( 
.A1(n_796),
.A2(n_212),
.B(n_214),
.Y(n_931)
);

AO22x2_ASAP7_75t_L g932 ( 
.A1(n_797),
.A2(n_215),
.B1(n_217),
.B2(n_219),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_781),
.B(n_759),
.Y(n_933)
);

NOR2xp67_ASAP7_75t_L g934 ( 
.A(n_757),
.B(n_758),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_760),
.B(n_232),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_802),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_695),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_762),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_818),
.Y(n_939)
);

NAND3xp33_ASAP7_75t_SL g940 ( 
.A(n_899),
.B(n_766),
.C(n_771),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_869),
.B(n_928),
.Y(n_941)
);

INVxp67_ASAP7_75t_L g942 ( 
.A(n_838),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_836),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_872),
.A2(n_711),
.B1(n_881),
.B2(n_860),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_860),
.B(n_862),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_887),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_855),
.B(n_842),
.Y(n_947)
);

INVx5_ASAP7_75t_L g948 ( 
.A(n_842),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_865),
.B(n_881),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_808),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_865),
.B(n_877),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_876),
.B(n_859),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_821),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_870),
.A2(n_834),
.B1(n_844),
.B2(n_825),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_887),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_833),
.A2(n_849),
.B(n_841),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_868),
.A2(n_911),
.B(n_918),
.C(n_902),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_936),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_938),
.B(n_840),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_926),
.A2(n_820),
.B(n_816),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_909),
.A2(n_929),
.B(n_924),
.Y(n_961)
);

BUFx8_ASAP7_75t_L g962 ( 
.A(n_831),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_856),
.B(n_858),
.Y(n_963)
);

AOI221xp5_ASAP7_75t_L g964 ( 
.A1(n_835),
.A2(n_871),
.B1(n_839),
.B2(n_812),
.C(n_866),
.Y(n_964)
);

CKINVDCx20_ASAP7_75t_R g965 ( 
.A(n_906),
.Y(n_965)
);

OA22x2_ASAP7_75t_L g966 ( 
.A1(n_892),
.A2(n_851),
.B1(n_853),
.B2(n_848),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_887),
.A2(n_901),
.B(n_870),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_810),
.B(n_875),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_867),
.B(n_873),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_826),
.A2(n_847),
.B(n_850),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_894),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_932),
.A2(n_889),
.B1(n_822),
.B2(n_823),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_829),
.B(n_879),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_814),
.A2(n_886),
.B(n_843),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_912),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_888),
.A2(n_912),
.B(n_914),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_874),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_846),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_861),
.A2(n_852),
.B(n_915),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_933),
.B(n_880),
.Y(n_980)
);

NAND2x1p5_ASAP7_75t_L g981 ( 
.A(n_907),
.B(n_923),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_917),
.Y(n_982)
);

OA22x2_ASAP7_75t_L g983 ( 
.A1(n_916),
.A2(n_878),
.B1(n_885),
.B2(n_884),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_895),
.A2(n_897),
.B1(n_903),
.B2(n_893),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_845),
.B(n_910),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_900),
.B(n_935),
.Y(n_986)
);

AO21x2_ASAP7_75t_L g987 ( 
.A1(n_930),
.A2(n_863),
.B(n_919),
.Y(n_987)
);

AOI221xp5_ASAP7_75t_L g988 ( 
.A1(n_882),
.A2(n_878),
.B1(n_883),
.B2(n_896),
.C(n_904),
.Y(n_988)
);

AOI21xp33_ASAP7_75t_L g989 ( 
.A1(n_932),
.A2(n_920),
.B(n_913),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_854),
.B(n_934),
.Y(n_990)
);

NOR2xp67_ASAP7_75t_L g991 ( 
.A(n_813),
.B(n_905),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_922),
.B(n_927),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_925),
.B(n_937),
.Y(n_993)
);

AO21x1_ASAP7_75t_L g994 ( 
.A1(n_890),
.A2(n_921),
.B(n_908),
.Y(n_994)
);

AO31x2_ASAP7_75t_L g995 ( 
.A1(n_890),
.A2(n_830),
.A3(n_837),
.B(n_931),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_824),
.A2(n_827),
.B1(n_836),
.B2(n_828),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_818),
.Y(n_997)
);

CKINVDCx8_ASAP7_75t_R g998 ( 
.A(n_853),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_832),
.A2(n_872),
.B(n_857),
.Y(n_999)
);

INVx5_ASAP7_75t_L g1000 ( 
.A(n_842),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_832),
.A2(n_872),
.B(n_857),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_838),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_824),
.B(n_827),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_832),
.A2(n_872),
.B(n_857),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_832),
.A2(n_872),
.B(n_857),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_824),
.B(n_827),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_832),
.A2(n_872),
.B(n_857),
.Y(n_1007)
);

AO21x2_ASAP7_75t_L g1008 ( 
.A1(n_830),
.A2(n_837),
.B(n_857),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_808),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_818),
.Y(n_1010)
);

AOI21xp33_ASAP7_75t_L g1011 ( 
.A1(n_889),
.A2(n_823),
.B(n_915),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_824),
.B(n_827),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_832),
.A2(n_872),
.B(n_857),
.Y(n_1013)
);

NAND2x1p5_ASAP7_75t_L g1014 ( 
.A(n_817),
.B(n_855),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_824),
.B(n_827),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_898),
.B(n_722),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_SL g1017 ( 
.A1(n_872),
.A2(n_881),
.B(n_827),
.Y(n_1017)
);

NAND2x1p5_ASAP7_75t_L g1018 ( 
.A(n_817),
.B(n_855),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_846),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_838),
.Y(n_1020)
);

BUFx10_ASAP7_75t_L g1021 ( 
.A(n_819),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_842),
.Y(n_1022)
);

AND3x4_ASAP7_75t_L g1023 ( 
.A(n_864),
.B(n_806),
.C(n_798),
.Y(n_1023)
);

OAI21xp33_ASAP7_75t_L g1024 ( 
.A1(n_872),
.A2(n_603),
.B(n_601),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_832),
.A2(n_872),
.B(n_857),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_818),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_846),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_824),
.A2(n_827),
.B1(n_836),
.B2(n_828),
.Y(n_1028)
);

AO31x2_ASAP7_75t_L g1029 ( 
.A1(n_830),
.A2(n_837),
.A3(n_931),
.B(n_832),
.Y(n_1029)
);

OR2x6_ASAP7_75t_L g1030 ( 
.A(n_842),
.B(n_677),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_872),
.A2(n_499),
.B1(n_513),
.B2(n_700),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_832),
.A2(n_857),
.B(n_815),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_824),
.B(n_827),
.Y(n_1033)
);

AOI211x1_ASAP7_75t_L g1034 ( 
.A1(n_891),
.A2(n_911),
.B(n_811),
.C(n_865),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_832),
.A2(n_857),
.B(n_815),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_824),
.B(n_827),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_824),
.B(n_827),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_824),
.B(n_827),
.Y(n_1038)
);

INVxp67_ASAP7_75t_SL g1039 ( 
.A(n_872),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_824),
.B(n_827),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_824),
.B(n_827),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_809),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_872),
.A2(n_499),
.B1(n_513),
.B2(n_700),
.Y(n_1043)
);

INVx4_ASAP7_75t_L g1044 ( 
.A(n_846),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_SL g1045 ( 
.A1(n_872),
.A2(n_860),
.B(n_827),
.Y(n_1045)
);

AOI221xp5_ASAP7_75t_L g1046 ( 
.A1(n_868),
.A2(n_685),
.B1(n_724),
.B2(n_586),
.C(n_688),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_898),
.B(n_722),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_887),
.Y(n_1048)
);

OR2x6_ASAP7_75t_L g1049 ( 
.A(n_842),
.B(n_677),
.Y(n_1049)
);

NOR2xp67_ASAP7_75t_L g1050 ( 
.A(n_818),
.B(n_831),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_842),
.B(n_827),
.Y(n_1051)
);

AOI21xp33_ASAP7_75t_L g1052 ( 
.A1(n_889),
.A2(n_823),
.B(n_915),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_824),
.B(n_827),
.Y(n_1053)
);

NOR2xp67_ASAP7_75t_L g1054 ( 
.A(n_818),
.B(n_831),
.Y(n_1054)
);

BUFx4_ASAP7_75t_SL g1055 ( 
.A(n_809),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_824),
.A2(n_827),
.B(n_836),
.C(n_828),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_824),
.B(n_827),
.Y(n_1057)
);

AO31x2_ASAP7_75t_L g1058 ( 
.A1(n_830),
.A2(n_837),
.A3(n_931),
.B(n_832),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_942),
.Y(n_1059)
);

NAND2x1p5_ASAP7_75t_L g1060 ( 
.A(n_948),
.B(n_1000),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_1024),
.B(n_1016),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_1055),
.Y(n_1062)
);

INVx1_ASAP7_75t_SL g1063 ( 
.A(n_1002),
.Y(n_1063)
);

OR2x6_ASAP7_75t_L g1064 ( 
.A(n_1014),
.B(n_1018),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1045),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1003),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1003),
.Y(n_1067)
);

AO22x2_ASAP7_75t_L g1068 ( 
.A1(n_972),
.A2(n_996),
.B1(n_1028),
.B2(n_1034),
.Y(n_1068)
);

BUFx10_ASAP7_75t_L g1069 ( 
.A(n_1010),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_996),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_1056),
.A2(n_957),
.B(n_999),
.Y(n_1071)
);

CKINVDCx16_ASAP7_75t_R g1072 ( 
.A(n_965),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_1042),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1001),
.A2(n_1005),
.B(n_1004),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1007),
.A2(n_1025),
.B(n_1013),
.Y(n_1075)
);

AOI221xp5_ASAP7_75t_L g1076 ( 
.A1(n_1046),
.A2(n_964),
.B1(n_1028),
.B2(n_1047),
.C(n_1020),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1006),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_SL g1078 ( 
.A1(n_979),
.A2(n_956),
.B(n_989),
.C(n_1011),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1006),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1036),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1036),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_1002),
.B(n_1020),
.Y(n_1082)
);

OAI211xp5_ASAP7_75t_L g1083 ( 
.A1(n_1031),
.A2(n_1043),
.B(n_988),
.C(n_984),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1037),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_959),
.B(n_952),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1037),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_948),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_1000),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1038),
.Y(n_1089)
);

NAND2x1p5_ASAP7_75t_L g1090 ( 
.A(n_1000),
.B(n_1051),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_966),
.A2(n_983),
.B1(n_975),
.B2(n_1053),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1012),
.A2(n_1057),
.B1(n_1033),
.B2(n_1041),
.Y(n_1092)
);

INVx6_ASAP7_75t_L g1093 ( 
.A(n_1019),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_1030),
.B(n_1049),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_1030),
.B(n_1049),
.Y(n_1095)
);

NOR2xp67_ASAP7_75t_L g1096 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_960),
.A2(n_951),
.B(n_1040),
.C(n_1015),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_954),
.A2(n_951),
.B(n_1052),
.C(n_1011),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_943),
.B(n_1022),
.Y(n_1099)
);

NOR2xp67_ASAP7_75t_L g1100 ( 
.A(n_1027),
.B(n_1044),
.Y(n_1100)
);

CKINVDCx6p67_ASAP7_75t_R g1101 ( 
.A(n_939),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_1014),
.Y(n_1102)
);

BUFx2_ASAP7_75t_SL g1103 ( 
.A(n_1050),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_953),
.Y(n_1104)
);

OAI21xp33_ASAP7_75t_L g1105 ( 
.A1(n_985),
.A2(n_1052),
.B(n_973),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_977),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_SL g1107 ( 
.A1(n_945),
.A2(n_970),
.B(n_1035),
.C(n_1032),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_985),
.A2(n_944),
.B(n_979),
.C(n_969),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_958),
.Y(n_1109)
);

INVx1_ASAP7_75t_SL g1110 ( 
.A(n_982),
.Y(n_1110)
);

CKINVDCx6p67_ASAP7_75t_R g1111 ( 
.A(n_997),
.Y(n_1111)
);

NOR2x1_ASAP7_75t_R g1112 ( 
.A(n_1044),
.B(n_1026),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1009),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_963),
.A2(n_969),
.B(n_973),
.C(n_974),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_963),
.A2(n_967),
.B(n_986),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_971),
.A2(n_940),
.B1(n_980),
.B2(n_986),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_1030),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_1049),
.B(n_947),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_SL g1119 ( 
.A(n_962),
.B(n_1054),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_962),
.Y(n_1120)
);

AO21x2_ASAP7_75t_L g1121 ( 
.A1(n_1008),
.A2(n_987),
.B(n_994),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_990),
.A2(n_968),
.B1(n_941),
.B2(n_950),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_978),
.B(n_991),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_992),
.Y(n_1124)
);

CKINVDCx6p67_ASAP7_75t_R g1125 ( 
.A(n_1021),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_981),
.Y(n_1126)
);

OA21x2_ASAP7_75t_L g1127 ( 
.A1(n_995),
.A2(n_1058),
.B(n_1029),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1023),
.A2(n_1021),
.B1(n_993),
.B2(n_955),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_998),
.Y(n_1129)
);

OA21x2_ASAP7_75t_L g1130 ( 
.A1(n_946),
.A2(n_976),
.B(n_961),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_1048),
.A2(n_957),
.B(n_949),
.C(n_1045),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_SL g1132 ( 
.A1(n_1045),
.A2(n_996),
.B1(n_1028),
.B2(n_1039),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_942),
.B(n_1002),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1017),
.A2(n_1045),
.B(n_1039),
.Y(n_1134)
);

AO32x2_ASAP7_75t_L g1135 ( 
.A1(n_972),
.A2(n_954),
.A3(n_1028),
.B1(n_996),
.B2(n_878),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_962),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_1046),
.A2(n_1039),
.B1(n_1045),
.B2(n_1028),
.Y(n_1137)
);

INVxp67_ASAP7_75t_L g1138 ( 
.A(n_1039),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_942),
.B(n_1002),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1045),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_942),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_942),
.B(n_1002),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1045),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1017),
.A2(n_1045),
.B(n_1039),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1067),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1076),
.B(n_1066),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1077),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1080),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_1136),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_1082),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1083),
.A2(n_1092),
.B(n_1108),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1086),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1089),
.Y(n_1153)
);

INVxp67_ASAP7_75t_L g1154 ( 
.A(n_1133),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_1060),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1065),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_1070),
.B(n_1079),
.Y(n_1157)
);

AO21x2_ASAP7_75t_L g1158 ( 
.A1(n_1074),
.A2(n_1075),
.B(n_1071),
.Y(n_1158)
);

AND2x6_ASAP7_75t_L g1159 ( 
.A(n_1140),
.B(n_1143),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1081),
.B(n_1084),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1104),
.B(n_1109),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1085),
.B(n_1059),
.Y(n_1162)
);

INVxp33_ASAP7_75t_L g1163 ( 
.A(n_1112),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1109),
.B(n_1113),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1083),
.A2(n_1108),
.B(n_1114),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1130),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_1070),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_1063),
.B(n_1139),
.Y(n_1168)
);

INVx4_ASAP7_75t_L g1169 ( 
.A(n_1090),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1110),
.B(n_1073),
.Y(n_1170)
);

AO21x1_ASAP7_75t_SL g1171 ( 
.A1(n_1137),
.A2(n_1091),
.B(n_1126),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1115),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1115),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1098),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1114),
.A2(n_1098),
.B(n_1097),
.Y(n_1175)
);

AOI21xp33_ASAP7_75t_L g1176 ( 
.A1(n_1105),
.A2(n_1078),
.B(n_1061),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1141),
.B(n_1142),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_1099),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1134),
.A2(n_1144),
.B(n_1131),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_1138),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1124),
.B(n_1061),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1157),
.B(n_1174),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1156),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1178),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1157),
.B(n_1174),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1163),
.B(n_1119),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1145),
.B(n_1068),
.Y(n_1187)
);

INVxp67_ASAP7_75t_SL g1188 ( 
.A(n_1166),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1159),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1147),
.B(n_1068),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1148),
.B(n_1132),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1153),
.B(n_1068),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1152),
.B(n_1132),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1180),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1165),
.B(n_1107),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1172),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1151),
.B(n_1137),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1172),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1173),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1162),
.B(n_1120),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1159),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1161),
.B(n_1135),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1161),
.B(n_1135),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1180),
.B(n_1127),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1164),
.B(n_1135),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1164),
.B(n_1121),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1160),
.B(n_1116),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1183),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1182),
.B(n_1175),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1182),
.B(n_1185),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1185),
.B(n_1167),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1183),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1206),
.B(n_1158),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1197),
.A2(n_1171),
.B1(n_1146),
.B2(n_1116),
.Y(n_1214)
);

NAND2x1_ASAP7_75t_SL g1215 ( 
.A(n_1189),
.B(n_1169),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1194),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1206),
.B(n_1202),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1202),
.B(n_1158),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1204),
.B(n_1158),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1203),
.B(n_1205),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1188),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1184),
.B(n_1191),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1191),
.B(n_1168),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1193),
.B(n_1168),
.Y(n_1224)
);

NOR2xp67_ASAP7_75t_L g1225 ( 
.A(n_1189),
.B(n_1155),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1208),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1222),
.B(n_1196),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1222),
.B(n_1207),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1221),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_1223),
.B(n_1196),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1208),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1212),
.Y(n_1232)
);

INVxp33_ASAP7_75t_L g1233 ( 
.A(n_1215),
.Y(n_1233)
);

OR2x6_ASAP7_75t_L g1234 ( 
.A(n_1225),
.B(n_1201),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1212),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1217),
.B(n_1187),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1217),
.B(n_1187),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_1223),
.B(n_1198),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_1224),
.B(n_1198),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1216),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1224),
.B(n_1199),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1217),
.B(n_1190),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1210),
.B(n_1207),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1210),
.B(n_1195),
.Y(n_1244)
);

INVxp67_ASAP7_75t_SL g1245 ( 
.A(n_1221),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1220),
.B(n_1190),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1220),
.B(n_1192),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1226),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1226),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1231),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1231),
.Y(n_1251)
);

OR2x2_ASAP7_75t_L g1252 ( 
.A(n_1228),
.B(n_1219),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1246),
.B(n_1220),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1227),
.B(n_1219),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1232),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1240),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1232),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1235),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1235),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1246),
.B(n_1247),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1229),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1247),
.B(n_1213),
.Y(n_1262)
);

OR2x6_ASAP7_75t_L g1263 ( 
.A(n_1234),
.B(n_1225),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1236),
.B(n_1213),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1236),
.B(n_1213),
.Y(n_1265)
);

INVxp67_ASAP7_75t_L g1266 ( 
.A(n_1229),
.Y(n_1266)
);

OAI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1263),
.A2(n_1233),
.B1(n_1234),
.B2(n_1245),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1256),
.A2(n_1214),
.B1(n_1243),
.B2(n_1244),
.Y(n_1268)
);

NOR4xp25_ASAP7_75t_L g1269 ( 
.A(n_1266),
.B(n_1214),
.C(n_1154),
.D(n_1170),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1254),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1261),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1254),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1263),
.A2(n_1234),
.B1(n_1227),
.B2(n_1230),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1261),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1252),
.A2(n_1200),
.B1(n_1218),
.B2(n_1209),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1249),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1252),
.A2(n_1218),
.B1(n_1209),
.B2(n_1197),
.Y(n_1277)
);

NOR2xp67_ASAP7_75t_SL g1278 ( 
.A(n_1263),
.B(n_1103),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1253),
.B(n_1237),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1262),
.A2(n_1218),
.B1(n_1186),
.B2(n_1237),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1249),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1253),
.B(n_1242),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1248),
.Y(n_1283)
);

NOR2x1_ASAP7_75t_L g1284 ( 
.A(n_1263),
.B(n_1234),
.Y(n_1284)
);

OAI21xp33_ASAP7_75t_L g1285 ( 
.A1(n_1262),
.A2(n_1238),
.B(n_1230),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1268),
.B(n_1260),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1271),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1276),
.Y(n_1288)
);

NOR2x1_ASAP7_75t_L g1289 ( 
.A(n_1284),
.B(n_1149),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1277),
.B(n_1260),
.Y(n_1290)
);

AOI21xp33_ASAP7_75t_L g1291 ( 
.A1(n_1267),
.A2(n_1278),
.B(n_1273),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1271),
.B(n_1264),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1275),
.B(n_1285),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1269),
.A2(n_1216),
.B(n_1179),
.Y(n_1294)
);

INVx1_ASAP7_75t_SL g1295 ( 
.A(n_1274),
.Y(n_1295)
);

AOI222xp33_ASAP7_75t_L g1296 ( 
.A1(n_1270),
.A2(n_1150),
.B1(n_1265),
.B2(n_1264),
.C1(n_1255),
.C2(n_1257),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_SL g1297 ( 
.A1(n_1289),
.A2(n_1280),
.B(n_1095),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1291),
.A2(n_1176),
.B(n_1177),
.C(n_1106),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1295),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1287),
.B(n_1296),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1293),
.A2(n_1283),
.B(n_1062),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1294),
.A2(n_1106),
.B(n_1272),
.C(n_1283),
.Y(n_1302)
);

OAI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1286),
.A2(n_1290),
.B1(n_1234),
.B2(n_1292),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1292),
.Y(n_1304)
);

AOI322xp5_ASAP7_75t_L g1305 ( 
.A1(n_1288),
.A2(n_1282),
.A3(n_1279),
.B1(n_1265),
.B2(n_1242),
.C1(n_1281),
.C2(n_1251),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1286),
.B(n_1250),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1289),
.A2(n_1062),
.B(n_1155),
.Y(n_1307)
);

AOI311xp33_ASAP7_75t_L g1308 ( 
.A1(n_1291),
.A2(n_1259),
.A3(n_1257),
.B(n_1250),
.C(n_1255),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1286),
.B(n_1251),
.Y(n_1309)
);

NOR3xp33_ASAP7_75t_L g1310 ( 
.A(n_1298),
.B(n_1072),
.C(n_1129),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1304),
.B(n_1259),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1299),
.B(n_1248),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1305),
.B(n_1258),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1301),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1300),
.Y(n_1315)
);

AND4x1_ASAP7_75t_L g1316 ( 
.A(n_1308),
.B(n_1101),
.C(n_1111),
.D(n_1125),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1306),
.Y(n_1317)
);

OAI322xp33_ASAP7_75t_L g1318 ( 
.A1(n_1303),
.A2(n_1241),
.A3(n_1239),
.B1(n_1238),
.B2(n_1181),
.C1(n_1211),
.C2(n_1195),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1309),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1314),
.B(n_1297),
.Y(n_1320)
);

NOR3xp33_ASAP7_75t_L g1321 ( 
.A(n_1315),
.B(n_1303),
.C(n_1302),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1317),
.B(n_1307),
.Y(n_1322)
);

NAND3xp33_ASAP7_75t_SL g1323 ( 
.A(n_1316),
.B(n_1128),
.C(n_1117),
.Y(n_1323)
);

AOI211xp5_ASAP7_75t_L g1324 ( 
.A1(n_1310),
.A2(n_1129),
.B(n_1100),
.C(n_1096),
.Y(n_1324)
);

NOR2xp67_ASAP7_75t_SL g1325 ( 
.A(n_1312),
.B(n_1087),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_1310),
.Y(n_1326)
);

NAND3xp33_ASAP7_75t_L g1327 ( 
.A(n_1319),
.B(n_1313),
.C(n_1311),
.Y(n_1327)
);

NOR2x1_ASAP7_75t_L g1328 ( 
.A(n_1318),
.B(n_1088),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1322),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1326),
.B(n_1258),
.Y(n_1330)
);

NOR2x1_ASAP7_75t_L g1331 ( 
.A(n_1323),
.B(n_1088),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1320),
.B(n_1239),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1328),
.Y(n_1333)
);

NOR3x2_ASAP7_75t_L g1334 ( 
.A(n_1324),
.B(n_1069),
.C(n_1093),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1321),
.B(n_1325),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1327),
.Y(n_1336)
);

NAND4xp25_ASAP7_75t_L g1337 ( 
.A(n_1326),
.B(n_1094),
.C(n_1122),
.D(n_1123),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1332),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1335),
.B(n_1069),
.Y(n_1339)
);

NOR2x1_ASAP7_75t_L g1340 ( 
.A(n_1329),
.B(n_1064),
.Y(n_1340)
);

XNOR2xp5_ASAP7_75t_L g1341 ( 
.A(n_1334),
.B(n_1123),
.Y(n_1341)
);

OAI22x1_ASAP7_75t_L g1342 ( 
.A1(n_1336),
.A2(n_1169),
.B1(n_1118),
.B2(n_1102),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1339),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_1342),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1338),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1343),
.B(n_1333),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_1346),
.Y(n_1347)
);

OAI21xp33_ASAP7_75t_L g1348 ( 
.A1(n_1346),
.A2(n_1343),
.B(n_1344),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1348),
.B(n_1330),
.Y(n_1349)
);

NOR4xp25_ASAP7_75t_SL g1350 ( 
.A(n_1349),
.B(n_1347),
.C(n_1345),
.D(n_1341),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1350),
.A2(n_1340),
.B(n_1331),
.Y(n_1351)
);

OR2x6_ASAP7_75t_L g1352 ( 
.A(n_1351),
.B(n_1093),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1352),
.A2(n_1337),
.B1(n_1093),
.B2(n_1064),
.Y(n_1353)
);


endmodule