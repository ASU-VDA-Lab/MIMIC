module fake_jpeg_3990_n_216 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_216);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx11_ASAP7_75t_SL g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_33),
.B(n_3),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_23),
.Y(n_51)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_43),
.Y(n_81)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_0),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_47),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_6),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_47),
.A2(n_24),
.B1(n_22),
.B2(n_19),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_48),
.A2(n_76),
.B1(n_13),
.B2(n_7),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_59),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_51),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_16),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_53),
.Y(n_102)
);

NAND2x1p5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_23),
.Y(n_54)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_60),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_20),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_32),
.A2(n_27),
.B1(n_24),
.B2(n_22),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_62),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_103)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_68),
.Y(n_95)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_17),
.Y(n_72)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_40),
.B(n_28),
.Y(n_75)
);

AO22x1_ASAP7_75t_SL g76 ( 
.A1(n_33),
.A2(n_26),
.B1(n_0),
.B2(n_2),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_28),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_35),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_84),
.Y(n_90)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_47),
.B(n_3),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_3),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_26),
.B1(n_4),
.B2(n_5),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_109),
.B1(n_76),
.B2(n_58),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_74),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_64),
.B1(n_61),
.B2(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_8),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_106),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_11),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_9),
.C(n_10),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_49),
.B(n_52),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_87),
.B(n_56),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_116),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_48),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_135),
.B1(n_119),
.B2(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_124),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_82),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_54),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_127),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_101),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_64),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_59),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_110),
.Y(n_128)
);

NOR4xp25_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_67),
.C(n_88),
.D(n_122),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_70),
.B(n_52),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_136),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_102),
.B(n_77),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_77),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

INVx3_ASAP7_75t_SL g155 ( 
.A(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_102),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_92),
.A2(n_70),
.B(n_67),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_156),
.C(n_157),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_140),
.B(n_153),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_107),
.B(n_79),
.C(n_61),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_144),
.B1(n_150),
.B2(n_130),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_57),
.Y(n_167)
);

NAND4xp25_ASAP7_75t_SL g148 ( 
.A(n_133),
.B(n_69),
.C(n_105),
.D(n_68),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_100),
.B1(n_111),
.B2(n_107),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_100),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_125),
.Y(n_161)
);

XNOR2x1_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_65),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_112),
.Y(n_158)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_127),
.B1(n_116),
.B2(n_129),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_164),
.B1(n_141),
.B2(n_144),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_136),
.B(n_131),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_152),
.B(n_143),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_171),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_167),
.B(n_168),
.Y(n_181)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_124),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_172),
.Y(n_183)
);

NOR4xp25_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_143),
.C(n_153),
.D(n_139),
.Y(n_170)
);

OAI322xp33_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_161),
.A3(n_171),
.B1(n_150),
.B2(n_162),
.C1(n_163),
.C2(n_165),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_115),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_176),
.B1(n_180),
.B2(n_151),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_164),
.A2(n_141),
.B1(n_142),
.B2(n_149),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_185),
.B(n_90),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_120),
.C(n_149),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_184),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_141),
.B1(n_113),
.B2(n_121),
.Y(n_180)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_151),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_SL g186 ( 
.A1(n_177),
.A2(n_170),
.B(n_158),
.C(n_155),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_186),
.A2(n_175),
.B(n_179),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_159),
.B1(n_168),
.B2(n_117),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_191),
.Y(n_200)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_188),
.B(n_189),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_192),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_181),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_173),
.A2(n_97),
.B1(n_99),
.B2(n_69),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_97),
.B1(n_99),
.B2(n_128),
.Y(n_194)
);

AOI31xp67_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_180),
.A3(n_155),
.B(n_148),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_195),
.A2(n_186),
.B(n_155),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_174),
.B(n_175),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_201),
.B(n_182),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_202),
.A2(n_205),
.A3(n_200),
.B1(n_186),
.B2(n_199),
.C1(n_185),
.C2(n_184),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_197),
.A2(n_186),
.B1(n_190),
.B2(n_182),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_206),
.B1(n_166),
.B2(n_11),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_208),
.C(n_105),
.Y(n_211)
);

AOI322xp5_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_200),
.A3(n_90),
.B1(n_166),
.B2(n_96),
.C1(n_57),
.C2(n_105),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

AOI21x1_ASAP7_75t_L g210 ( 
.A1(n_203),
.A2(n_105),
.B(n_10),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_210),
.A2(n_91),
.B(n_93),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_211),
.A2(n_93),
.B(n_213),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_91),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_215),
.Y(n_216)
);


endmodule