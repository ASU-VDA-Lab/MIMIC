module fake_jpeg_19175_n_319 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_319);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx11_ASAP7_75t_SL g12 ( 
.A(n_5),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_23),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_26),
.Y(n_44)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_18),
.B(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_31),
.B(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_58),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_30),
.Y(n_48)
);

FAx1_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_41),
.CI(n_12),
.CON(n_63),
.SN(n_63)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_20),
.B1(n_17),
.B2(n_13),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_28),
.B1(n_39),
.B2(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_52),
.B(n_53),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_25),
.B1(n_33),
.B2(n_27),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_43),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_26),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_33),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_79),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_25),
.B1(n_32),
.B2(n_30),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_48),
.B1(n_46),
.B2(n_27),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_28),
.B1(n_56),
.B2(n_60),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_13),
.B1(n_20),
.B2(n_25),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_76),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_38),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_58),
.B(n_59),
.Y(n_90)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_47),
.B(n_13),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_78),
.Y(n_89)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_62),
.B1(n_52),
.B2(n_55),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_69),
.B1(n_63),
.B2(n_29),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_SL g122 ( 
.A1(n_88),
.A2(n_94),
.B(n_64),
.C(n_63),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_92),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_68),
.Y(n_111)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_51),
.B(n_54),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_71),
.B(n_75),
.Y(n_117)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_61),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_96),
.B(n_98),
.Y(n_115)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_32),
.C(n_29),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_63),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_20),
.B1(n_35),
.B2(n_23),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_104),
.B(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_81),
.B1(n_66),
.B2(n_69),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_118),
.B1(n_101),
.B2(n_92),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_108),
.B(n_109),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_65),
.B1(n_56),
.B2(n_77),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_39),
.B1(n_49),
.B2(n_42),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_111),
.A2(n_112),
.B(n_117),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_81),
.B(n_78),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_86),
.B(n_82),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_116),
.B(n_128),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_69),
.B1(n_71),
.B2(n_68),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_121),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_39),
.B(n_35),
.C(n_43),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_101),
.B(n_63),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_84),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_49),
.Y(n_157)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_130),
.B(n_139),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_140),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_138),
.A2(n_141),
.B1(n_147),
.B2(n_40),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_103),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_80),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_95),
.B1(n_98),
.B2(n_85),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_106),
.A2(n_77),
.B1(n_65),
.B2(n_36),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_153),
.B1(n_159),
.B2(n_40),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_80),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_149),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_120),
.B(n_106),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_145),
.Y(n_184)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_65),
.B1(n_56),
.B2(n_60),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_148),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_127),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_154),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_65),
.C(n_10),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_158),
.C(n_9),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_157),
.Y(n_175)
);

AOI32xp33_ASAP7_75t_L g158 ( 
.A1(n_109),
.A2(n_17),
.A3(n_28),
.B1(n_16),
.B2(n_19),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_28),
.B1(n_18),
.B2(n_15),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_17),
.B1(n_18),
.B2(n_16),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_164),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_122),
.B(n_22),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_161),
.B(n_22),
.Y(n_169)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_122),
.A2(n_16),
.B(n_22),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_122),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_183),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_166),
.A2(n_137),
.B1(n_159),
.B2(n_133),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_38),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_136),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_170),
.B(n_186),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_179),
.B1(n_190),
.B2(n_194),
.Y(n_201)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_16),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_151),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_135),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_135),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_134),
.B(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_143),
.B(n_16),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_164),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_15),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_165),
.B(n_131),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_195),
.B(n_199),
.Y(n_241)
);

HAxp5_ASAP7_75t_SL g198 ( 
.A(n_173),
.B(n_189),
.CON(n_198),
.SN(n_198)
);

NOR2x1_ASAP7_75t_R g229 ( 
.A(n_198),
.B(n_211),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_183),
.B(n_138),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_207),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_204),
.B(n_209),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_182),
.B1(n_172),
.B2(n_178),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_137),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_181),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_144),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_216),
.Y(n_226)
);

XOR2x1_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_162),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_192),
.C(n_167),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_219),
.C(n_185),
.Y(n_235)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_133),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_217),
.Y(n_224)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_166),
.B(n_141),
.C(n_150),
.Y(n_219)
);

NOR3xp33_ASAP7_75t_SL g222 ( 
.A(n_211),
.B(n_176),
.C(n_190),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_230),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_228),
.A2(n_148),
.B1(n_1),
.B2(n_2),
.Y(n_257)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_175),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_232),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_182),
.B1(n_178),
.B2(n_176),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_236),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_238),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_191),
.C(n_168),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_216),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_239),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_168),
.Y(n_238)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_199),
.B(n_179),
.CI(n_147),
.CON(n_239),
.SN(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_184),
.B(n_188),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_242),
.B(n_9),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_197),
.A2(n_145),
.B(n_130),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_198),
.B(n_210),
.Y(n_243)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_206),
.B(n_203),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_244),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_241),
.B(n_196),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_249),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_196),
.C(n_201),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_238),
.B(n_226),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_200),
.Y(n_249)
);

INVx13_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_253),
.Y(n_262)
);

INVx13_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

INVx13_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_259),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_257),
.A2(n_260),
.B1(n_225),
.B2(n_239),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_16),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_22),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_235),
.A2(n_21),
.B1(n_40),
.B2(n_8),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_236),
.C(n_223),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_261),
.B(n_266),
.Y(n_283)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_264),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_226),
.C(n_239),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_222),
.C(n_34),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_273),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_258),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_248),
.A2(n_19),
.B1(n_21),
.B2(n_14),
.Y(n_271)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_252),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_244),
.B(n_251),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_34),
.C(n_38),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_250),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_278),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_255),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_281),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_257),
.B1(n_243),
.B2(n_260),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_268),
.B1(n_265),
.B2(n_8),
.Y(n_289)
);

AOI21x1_ASAP7_75t_SL g285 ( 
.A1(n_274),
.A2(n_253),
.B(n_249),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_277),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_19),
.B(n_22),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_4),
.B(n_6),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_21),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_34),
.C(n_38),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_267),
.C(n_273),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_290),
.Y(n_307)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_34),
.C(n_38),
.Y(n_290)
);

OAI21x1_ASAP7_75t_SL g292 ( 
.A1(n_275),
.A2(n_21),
.B(n_5),
.Y(n_292)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_293),
.B(n_294),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_6),
.B1(n_8),
.B2(n_4),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_6),
.B1(n_7),
.B2(n_4),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_297),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_285),
.B1(n_281),
.B2(n_7),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_38),
.C(n_14),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_7),
.B(n_6),
.Y(n_300)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_305),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_14),
.C(n_7),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_298),
.B(n_3),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_0),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_310),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_301),
.A2(n_296),
.B1(n_308),
.B2(n_288),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_307),
.A3(n_302),
.B1(n_304),
.B2(n_290),
.C1(n_1),
.C2(n_3),
.Y(n_314)
);

NAND4xp25_ASAP7_75t_SL g315 ( 
.A(n_314),
.B(n_309),
.C(n_311),
.D(n_312),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_313),
.B(n_307),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_0),
.C(n_3),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_3),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_3),
.Y(n_319)
);


endmodule