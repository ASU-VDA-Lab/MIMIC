module fake_jpeg_31416_n_90 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_90);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_90;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx4f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_6),
.B(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_15),
.Y(n_43)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_29),
.A2(n_23),
.B1(n_20),
.B2(n_16),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_21),
.B1(n_20),
.B2(n_22),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_51),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_30),
.B(n_31),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_53),
.B(n_55),
.C(n_37),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_30),
.B1(n_33),
.B2(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_52),
.Y(n_67)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_26),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_21),
.B1(n_32),
.B2(n_27),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_57),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

AOI22x1_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_53),
.B1(n_46),
.B2(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_40),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_54),
.B(n_56),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_67),
.B(n_62),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_13),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_72),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_44),
.C(n_34),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_76),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_66),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_66),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_0),
.B(n_1),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_38),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_73),
.C(n_38),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_77),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_85),
.C(n_86),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_82),
.C(n_32),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_32),
.B(n_7),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_87),
.C(n_10),
.Y(n_90)
);


endmodule