module fake_jpeg_31594_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

INVx11_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_35),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_3),
.B(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_56),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_49),
.B(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_60),
.Y(n_74)
);

AND2x4_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_2),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_61),
.B(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_46),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_73),
.Y(n_85)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_4),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_70),
.B1(n_66),
.B2(n_51),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_89),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_39),
.B(n_43),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_84),
.B(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_65),
.B(n_47),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_46),
.B(n_38),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_45),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_50),
.Y(n_89)
);

BUFx16f_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_88),
.B(n_3),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_94),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_41),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_13),
.C(n_14),
.Y(n_109)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_96),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_5),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_5),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_36),
.B1(n_41),
.B2(n_11),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_103),
.A2(n_22),
.B1(n_26),
.B2(n_29),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_8),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_108),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_106),
.A2(n_15),
.B(n_19),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_78),
.B(n_9),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_113),
.C(n_118),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_20),
.C(n_21),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_30),
.C(n_31),
.Y(n_118)
);

AOI221xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_103),
.B1(n_100),
.B2(n_101),
.C(n_107),
.Y(n_119)
);

BUFx12f_ASAP7_75t_SL g125 ( 
.A(n_119),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_101),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_116),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_126),
.Y(n_127)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_125),
.C(n_122),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_117),
.C(n_123),
.Y(n_129)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_116),
.B(n_115),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_131),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_100),
.Y(n_133)
);


endmodule