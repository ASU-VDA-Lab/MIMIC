module fake_jpeg_11867_n_363 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_363);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_363;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_22),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g152 ( 
.A(n_54),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_57),
.Y(n_140)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_39),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_66),
.B(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

BUFx4f_ASAP7_75t_SL g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_20),
.B(n_7),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_73),
.A2(n_78),
.B(n_83),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_22),
.Y(n_74)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_75),
.Y(n_156)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_22),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_20),
.B(n_7),
.Y(n_78)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_38),
.B(n_7),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_80),
.B(n_89),
.Y(n_142)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_27),
.B(n_34),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_42),
.B(n_0),
.Y(n_93)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_27),
.B(n_9),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_96),
.Y(n_110)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_98),
.Y(n_113)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_29),
.B(n_13),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_103),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_33),
.B(n_1),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_54),
.A2(n_42),
.B1(n_40),
.B2(n_24),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_105),
.A2(n_125),
.B1(n_127),
.B2(n_133),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_34),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_124),
.B(n_126),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_74),
.A2(n_42),
.B1(n_24),
.B2(n_44),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_73),
.A2(n_29),
.B(n_47),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_90),
.A2(n_53),
.B1(n_44),
.B2(n_41),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_66),
.A2(n_47),
.B1(n_41),
.B2(n_46),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_78),
.B(n_46),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_135),
.B(n_139),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_90),
.A2(n_53),
.B1(n_48),
.B2(n_45),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_136),
.A2(n_138),
.B1(n_145),
.B2(n_31),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_62),
.A2(n_48),
.B1(n_45),
.B2(n_43),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_23),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_23),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_149),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_65),
.A2(n_43),
.B1(n_52),
.B2(n_51),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_93),
.B(n_51),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_147),
.B(n_150),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_52),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_80),
.B(n_49),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_55),
.A2(n_50),
.B1(n_49),
.B2(n_36),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_153),
.B(n_105),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_57),
.B(n_36),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_162),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_68),
.A2(n_50),
.B1(n_26),
.B2(n_3),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_60),
.B(n_26),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_164),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_107),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_165),
.A2(n_196),
.B(n_199),
.Y(n_255)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_167),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_86),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_170),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_149),
.A2(n_63),
.B1(n_85),
.B2(n_82),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_171),
.A2(n_179),
.B1(n_187),
.B2(n_205),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_163),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_172),
.B(n_173),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_110),
.B(n_69),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_118),
.B(n_10),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_174),
.B(n_182),
.Y(n_229)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_138),
.A2(n_79),
.B1(n_99),
.B2(n_31),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_180),
.Y(n_256)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_117),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_183),
.B(n_185),
.Y(n_239)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_184),
.A2(n_193),
.B(n_194),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_116),
.B(n_12),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_186),
.B(n_190),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_145),
.A2(n_31),
.B1(n_12),
.B2(n_11),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_188),
.A2(n_189),
.B1(n_123),
.B2(n_119),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_121),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_191),
.A2(n_195),
.B1(n_198),
.B2(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_106),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_125),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_197),
.Y(n_220)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_129),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_163),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_204),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_127),
.B1(n_148),
.B2(n_111),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_136),
.Y(n_203)
);

NOR3xp33_ASAP7_75t_SL g254 ( 
.A(n_203),
.B(n_204),
.C(n_195),
.Y(n_254)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_152),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_120),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_207),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_142),
.B(n_4),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_142),
.B(n_152),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_209),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_152),
.B(n_144),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_141),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_212),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_158),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_114),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_106),
.Y(n_231)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_114),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_112),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_216),
.A2(n_146),
.B(n_108),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_203),
.B1(n_216),
.B2(n_168),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_218),
.A2(n_228),
.B1(n_237),
.B2(n_241),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_224),
.B(n_225),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_175),
.A2(n_151),
.B1(n_109),
.B2(n_119),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_231),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_232),
.A2(n_242),
.B(n_220),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_188),
.A2(n_112),
.B1(n_151),
.B2(n_109),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_244),
.B1(n_167),
.B2(n_180),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_176),
.B(n_146),
.C(n_160),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_236),
.C(n_240),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_111),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_181),
.A2(n_123),
.B1(n_160),
.B2(n_148),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_192),
.B(n_158),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_196),
.A2(n_131),
.B1(n_140),
.B2(n_158),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_166),
.A2(n_131),
.B(n_140),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_189),
.A2(n_202),
.B1(n_193),
.B2(n_178),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_192),
.A2(n_211),
.B(n_165),
.C(n_177),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_218),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_202),
.A2(n_206),
.B1(n_215),
.B2(n_198),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_202),
.A2(n_200),
.B1(n_191),
.B2(n_210),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_182),
.A2(n_190),
.B1(n_183),
.B2(n_199),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_164),
.A2(n_186),
.B1(n_214),
.B2(n_194),
.Y(n_251)
);

NOR3xp33_ASAP7_75t_SL g265 ( 
.A(n_254),
.B(n_243),
.C(n_230),
.Y(n_265)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_258),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_259),
.A2(n_286),
.B1(n_241),
.B2(n_257),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_184),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_260),
.B(n_266),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_170),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_261),
.B(n_270),
.C(n_288),
.Y(n_305)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_227),
.Y(n_263)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_264),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_SL g295 ( 
.A1(n_265),
.A2(n_268),
.A3(n_269),
.B1(n_281),
.B2(n_242),
.C1(n_219),
.C2(n_231),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_229),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_222),
.B(n_243),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_222),
.B(n_236),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_275),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_272),
.A2(n_281),
.B(n_275),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_247),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_279),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_238),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_234),
.B(n_238),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_278),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_223),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_234),
.B(n_226),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_228),
.A2(n_249),
.B1(n_248),
.B2(n_220),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_280),
.A2(n_277),
.B1(n_262),
.B2(n_282),
.Y(n_291)
);

NOR4xp25_ASAP7_75t_L g281 ( 
.A(n_232),
.B(n_223),
.C(n_255),
.D(n_254),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_221),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_283),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_221),
.B(n_252),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_250),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_285),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_237),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_224),
.A2(n_219),
.B1(n_217),
.B2(n_225),
.Y(n_286)
);

INVx3_ASAP7_75t_SL g287 ( 
.A(n_253),
.Y(n_287)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_287),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_256),
.B(n_235),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_261),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_291),
.B(n_301),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_294),
.A2(n_302),
.B(n_296),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_253),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_296),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_276),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_280),
.A2(n_245),
.B1(n_277),
.B2(n_273),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_272),
.A2(n_271),
.B(n_278),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_308),
.B(n_309),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_304),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_310),
.C(n_308),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_283),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_274),
.A2(n_270),
.B(n_267),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_268),
.A2(n_269),
.B(n_266),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_310),
.B(n_311),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_260),
.Y(n_311)
);

OAI32xp33_ASAP7_75t_SL g314 ( 
.A1(n_303),
.A2(n_262),
.A3(n_265),
.B1(n_286),
.B2(n_267),
.Y(n_314)
);

AOI321xp33_ASAP7_75t_L g330 ( 
.A1(n_314),
.A2(n_293),
.A3(n_295),
.B1(n_305),
.B2(n_296),
.C(n_297),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_291),
.A2(n_258),
.B1(n_263),
.B2(n_287),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_315),
.A2(n_316),
.B(n_320),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_308),
.A2(n_264),
.B(n_287),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_289),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_323),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_307),
.C(n_313),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g322 ( 
.A1(n_302),
.A2(n_294),
.B(n_292),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_322),
.A2(n_298),
.B1(n_307),
.B2(n_324),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_299),
.B(n_300),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_300),
.B(n_290),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_325),
.B(n_322),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_L g327 ( 
.A1(n_292),
.A2(n_312),
.B(n_306),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_305),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_314),
.Y(n_345)
);

XNOR2x1_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_338),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_324),
.A2(n_289),
.B1(n_297),
.B2(n_296),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_332),
.A2(n_318),
.B1(n_326),
.B2(n_331),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_333),
.Y(n_341)
);

AOI322xp5_ASAP7_75t_L g334 ( 
.A1(n_319),
.A2(n_298),
.A3(n_307),
.B1(n_323),
.B2(n_317),
.C1(n_320),
.C2(n_314),
.Y(n_334)
);

INVx6_ASAP7_75t_L g344 ( 
.A(n_334),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_336),
.C(n_322),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_316),
.C(n_322),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_345),
.Y(n_351)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_328),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_342),
.B(n_343),
.Y(n_350)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_332),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_315),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_346),
.B(n_345),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_337),
.A2(n_326),
.B(n_336),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_348),
.B(n_347),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_341),
.A2(n_335),
.B1(n_337),
.B2(n_330),
.Y(n_349)
);

OAI21x1_ASAP7_75t_L g358 ( 
.A1(n_352),
.A2(n_353),
.B(n_354),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_340),
.Y(n_354)
);

AOI31xp67_ASAP7_75t_SL g355 ( 
.A1(n_350),
.A2(n_339),
.A3(n_348),
.B(n_346),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_355),
.B(n_356),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_349),
.A2(n_339),
.B(n_353),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_351),
.B(n_329),
.C(n_340),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_358),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_359),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_361),
.B(n_357),
.C(n_360),
.Y(n_362)
);

INVxp33_ASAP7_75t_L g363 ( 
.A(n_362),
.Y(n_363)
);


endmodule