module fake_jpeg_2004_n_192 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_192);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_36),
.Y(n_55)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_12),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_22),
.B(n_11),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_11),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_18),
.B(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_16),
.B1(n_25),
.B2(n_26),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_53),
.A2(n_58),
.B1(n_73),
.B2(n_21),
.Y(n_86)
);

CKINVDCx12_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_80),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_22),
.B1(n_20),
.B2(n_25),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_29),
.B1(n_27),
.B2(n_15),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_60),
.A2(n_32),
.B(n_6),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_61),
.B(n_65),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_15),
.C(n_26),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_72),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_79),
.Y(n_83)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_27),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_33),
.A2(n_16),
.B1(n_29),
.B2(n_27),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_74),
.B(n_10),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_35),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_32),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_10),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_38),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_1),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_85),
.B(n_91),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_52),
.B1(n_76),
.B2(n_32),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_77),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_72),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_4),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_105),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_57),
.B(n_5),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_97),
.Y(n_121)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_5),
.Y(n_97)
);

OR2x4_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_21),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_98),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_101),
.A2(n_72),
.B1(n_75),
.B2(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_74),
.B(n_6),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_104),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_77),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_7),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_98),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_106),
.B(n_119),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_62),
.C(n_50),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_113),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_71),
.B1(n_70),
.B2(n_76),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_112),
.B1(n_120),
.B2(n_125),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_75),
.C(n_63),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_116),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_82),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_115),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_55),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_59),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_89),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_122),
.B(n_104),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_86),
.A2(n_67),
.B1(n_78),
.B2(n_7),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_123),
.A2(n_94),
.B1(n_101),
.B2(n_105),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_128),
.B1(n_132),
.B2(n_135),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_125),
.A2(n_91),
.B1(n_96),
.B2(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_136),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_100),
.B1(n_83),
.B2(n_90),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_88),
.B1(n_67),
.B2(n_87),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_110),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_87),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_144),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_92),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_140),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_143),
.Y(n_149)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_134),
.A2(n_115),
.B(n_113),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_145),
.A2(n_133),
.B(n_128),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_115),
.C(n_114),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_151),
.C(n_142),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_144),
.A2(n_113),
.B1(n_117),
.B2(n_107),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_156),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_119),
.C(n_117),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_153),
.B(n_127),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_88),
.B1(n_99),
.B2(n_78),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_158),
.A2(n_161),
.B(n_165),
.Y(n_171)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_152),
.B(n_129),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_142),
.C(n_137),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_138),
.C(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_155),
.B1(n_150),
.B2(n_149),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_145),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_163),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_146),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_178),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_177),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_173),
.A2(n_153),
.B1(n_146),
.B2(n_156),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_155),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_168),
.C(n_171),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_78),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_173),
.B(n_157),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_170),
.B(n_157),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_175),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_186),
.Y(n_188)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

OAI21x1_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_180),
.B(n_182),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_187),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_99),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_7),
.Y(n_192)
);


endmodule