module fake_jpeg_6056_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_37),
.C(n_41),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_43),
.Y(n_63)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_44),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_46),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_21),
.B1(n_23),
.B2(n_28),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_49),
.A2(n_66),
.B1(n_70),
.B2(n_28),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_23),
.B1(n_21),
.B2(n_29),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_73)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_55),
.Y(n_74)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_34),
.A2(n_21),
.B1(n_23),
.B2(n_29),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_64),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_23),
.B1(n_26),
.B2(n_18),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_26),
.B1(n_18),
.B2(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_28),
.B1(n_31),
.B2(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_22),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_69),
.Y(n_94)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_71),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_42),
.B(n_41),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_83),
.B(n_19),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_42),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_86),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_44),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_84),
.C(n_85),
.Y(n_101)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_88),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_35),
.C(n_31),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_24),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_31),
.B(n_35),
.C(n_33),
.Y(n_83)
);

OR2x2_ASAP7_75t_SL g84 ( 
.A(n_62),
.B(n_14),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_64),
.B(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_30),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_50),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_93),
.A2(n_52),
.B1(n_57),
.B2(n_45),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_112),
.B1(n_118),
.B2(n_77),
.Y(n_129)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_67),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_121),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_116),
.B(n_76),
.Y(n_123)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_104),
.B(n_115),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_73),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_105),
.A2(n_107),
.B1(n_119),
.B2(n_78),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_65),
.B1(n_70),
.B2(n_45),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_19),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_111),
.B(n_113),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_85),
.A2(n_70),
.B1(n_45),
.B2(n_58),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_30),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_30),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_58),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_76),
.A2(n_24),
.B(n_46),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_82),
.Y(n_117)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_32),
.B1(n_25),
.B2(n_35),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_35),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_127),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_125),
.B(n_138),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_81),
.C(n_76),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_130),
.C(n_140),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_85),
.B(n_83),
.Y(n_125)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_126),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_136),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_129),
.A2(n_142),
.B1(n_117),
.B2(n_103),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_71),
.C(n_83),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_84),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_96),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_101),
.A2(n_94),
.B(n_91),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_113),
.B(n_114),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_99),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_74),
.B1(n_91),
.B2(n_77),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_137),
.A2(n_141),
.B1(n_143),
.B2(n_119),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_116),
.A2(n_88),
.B(n_35),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_87),
.C(n_68),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_89),
.B1(n_32),
.B2(n_25),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_110),
.A2(n_78),
.B1(n_32),
.B2(n_25),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_101),
.A2(n_24),
.B(n_33),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_144),
.A2(n_111),
.B(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_105),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_149),
.A2(n_159),
.B(n_163),
.Y(n_196)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_139),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_97),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_167),
.Y(n_185)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_168),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_158),
.B1(n_162),
.B2(n_172),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_119),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_160),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_107),
.B1(n_109),
.B2(n_118),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_131),
.B(n_118),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_147),
.A2(n_107),
.B1(n_118),
.B2(n_96),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_131),
.B(n_104),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_169),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_123),
.A2(n_106),
.B(n_115),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_173),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_SL g171 ( 
.A1(n_138),
.A2(n_24),
.B(n_33),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_24),
.Y(n_197)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_87),
.C(n_90),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_152),
.C(n_160),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_166),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_176),
.B(n_180),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_170),
.A2(n_130),
.B1(n_142),
.B2(n_141),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_193),
.B1(n_89),
.B2(n_32),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_153),
.Y(n_179)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_150),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_183),
.C(n_156),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_127),
.C(n_128),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_167),
.A2(n_134),
.B(n_132),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_184),
.A2(n_24),
.B1(n_27),
.B2(n_33),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_146),
.Y(n_186)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_134),
.C(n_146),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_190),
.Y(n_203)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_192),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_162),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_168),
.A2(n_145),
.B1(n_103),
.B2(n_122),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_197),
.Y(n_218)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_149),
.B(n_145),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_200),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_161),
.B1(n_159),
.B2(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_187),
.A2(n_161),
.B1(n_159),
.B2(n_158),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_217),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_212),
.Y(n_229)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_211),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_210),
.C(n_222),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_165),
.C(n_90),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_90),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_214),
.A2(n_196),
.B(n_185),
.Y(n_226)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_220),
.Y(n_231)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_223),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_139),
.C(n_89),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_179),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_139),
.C(n_33),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_178),
.C(n_175),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_196),
.B(n_191),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_214),
.Y(n_247)
);

NAND2xp33_ASAP7_75t_SL g255 ( 
.A(n_226),
.B(n_230),
.Y(n_255)
);

INVxp33_ASAP7_75t_SL g227 ( 
.A(n_223),
.Y(n_227)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

NOR2xp67_ASAP7_75t_SL g230 ( 
.A(n_222),
.B(n_210),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_181),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_234),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_181),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_184),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_206),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_239),
.C(n_241),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_213),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_238),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_188),
.C(n_197),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_179),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_33),
.C(n_27),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_244),
.C(n_206),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_27),
.C(n_25),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_204),
.B(n_10),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_245),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_256),
.C(n_261),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_209),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

OAI321xp33_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_217),
.A3(n_209),
.B1(n_203),
.B2(n_218),
.C(n_216),
.Y(n_251)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_237),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_258),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_203),
.Y(n_254)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_228),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_260),
.Y(n_276)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_223),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_229),
.B(n_216),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_239),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_27),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_266),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_232),
.C(n_229),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_268),
.C(n_272),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_232),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_244),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_270),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_255),
.B(n_242),
.Y(n_268)
);

BUFx24_ASAP7_75t_SL g270 ( 
.A(n_249),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_246),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_271),
.A2(n_278),
.B1(n_254),
.B2(n_274),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_27),
.C(n_4),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_277),
.A2(n_12),
.B(n_5),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_256),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_284),
.B(n_285),
.Y(n_291)
);

O2A1O1Ixp33_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_248),
.B(n_255),
.C(n_246),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_282),
.B(n_283),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_263),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_290),
.Y(n_294)
);

NOR2x1_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_257),
.Y(n_289)
);

NOR3xp33_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_10),
.C(n_5),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_272),
.B(n_11),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_265),
.C(n_5),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_299),
.B(n_300),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_287),
.B(n_11),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_298),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_11),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_297),
.B(n_295),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_3),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_6),
.C(n_7),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_279),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_304),
.B(n_306),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_15),
.B(n_13),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_279),
.B(n_289),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_292),
.A2(n_3),
.B(n_6),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_7),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_307),
.A2(n_308),
.B(n_15),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_305),
.C(n_12),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_311),
.B(n_312),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_7),
.C(n_12),
.Y(n_311)
);

AO21x1_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_13),
.B(n_14),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_314),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_316),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_315),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_310),
.Y(n_319)
);


endmodule