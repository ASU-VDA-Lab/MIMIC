module real_aes_4020_n_407 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_401, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_399, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_400, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_398, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_405, n_368, n_250, n_85, n_406, n_45, n_5, n_244, n_118, n_139, n_402, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_404, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_1349, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_403, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_407);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_401;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_399;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_400;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_398;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_405;
input n_368;
input n_250;
input n_85;
input n_406;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_402;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_404;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_1349;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_403;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_407;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_592;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_795;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1325;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_417;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_1342;
wire n_1346;
wire n_552;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_829;
wire n_1030;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_994;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_617;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_1298;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_905;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_816;
wire n_625;
wire n_953;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_632;
wire n_1344;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_1083;
wire n_727;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1240;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_698;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_483;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_1236;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_0), .A2(n_283), .B1(n_846), .B2(n_855), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g1319 ( .A1(n_1), .A2(n_6), .B1(n_1320), .B2(n_1321), .Y(n_1319) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_2), .A2(n_60), .B1(n_882), .B2(n_1024), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_3), .A2(n_209), .B1(n_847), .B2(n_853), .Y(n_1137) );
AOI22xp5_ASAP7_75t_L g1220 ( .A1(n_4), .A2(n_216), .B1(n_880), .B2(n_962), .Y(n_1220) );
AOI22xp33_ASAP7_75t_L g1234 ( .A1(n_5), .A2(n_162), .B1(n_849), .B2(n_850), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_7), .A2(n_176), .B1(n_805), .B2(n_806), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_8), .A2(n_351), .B1(n_847), .B2(n_853), .Y(n_1010) );
INVx1_ASAP7_75t_L g1041 ( .A(n_9), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_10), .A2(n_179), .B1(n_707), .B2(n_894), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1281 ( .A1(n_11), .A2(n_101), .B1(n_660), .B2(n_882), .Y(n_1281) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_12), .A2(n_48), .B1(n_713), .B2(n_893), .Y(n_1027) );
INVx1_ASAP7_75t_L g937 ( .A(n_13), .Y(n_937) );
AOI21x1_ASAP7_75t_L g1035 ( .A1(n_14), .A2(n_1036), .B(n_1040), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_15), .A2(n_367), .B1(n_805), .B2(n_964), .Y(n_1240) );
INVx1_ASAP7_75t_L g957 ( .A(n_16), .Y(n_957) );
AOI22xp5_ASAP7_75t_L g1246 ( .A1(n_17), .A2(n_329), .B1(n_746), .B2(n_812), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_18), .A2(n_35), .B1(n_703), .B2(n_898), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g1282 ( .A1(n_19), .A2(n_103), .B1(n_805), .B2(n_1283), .Y(n_1282) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_20), .A2(n_116), .B1(n_722), .B2(n_962), .Y(n_1059) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_21), .B(n_666), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_22), .A2(n_212), .B1(n_746), .B2(n_815), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1323 ( .A1(n_23), .A2(n_287), .B1(n_1324), .B2(n_1325), .Y(n_1323) );
CKINVDCx20_ASAP7_75t_R g1117 ( .A(n_24), .Y(n_1117) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_25), .A2(n_370), .B1(n_427), .B2(n_435), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_26), .A2(n_267), .B1(n_849), .B2(n_850), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_27), .B(n_913), .Y(n_912) );
AOI22xp5_ASAP7_75t_L g1080 ( .A1(n_28), .A2(n_222), .B1(n_834), .B2(n_856), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_29), .A2(n_256), .B1(n_808), .B2(n_924), .Y(n_966) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_30), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_31), .A2(n_369), .B1(n_951), .B2(n_1034), .Y(n_1208) );
AOI22xp5_ASAP7_75t_L g908 ( .A1(n_32), .A2(n_76), .B1(n_909), .B2(n_911), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g1244 ( .A1(n_33), .A2(n_160), .B1(n_882), .B2(n_1024), .Y(n_1244) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_34), .A2(n_45), .B1(n_659), .B2(n_685), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g1272 ( .A1(n_36), .A2(n_239), .B1(n_735), .B2(n_905), .Y(n_1272) );
INVx1_ASAP7_75t_L g889 ( .A(n_37), .Y(n_889) );
INVx1_ASAP7_75t_L g1267 ( .A(n_38), .Y(n_1267) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_39), .A2(n_300), .B1(n_962), .B2(n_964), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_40), .B(n_959), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_41), .A2(n_107), .B1(n_855), .B2(n_856), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_42), .A2(n_403), .B1(n_834), .B2(n_856), .Y(n_1235) );
XOR2x2_ASAP7_75t_L g1071 ( .A(n_43), .B(n_1072), .Y(n_1071) );
AOI22xp33_ASAP7_75t_SL g1134 ( .A1(n_44), .A2(n_390), .B1(n_835), .B2(n_951), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_46), .A2(n_157), .B1(n_805), .B2(n_924), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_47), .A2(n_115), .B1(n_746), .B2(n_815), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_49), .A2(n_142), .B1(n_746), .B2(n_815), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_50), .A2(n_168), .B1(n_875), .B2(n_1210), .Y(n_1209) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_51), .A2(n_345), .B1(n_718), .B2(n_721), .Y(n_1025) );
INVx1_ASAP7_75t_L g1174 ( .A(n_52), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_53), .A2(n_150), .B1(n_808), .B2(n_884), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_54), .A2(n_177), .B1(n_660), .B2(n_699), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_55), .A2(n_113), .B1(n_849), .B2(n_850), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g1260 ( .A1(n_56), .A2(n_204), .B1(n_718), .B2(n_721), .Y(n_1260) );
OA22x2_ASAP7_75t_L g672 ( .A1(n_57), .A2(n_174), .B1(n_666), .B2(n_670), .Y(n_672) );
INVx1_ASAP7_75t_L g693 ( .A(n_57), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_58), .A2(n_229), .B1(n_434), .B2(n_461), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_59), .A2(n_68), .B1(n_755), .B2(n_765), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_61), .A2(n_63), .B1(n_849), .B2(n_850), .Y(n_1083) );
AOI22xp5_ASAP7_75t_L g1078 ( .A1(n_62), .A2(n_322), .B1(n_880), .B2(n_962), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1247 ( .A1(n_64), .A2(n_387), .B1(n_955), .B2(n_988), .Y(n_1247) );
AOI22xp33_ASAP7_75t_L g1205 ( .A1(n_65), .A2(n_281), .B1(n_699), .B2(n_924), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_66), .A2(n_206), .B1(n_418), .B2(n_440), .Y(n_451) );
XNOR2x2_ASAP7_75t_L g859 ( .A(n_67), .B(n_860), .Y(n_859) );
XOR2x2_ASAP7_75t_L g1020 ( .A(n_69), .B(n_1021), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_70), .A2(n_276), .B1(n_837), .B2(n_838), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_71), .A2(n_328), .B1(n_849), .B2(n_850), .Y(n_1309) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_72), .A2(n_284), .B1(n_964), .B2(n_1157), .Y(n_1204) );
INVx1_ASAP7_75t_L g981 ( .A(n_73), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_74), .A2(n_112), .B1(n_880), .B2(n_1157), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1307 ( .A1(n_75), .A2(n_286), .B1(n_834), .B2(n_856), .Y(n_1307) );
AOI221xp5_ASAP7_75t_L g1073 ( .A1(n_77), .A2(n_199), .B1(n_914), .B2(n_943), .C(n_1074), .Y(n_1073) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_78), .B(n_194), .Y(n_652) );
INVx1_ASAP7_75t_L g669 ( .A(n_78), .Y(n_669) );
OAI21xp33_ASAP7_75t_L g694 ( .A1(n_78), .A2(n_174), .B(n_695), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g904 ( .A1(n_79), .A2(n_905), .B(n_906), .Y(n_904) );
AO221x2_ASAP7_75t_L g432 ( .A1(n_80), .A2(n_371), .B1(n_418), .B2(n_424), .C(n_433), .Y(n_432) );
AOI22xp33_ASAP7_75t_SL g874 ( .A1(n_81), .A2(n_161), .B1(n_822), .B2(n_875), .Y(n_874) );
AOI221xp5_ASAP7_75t_L g1066 ( .A1(n_82), .A2(n_341), .B1(n_905), .B2(n_1067), .C(n_1068), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_83), .A2(n_382), .B1(n_849), .B2(n_850), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_84), .A2(n_325), .B1(n_835), .B2(n_837), .Y(n_1232) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_85), .A2(n_131), .B1(n_898), .B2(n_1029), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_86), .A2(n_302), .B1(n_718), .B2(n_721), .Y(n_899) );
INVx1_ASAP7_75t_L g1305 ( .A(n_87), .Y(n_1305) );
AOI22xp5_ASAP7_75t_L g1155 ( .A1(n_88), .A2(n_197), .B1(n_801), .B2(n_1057), .Y(n_1155) );
AOI22xp33_ASAP7_75t_SL g900 ( .A1(n_89), .A2(n_230), .B1(n_801), .B2(n_882), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_90), .A2(n_363), .B1(n_911), .B2(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1213 ( .A(n_91), .Y(n_1213) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_92), .A2(n_360), .B1(n_438), .B2(n_440), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_93), .A2(n_134), .B1(n_698), .B2(n_703), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_94), .A2(n_375), .B1(n_427), .B2(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_95), .B(n_988), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_96), .A2(n_376), .B1(n_741), .B2(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g423 ( .A(n_97), .Y(n_423) );
AND2x4_ASAP7_75t_L g428 ( .A(n_97), .B(n_298), .Y(n_428) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_97), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_98), .A2(n_346), .B1(n_834), .B2(n_856), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_99), .A2(n_260), .B1(n_806), .B2(n_882), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_100), .A2(n_220), .B1(n_1005), .B2(n_1108), .Y(n_1107) );
AO22x1_ASAP7_75t_L g433 ( .A1(n_102), .A2(n_205), .B1(n_434), .B2(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g1251 ( .A(n_102), .Y(n_1251) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_104), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g892 ( .A1(n_105), .A2(n_106), .B1(n_893), .B2(n_894), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_108), .A2(n_211), .B1(n_838), .B2(n_1003), .Y(n_1231) );
INVx1_ASAP7_75t_L g1340 ( .A(n_109), .Y(n_1340) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_110), .A2(n_147), .B1(n_429), .B2(n_442), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g1248 ( .A1(n_111), .A2(n_114), .B1(n_741), .B2(n_1226), .C(n_1249), .Y(n_1248) );
XNOR2x1_ASAP7_75t_L g976 ( .A(n_117), .B(n_977), .Y(n_976) );
AOI21xp5_ASAP7_75t_L g1225 ( .A1(n_118), .A2(n_1226), .B(n_1228), .Y(n_1225) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_119), .A2(n_352), .B1(n_852), .B2(n_853), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_120), .B(n_1148), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_121), .A2(n_163), .B1(n_878), .B2(n_1318), .Y(n_1317) );
AOI21xp5_ASAP7_75t_L g1264 ( .A1(n_122), .A2(n_1265), .B(n_1266), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_123), .A2(n_164), .B1(n_808), .B2(n_809), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g1112 ( .A1(n_124), .A2(n_155), .B1(n_1113), .B2(n_1114), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1302 ( .A1(n_125), .A2(n_193), .B1(n_835), .B2(n_838), .Y(n_1302) );
INVx1_ASAP7_75t_L g1250 ( .A(n_126), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_127), .A2(n_148), .B1(n_686), .B2(n_1024), .Y(n_1201) );
INVx1_ASAP7_75t_L g421 ( .A(n_128), .Y(n_421) );
AND2x4_ASAP7_75t_L g425 ( .A(n_128), .B(n_420), .Y(n_425) );
INVx1_ASAP7_75t_SL g439 ( .A(n_128), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_129), .A2(n_282), .B1(n_746), .B2(n_1003), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_130), .A2(n_188), .B1(n_1179), .B2(n_1181), .Y(n_1178) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_132), .A2(n_207), .B1(n_871), .B2(n_872), .Y(n_870) );
XNOR2x1_ASAP7_75t_L g920 ( .A(n_133), .B(n_921), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_135), .A2(n_305), .B1(n_721), .B2(n_1111), .Y(n_1110) );
INVx1_ASAP7_75t_L g1013 ( .A(n_136), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_137), .A2(n_170), .B1(n_427), .B2(n_435), .Y(n_450) );
INVx1_ASAP7_75t_L g824 ( .A(n_138), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_139), .B(n_1067), .Y(n_1214) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_140), .A2(n_290), .B1(n_808), .B2(n_924), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g1301 ( .A1(n_141), .A2(n_386), .B1(n_837), .B2(n_852), .Y(n_1301) );
AOI221xp5_ASAP7_75t_L g940 ( .A1(n_143), .A2(n_393), .B1(n_941), .B2(n_943), .C(n_944), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_144), .A2(n_775), .B1(n_776), .B2(n_777), .Y(n_774) );
CKINVDCx5p33_ASAP7_75t_R g777 ( .A(n_144), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_145), .A2(n_159), .B1(n_805), .B2(n_880), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_146), .A2(n_311), .B1(n_746), .B2(n_951), .Y(n_950) );
XNOR2x1_ASAP7_75t_L g1217 ( .A(n_147), .B(n_1218), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g1289 ( .A1(n_149), .A2(n_215), .B1(n_875), .B2(n_905), .Y(n_1289) );
INVx1_ASAP7_75t_L g1224 ( .A(n_151), .Y(n_1224) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_152), .A2(n_191), .B1(n_846), .B2(n_855), .Y(n_1011) );
AOI22xp5_ASAP7_75t_L g1007 ( .A1(n_153), .A2(n_392), .B1(n_849), .B2(n_850), .Y(n_1007) );
AOI21xp5_ASAP7_75t_L g1150 ( .A1(n_154), .A2(n_905), .B(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g932 ( .A(n_156), .Y(n_932) );
AOI22xp5_ASAP7_75t_L g1164 ( .A1(n_158), .A2(n_185), .B1(n_721), .B2(n_1165), .Y(n_1164) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_165), .A2(n_238), .B1(n_875), .B2(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g1069 ( .A(n_166), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_167), .A2(n_250), .B1(n_735), .B2(n_1065), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_169), .A2(n_327), .B1(n_798), .B2(n_799), .Y(n_797) );
INVx1_ASAP7_75t_L g1273 ( .A(n_170), .Y(n_1273) );
AOI22xp5_ASAP7_75t_L g1008 ( .A1(n_171), .A2(n_378), .B1(n_834), .B2(n_856), .Y(n_1008) );
INVx1_ASAP7_75t_L g684 ( .A(n_172), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_172), .B(n_235), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_172), .B(n_691), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_173), .A2(n_245), .B1(n_458), .B2(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_174), .B(n_310), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g965 ( .A1(n_175), .A2(n_249), .B1(n_799), .B2(n_878), .Y(n_965) );
INVx1_ASAP7_75t_L g907 ( .A(n_178), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_180), .A2(n_280), .B1(n_869), .B2(n_988), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_181), .A2(n_189), .B1(n_812), .B2(n_813), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_182), .A2(n_335), .B1(n_799), .B2(n_878), .Y(n_877) );
AOI221xp5_ASAP7_75t_L g995 ( .A1(n_183), .A2(n_195), .B1(n_741), .B2(n_818), .C(n_996), .Y(n_995) );
AOI22xp5_ASAP7_75t_L g1243 ( .A1(n_184), .A2(n_262), .B1(n_799), .B2(n_878), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1326 ( .A1(n_186), .A2(n_340), .B1(n_659), .B2(n_1327), .Y(n_1326) );
INVx1_ASAP7_75t_L g1152 ( .A(n_187), .Y(n_1152) );
AOI21xp5_ASAP7_75t_L g1127 ( .A1(n_190), .A2(n_832), .B(n_1128), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1287 ( .A(n_192), .B(n_1288), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_194), .B(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_196), .A2(n_227), .B1(n_699), .B2(n_924), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_198), .A2(n_404), .B1(n_799), .B2(n_878), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_200), .A2(n_405), .B1(n_799), .B2(n_893), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_201), .A2(n_248), .B1(n_660), .B2(n_882), .Y(n_881) );
AO22x2_ASAP7_75t_L g1121 ( .A1(n_202), .A2(n_1122), .B1(n_1140), .B2(n_1141), .Y(n_1121) );
INVxp67_ASAP7_75t_SL g1140 ( .A(n_202), .Y(n_1140) );
INVx1_ASAP7_75t_L g1229 ( .A(n_203), .Y(n_1229) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_208), .A2(n_326), .B1(n_808), .B2(n_884), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_210), .B(n_867), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_213), .A2(n_380), .B1(n_812), .B2(n_1065), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_214), .A2(n_219), .B1(n_926), .B2(n_1057), .Y(n_1056) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_217), .A2(n_794), .B1(n_795), .B2(n_827), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_217), .Y(n_794) );
AOI21xp33_ASAP7_75t_L g1211 ( .A1(n_218), .A2(n_1003), .B(n_1212), .Y(n_1211) );
AOI22xp33_ASAP7_75t_L g1290 ( .A1(n_221), .A2(n_253), .B1(n_741), .B2(n_911), .Y(n_1290) );
AOI22xp33_ASAP7_75t_L g1284 ( .A1(n_223), .A2(n_400), .B1(n_798), .B2(n_799), .Y(n_1284) );
AOI22xp33_ASAP7_75t_L g1332 ( .A1(n_224), .A2(n_394), .B1(n_1333), .B2(n_1334), .Y(n_1332) );
BUFx2_ASAP7_75t_L g1130 ( .A(n_225), .Y(n_1130) );
XNOR2x1_ASAP7_75t_L g947 ( .A(n_226), .B(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g1170 ( .A(n_228), .Y(n_1170) );
INVx1_ASAP7_75t_L g997 ( .A(n_231), .Y(n_997) );
AOI22xp5_ASAP7_75t_L g1221 ( .A1(n_232), .A2(n_377), .B1(n_699), .B2(n_1222), .Y(n_1221) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_233), .A2(n_255), .B1(n_418), .B2(n_424), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_234), .A2(n_406), .B1(n_905), .B2(n_1032), .Y(n_1031) );
INVx1_ASAP7_75t_L g667 ( .A(n_235), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_236), .A2(n_273), .B1(n_898), .B2(n_1029), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g1202 ( .A1(n_237), .A2(n_366), .B1(n_1184), .B2(n_1203), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_240), .A2(n_342), .B1(n_418), .B2(n_440), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_241), .A2(n_399), .B1(n_707), .B2(n_713), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g1261 ( .A1(n_242), .A2(n_272), .B1(n_713), .B2(n_893), .Y(n_1261) );
XNOR2x1_ASAP7_75t_L g828 ( .A(n_243), .B(n_829), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_244), .A2(n_373), .B1(n_916), .B2(n_917), .Y(n_915) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_246), .A2(n_288), .B1(n_418), .B2(n_440), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_247), .A2(n_343), .B1(n_808), .B2(n_1061), .Y(n_1060) );
AOI22xp5_ASAP7_75t_L g1004 ( .A1(n_251), .A2(n_261), .B1(n_875), .B2(n_1005), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_252), .B(n_832), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_254), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_257), .A2(n_338), .B1(n_418), .B2(n_458), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_258), .A2(n_333), .B1(n_434), .B2(n_435), .Y(n_454) );
OR2x2_ASAP7_75t_L g1206 ( .A(n_258), .B(n_1207), .Y(n_1206) );
INVxp67_ASAP7_75t_L g1216 ( .A(n_258), .Y(n_1216) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_259), .A2(n_319), .B1(n_718), .B2(n_884), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1285 ( .A1(n_263), .A2(n_313), .B1(n_699), .B2(n_809), .Y(n_1285) );
AOI22xp5_ASAP7_75t_L g1077 ( .A1(n_264), .A2(n_285), .B1(n_846), .B2(n_855), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_265), .A2(n_337), .B1(n_801), .B2(n_802), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_266), .A2(n_318), .B1(n_847), .B2(n_853), .Y(n_928) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_268), .A2(n_368), .B1(n_427), .B2(n_429), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g1055 ( .A1(n_269), .A2(n_270), .B1(n_713), .B2(n_878), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_271), .A2(n_347), .B1(n_905), .B2(n_1103), .Y(n_1102) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_274), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_275), .A2(n_316), .B1(n_837), .B2(n_838), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g1291 ( .A1(n_277), .A2(n_308), .B1(n_813), .B2(n_1292), .Y(n_1291) );
AOI22xp5_ASAP7_75t_L g1182 ( .A1(n_278), .A2(n_348), .B1(n_707), .B2(n_1183), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_279), .A2(n_385), .B1(n_802), .B2(n_926), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_289), .B(n_1269), .Y(n_1268) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_291), .A2(n_398), .B1(n_1100), .B2(n_1101), .Y(n_1099) );
AOI221xp5_ASAP7_75t_L g1335 ( .A1(n_292), .A2(n_294), .B1(n_1005), .B2(n_1336), .C(n_1339), .Y(n_1335) );
INVx1_ASAP7_75t_L g1043 ( .A(n_293), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_295), .A2(n_330), .B1(n_846), .B2(n_847), .Y(n_845) );
INVx1_ASAP7_75t_L g939 ( .A(n_296), .Y(n_939) );
AOI22x1_ASAP7_75t_L g1051 ( .A1(n_297), .A2(n_1052), .B1(n_1053), .B2(n_1070), .Y(n_1051) );
INVx1_ASAP7_75t_L g1070 ( .A(n_297), .Y(n_1070) );
AND2x4_ASAP7_75t_L g422 ( .A(n_298), .B(n_423), .Y(n_422) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_298), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_299), .B(n_818), .Y(n_817) );
XNOR2x2_ASAP7_75t_L g1314 ( .A(n_301), .B(n_1315), .Y(n_1314) );
AOI22xp33_ASAP7_75t_L g1310 ( .A1(n_303), .A2(n_334), .B1(n_846), .B2(n_855), .Y(n_1310) );
INVx1_ASAP7_75t_L g983 ( .A(n_304), .Y(n_983) );
XOR2x2_ASAP7_75t_L g1161 ( .A(n_306), .B(n_1162), .Y(n_1161) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_307), .A2(n_359), .B1(n_835), .B2(n_852), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_309), .A2(n_324), .B1(n_718), .B2(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g682 ( .A(n_310), .Y(n_682) );
INVxp67_ASAP7_75t_L g764 ( .A(n_310), .Y(n_764) );
AOI21xp33_ASAP7_75t_SL g1124 ( .A1(n_312), .A2(n_1003), .B(n_1125), .Y(n_1124) );
INVx1_ASAP7_75t_L g1075 ( .A(n_314), .Y(n_1075) );
INVx1_ASAP7_75t_L g1017 ( .A(n_315), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1308 ( .A1(n_317), .A2(n_336), .B1(n_847), .B2(n_853), .Y(n_1308) );
INVx2_ASAP7_75t_L g420 ( .A(n_320), .Y(n_420) );
INVx1_ASAP7_75t_L g1172 ( .A(n_321), .Y(n_1172) );
AOI21xp5_ASAP7_75t_L g862 ( .A1(n_323), .A2(n_863), .B(n_864), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g833 ( .A1(n_331), .A2(n_332), .B1(n_834), .B2(n_835), .Y(n_833) );
INVx1_ASAP7_75t_L g1187 ( .A(n_339), .Y(n_1187) );
INVx1_ASAP7_75t_L g1175 ( .A(n_344), .Y(n_1175) );
INVx1_ASAP7_75t_L g945 ( .A(n_349), .Y(n_945) );
INVx1_ASAP7_75t_L g1126 ( .A(n_350), .Y(n_1126) );
AOI21xp33_ASAP7_75t_L g839 ( .A1(n_353), .A2(n_840), .B(n_841), .Y(n_839) );
INVx1_ASAP7_75t_L g842 ( .A(n_354), .Y(n_842) );
INVx1_ASAP7_75t_L g985 ( .A(n_355), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_356), .B(n_1105), .Y(n_1104) );
AOI21xp33_ASAP7_75t_L g954 ( .A1(n_357), .A2(n_955), .B(n_956), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_358), .A2(n_361), .B1(n_686), .B2(n_926), .Y(n_967) );
INVx1_ASAP7_75t_L g1143 ( .A(n_362), .Y(n_1143) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_364), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_365), .B(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g1296 ( .A(n_368), .Y(n_1296) );
XNOR2x2_ASAP7_75t_L g656 ( .A(n_370), .B(n_657), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_370), .A2(n_773), .B1(n_778), .B2(n_780), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_372), .A2(n_389), .B1(n_718), .B2(n_721), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_374), .A2(n_396), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
INVx1_ASAP7_75t_SL g1293 ( .A(n_375), .Y(n_1293) );
INVx1_ASAP7_75t_L g1018 ( .A(n_379), .Y(n_1018) );
BUFx2_ASAP7_75t_L g1132 ( .A(n_381), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_383), .B(n_1300), .Y(n_1299) );
AOI22xp33_ASAP7_75t_L g1259 ( .A1(n_384), .A2(n_401), .B1(n_660), .B2(n_882), .Y(n_1259) );
AOI21xp5_ASAP7_75t_L g1015 ( .A1(n_388), .A2(n_942), .B(n_1016), .Y(n_1015) );
INVx1_ASAP7_75t_L g865 ( .A(n_391), .Y(n_865) );
AOI21xp33_ASAP7_75t_L g1303 ( .A1(n_395), .A2(n_840), .B(n_1304), .Y(n_1303) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_397), .Y(n_726) );
AOI21xp33_ASAP7_75t_SL g821 ( .A1(n_402), .A2(n_822), .B(n_823), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_1191), .B1(n_1344), .B2(n_1346), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_785), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_409), .B(n_1347), .Y(n_1346) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI221xp5_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_642), .B1(n_644), .B2(n_655), .C(n_772), .Y(n_410) );
AND5x1_ASAP7_75t_L g411 ( .A(n_412), .B(n_604), .C(n_613), .D(n_628), .E(n_638), .Y(n_411) );
OAI33xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_507), .A3(n_533), .B1(n_557), .B2(n_572), .B3(n_581), .Y(n_412) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_481), .C(n_492), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_443), .B1(n_462), .B2(n_468), .C(n_471), .Y(n_414) );
INVx1_ASAP7_75t_L g597 ( .A(n_415), .Y(n_597) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_430), .Y(n_415) );
AND2x2_ASAP7_75t_L g478 ( .A(n_416), .B(n_463), .Y(n_478) );
CKINVDCx6p67_ASAP7_75t_R g491 ( .A(n_416), .Y(n_491) );
AND2x2_ASAP7_75t_L g504 ( .A(n_416), .B(n_476), .Y(n_504) );
AND2x2_ASAP7_75t_L g513 ( .A(n_416), .B(n_486), .Y(n_513) );
AND2x2_ASAP7_75t_L g523 ( .A(n_416), .B(n_436), .Y(n_523) );
AND2x2_ASAP7_75t_L g545 ( .A(n_416), .B(n_517), .Y(n_545) );
AND2x2_ASAP7_75t_L g576 ( .A(n_416), .B(n_485), .Y(n_576) );
AND2x2_ASAP7_75t_L g584 ( .A(n_416), .B(n_537), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_416), .B(n_495), .Y(n_587) );
OAI332xp33_ASAP7_75t_L g589 ( .A1(n_416), .A2(n_470), .A3(n_491), .B1(n_590), .B2(n_591), .B3(n_592), .C1(n_594), .C2(n_595), .Y(n_589) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_426), .Y(n_416) );
INVx3_ASAP7_75t_L g555 ( .A(n_418), .Y(n_555) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_422), .Y(n_418) );
AND2x2_ASAP7_75t_L g427 ( .A(n_419), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g434 ( .A(n_419), .B(n_428), .Y(n_434) );
AND2x2_ASAP7_75t_L g442 ( .A(n_419), .B(n_428), .Y(n_442) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
AND3x4_ASAP7_75t_L g438 ( .A(n_420), .B(n_422), .C(n_439), .Y(n_438) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_420), .Y(n_654) );
AND2x4_ASAP7_75t_L g424 ( .A(n_422), .B(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_L g440 ( .A(n_422), .B(n_425), .Y(n_440) );
AND2x2_ASAP7_75t_L g429 ( .A(n_425), .B(n_428), .Y(n_429) );
AND2x2_ASAP7_75t_L g435 ( .A(n_425), .B(n_428), .Y(n_435) );
AND2x4_ASAP7_75t_L g461 ( .A(n_425), .B(n_428), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_430), .B(n_496), .Y(n_531) );
AND2x2_ASAP7_75t_L g550 ( .A(n_430), .B(n_490), .Y(n_550) );
NAND3xp33_ASAP7_75t_L g569 ( .A(n_430), .B(n_548), .C(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g621 ( .A(n_430), .B(n_478), .Y(n_621) );
AND2x2_ASAP7_75t_L g630 ( .A(n_430), .B(n_491), .Y(n_630) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NOR2x1_ASAP7_75t_L g462 ( .A(n_431), .B(n_463), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_431), .B(n_543), .Y(n_599) );
OR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_436), .Y(n_431) );
AND2x2_ASAP7_75t_L g476 ( .A(n_432), .B(n_436), .Y(n_476) );
AND2x2_ASAP7_75t_L g485 ( .A(n_432), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g495 ( .A(n_432), .Y(n_495) );
AND2x2_ASAP7_75t_L g627 ( .A(n_432), .B(n_491), .Y(n_627) );
BUFx2_ASAP7_75t_L g643 ( .A(n_434), .Y(n_643) );
INVx1_ASAP7_75t_L g486 ( .A(n_436), .Y(n_486) );
AND2x2_ASAP7_75t_L g517 ( .A(n_436), .B(n_495), .Y(n_517) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_441), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g784 ( .A1(n_439), .A2(n_648), .B(n_653), .Y(n_784) );
INVx2_ASAP7_75t_SL g459 ( .A(n_440), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_452), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_444), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_446), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_446), .B(n_543), .Y(n_637) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g502 ( .A(n_447), .Y(n_502) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g469 ( .A(n_448), .Y(n_469) );
OR2x2_ASAP7_75t_L g526 ( .A(n_448), .B(n_480), .Y(n_526) );
INVx4_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g498 ( .A(n_449), .B(n_480), .Y(n_498) );
AND2x2_ASAP7_75t_L g535 ( .A(n_449), .B(n_480), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_449), .B(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g564 ( .A(n_449), .B(n_453), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_449), .B(n_543), .Y(n_570) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
AOI222xp33_ASAP7_75t_L g518 ( .A1(n_452), .A2(n_519), .B1(n_524), .B2(n_527), .C1(n_528), .C2(n_529), .Y(n_518) );
AOI211xp5_ASAP7_75t_L g567 ( .A1(n_452), .A2(n_511), .B(n_568), .C(n_571), .Y(n_567) );
AND2x2_ASAP7_75t_L g588 ( .A(n_452), .B(n_528), .Y(n_588) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .Y(n_452) );
INVx2_ASAP7_75t_L g480 ( .A(n_453), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
INVx4_ASAP7_75t_L g470 ( .A(n_456), .Y(n_470) );
INVx1_ASAP7_75t_L g506 ( .A(n_456), .Y(n_506) );
AND2x2_ASAP7_75t_L g549 ( .A(n_456), .B(n_525), .Y(n_549) );
AND2x2_ASAP7_75t_L g577 ( .A(n_456), .B(n_469), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_456), .B(n_502), .Y(n_600) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_460), .Y(n_456) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_462), .B(n_491), .Y(n_566) );
AND2x2_ASAP7_75t_L g514 ( .A(n_463), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_463), .B(n_497), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_463), .B(n_517), .Y(n_595) );
INVx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g496 ( .A(n_464), .B(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g537 ( .A(n_464), .B(n_476), .Y(n_537) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g474 ( .A(n_465), .Y(n_474) );
AND2x2_ASAP7_75t_L g490 ( .A(n_465), .B(n_491), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_465), .B(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g543 ( .A(n_465), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_465), .B(n_470), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_465), .B(n_535), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_465), .B(n_513), .Y(n_619) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g594 ( .A(n_468), .Y(n_594) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_469), .A2(n_472), .B(n_477), .C(n_479), .Y(n_471) );
AND2x2_ASAP7_75t_L g484 ( .A(n_470), .B(n_480), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_470), .B(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g547 ( .A(n_470), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_470), .B(n_497), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g616 ( .A1(n_470), .A2(n_617), .B(n_620), .C(n_622), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_470), .B(n_564), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g638 ( .A1(n_470), .A2(n_523), .B(n_639), .C(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_473), .B(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_474), .A2(n_484), .B(n_509), .C(n_514), .Y(n_508) );
AND2x2_ASAP7_75t_L g524 ( .A(n_474), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_474), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g575 ( .A(n_474), .B(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_474), .B(n_608), .Y(n_607) );
O2A1O1Ixp33_ASAP7_75t_SL g611 ( .A1(n_474), .A2(n_483), .B(n_530), .C(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_476), .B(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g511 ( .A(n_476), .B(n_491), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_476), .B(n_490), .Y(n_633) );
INVx1_ASAP7_75t_L g527 ( .A(n_477), .Y(n_527) );
INVx3_ASAP7_75t_SL g505 ( .A(n_479), .Y(n_505) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_L g548 ( .A(n_480), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_485), .B(n_487), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g573 ( .A(n_484), .Y(n_573) );
AND2x2_ASAP7_75t_L g489 ( .A(n_485), .B(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g521 ( .A(n_485), .B(n_491), .Y(n_521) );
INVx1_ASAP7_75t_L g530 ( .A(n_485), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_486), .B(n_491), .Y(n_561) );
AOI211xp5_ASAP7_75t_L g604 ( .A1(n_487), .A2(n_525), .B(n_605), .C(n_611), .Y(n_604) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_491), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_491), .B(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_491), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_491), .B(n_543), .Y(n_624) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_496), .B(n_499), .C(n_506), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_494), .B(n_603), .Y(n_602) );
OAI22xp33_ASAP7_75t_L g631 ( .A1(n_494), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_496), .B(n_513), .Y(n_532) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AOI21xp33_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_503), .B(n_505), .Y(n_499) );
INVxp67_ASAP7_75t_SL g614 ( .A(n_500), .Y(n_614) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_504), .B(n_525), .Y(n_641) );
INVx1_ASAP7_75t_L g582 ( .A(n_505), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_505), .B(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_506), .B(n_540), .Y(n_539) );
NAND4xp25_ASAP7_75t_SL g507 ( .A(n_508), .B(n_518), .C(n_531), .D(n_532), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_510), .B(n_512), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_514), .A2(n_535), .B1(n_629), .B2(n_630), .C(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_516), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g593 ( .A(n_517), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_520), .B(n_522), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_521), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g580 ( .A(n_524), .Y(n_580) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_528), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g609 ( .A(n_529), .Y(n_609) );
AND2x2_ASAP7_75t_L g592 ( .A(n_530), .B(n_593), .Y(n_592) );
OAI211xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_536), .B(n_538), .C(n_544), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OAI211xp5_ASAP7_75t_L g622 ( .A1(n_537), .A2(n_623), .B(n_625), .C(n_626), .Y(n_622) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI211xp5_ASAP7_75t_L g572 ( .A1(n_540), .A2(n_573), .B(n_574), .C(n_578), .Y(n_572) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp33_ASAP7_75t_L g546 ( .A(n_542), .B(n_547), .Y(n_546) );
AOI221xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .B1(n_549), .B2(n_550), .C(n_551), .Y(n_544) );
INVx1_ASAP7_75t_L g608 ( .A(n_545), .Y(n_608) );
INVx1_ASAP7_75t_L g615 ( .A(n_547), .Y(n_615) );
INVx1_ASAP7_75t_L g610 ( .A(n_549), .Y(n_610) );
INVx2_ASAP7_75t_L g571 ( .A(n_551), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_556), .Y(n_552) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OAI211xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B(n_562), .C(n_567), .Y(n_557) );
INVx1_ASAP7_75t_L g629 ( .A(n_558), .Y(n_629) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OAI21xp5_ASAP7_75t_SL g574 ( .A1(n_565), .A2(n_575), .B(n_577), .Y(n_574) );
O2A1O1Ixp33_ASAP7_75t_L g613 ( .A1(n_565), .A2(n_614), .B(n_615), .C(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVxp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_573), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g612 ( .A(n_576), .Y(n_612) );
INVxp67_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
OAI211xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .B(n_585), .C(n_601), .Y(n_581) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI211xp5_ASAP7_75t_SL g585 ( .A1(n_586), .A2(n_588), .B(n_589), .C(n_596), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g632 ( .A(n_588), .Y(n_632) );
INVx1_ASAP7_75t_L g639 ( .A(n_590), .Y(n_639) );
AOI21xp33_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_598), .B(n_600), .Y(n_596) );
INVxp33_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
AOI21xp33_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_609), .B(n_610), .Y(n_605) );
INVxp33_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVxp67_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
INVxp67_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVxp33_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVxp33_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVxp67_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g642 ( .A(n_643), .Y(n_642) );
CKINVDCx16_ASAP7_75t_R g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_653), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
AND2x2_ASAP7_75t_L g779 ( .A(n_647), .B(n_653), .Y(n_779) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g787 ( .A(n_648), .B(n_649), .C(n_653), .Y(n_787) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AO21x2_ASAP7_75t_L g768 ( .A1(n_650), .A2(n_769), .B(n_770), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AO21x1_ASAP7_75t_L g781 ( .A1(n_654), .A2(n_782), .B(n_784), .Y(n_781) );
BUFx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_657), .Y(n_776) );
NAND3xp33_ASAP7_75t_SL g657 ( .A(n_658), .B(n_696), .C(n_724), .Y(n_657) );
BUFx3_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx6f_ASAP7_75t_L g801 ( .A(n_661), .Y(n_801) );
BUFx6f_ASAP7_75t_L g926 ( .A(n_661), .Y(n_926) );
BUFx6f_ASAP7_75t_L g1024 ( .A(n_661), .Y(n_1024) );
AND2x4_ASAP7_75t_L g661 ( .A(n_662), .B(n_673), .Y(n_661) );
AND2x4_ASAP7_75t_L g700 ( .A(n_662), .B(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g710 ( .A(n_662), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g714 ( .A(n_662), .B(n_715), .Y(n_714) );
AND2x4_ASAP7_75t_L g834 ( .A(n_662), .B(n_723), .Y(n_834) );
AND2x4_ASAP7_75t_L g846 ( .A(n_662), .B(n_701), .Y(n_846) );
AND2x4_ASAP7_75t_L g849 ( .A(n_662), .B(n_711), .Y(n_849) );
AND2x4_ASAP7_75t_L g850 ( .A(n_662), .B(n_715), .Y(n_850) );
AND2x4_ASAP7_75t_L g662 ( .A(n_663), .B(n_671), .Y(n_662) );
AND2x2_ASAP7_75t_L g731 ( .A(n_663), .B(n_672), .Y(n_731) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g720 ( .A(n_664), .B(n_672), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_668), .Y(n_664) );
NAND2xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
INVx2_ASAP7_75t_L g670 ( .A(n_666), .Y(n_670) );
INVx3_ASAP7_75t_L g677 ( .A(n_666), .Y(n_677) );
NAND2xp33_ASAP7_75t_L g683 ( .A(n_666), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g695 ( .A(n_666), .Y(n_695) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_666), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_667), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
OAI21xp5_ASAP7_75t_L g763 ( .A1(n_669), .A2(n_695), .B(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g762 ( .A(n_672), .B(n_763), .Y(n_762) );
AND2x4_ASAP7_75t_L g688 ( .A(n_673), .B(n_689), .Y(n_688) );
AND2x4_ASAP7_75t_L g847 ( .A(n_673), .B(n_720), .Y(n_847) );
AND2x4_ASAP7_75t_L g856 ( .A(n_673), .B(n_689), .Y(n_856) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g723 ( .A(n_674), .Y(n_723) );
OR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_679), .Y(n_674) );
AND2x4_ASAP7_75t_L g701 ( .A(n_675), .B(n_702), .Y(n_701) );
AND2x4_ASAP7_75t_L g711 ( .A(n_675), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g716 ( .A(n_675), .Y(n_716) );
AND2x2_ASAP7_75t_L g758 ( .A(n_675), .B(n_759), .Y(n_758) );
AND2x4_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_677), .B(n_682), .Y(n_681) );
INVxp67_ASAP7_75t_L g691 ( .A(n_677), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g770 ( .A(n_678), .B(n_690), .C(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g702 ( .A(n_679), .Y(n_702) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g712 ( .A(n_680), .Y(n_712) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .Y(n_680) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx5_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx3_ASAP7_75t_L g802 ( .A(n_687), .Y(n_802) );
INVx2_ASAP7_75t_L g1057 ( .A(n_687), .Y(n_1057) );
INVx1_ASAP7_75t_L g1111 ( .A(n_687), .Y(n_1111) );
INVx6_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
BUFx12f_ASAP7_75t_L g882 ( .A(n_688), .Y(n_882) );
AND2x4_ASAP7_75t_L g705 ( .A(n_689), .B(n_701), .Y(n_705) );
AND2x4_ASAP7_75t_L g747 ( .A(n_689), .B(n_715), .Y(n_747) );
AND2x4_ASAP7_75t_L g835 ( .A(n_689), .B(n_715), .Y(n_835) );
AND2x4_ASAP7_75t_L g855 ( .A(n_689), .B(n_701), .Y(n_855) );
AND2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_694), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
AND3x1_ASAP7_75t_L g696 ( .A(n_697), .B(n_706), .C(n_717), .Y(n_696) );
BUFx12f_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
BUFx6f_ASAP7_75t_L g1113 ( .A(n_699), .Y(n_1113) );
INVx1_ASAP7_75t_L g1180 ( .A(n_699), .Y(n_1180) );
BUFx12f_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
BUFx6f_ASAP7_75t_L g808 ( .A(n_700), .Y(n_808) );
BUFx6f_ASAP7_75t_L g898 ( .A(n_700), .Y(n_898) );
AND2x2_ASAP7_75t_L g719 ( .A(n_701), .B(n_720), .Y(n_719) );
AND2x4_ASAP7_75t_L g853 ( .A(n_701), .B(n_720), .Y(n_853) );
AND2x2_ASAP7_75t_L g963 ( .A(n_701), .B(n_720), .Y(n_963) );
INVx4_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g809 ( .A(n_704), .Y(n_809) );
INVx4_ASAP7_75t_L g884 ( .A(n_704), .Y(n_884) );
INVx2_ASAP7_75t_L g924 ( .A(n_704), .Y(n_924) );
INVx1_ASAP7_75t_L g1029 ( .A(n_704), .Y(n_1029) );
INVx4_ASAP7_75t_L g1061 ( .A(n_704), .Y(n_1061) );
INVx1_ASAP7_75t_L g1167 ( .A(n_704), .Y(n_1167) );
INVx1_ASAP7_75t_L g1222 ( .A(n_704), .Y(n_1222) );
INVx8_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
BUFx4f_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g798 ( .A(n_709), .Y(n_798) );
INVx1_ASAP7_75t_L g1203 ( .A(n_709), .Y(n_1203) );
INVx3_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
BUFx12f_ASAP7_75t_L g878 ( .A(n_710), .Y(n_878) );
BUFx6f_ASAP7_75t_L g893 ( .A(n_710), .Y(n_893) );
AND2x4_ASAP7_75t_L g730 ( .A(n_711), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g737 ( .A(n_711), .B(n_720), .Y(n_737) );
AND2x4_ASAP7_75t_L g837 ( .A(n_711), .B(n_720), .Y(n_837) );
AND2x4_ASAP7_75t_L g852 ( .A(n_711), .B(n_731), .Y(n_852) );
AND2x4_ASAP7_75t_L g715 ( .A(n_712), .B(n_716), .Y(n_715) );
BUFx3_ASAP7_75t_L g1318 ( .A(n_713), .Y(n_1318) );
BUFx5_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
BUFx6f_ASAP7_75t_L g799 ( .A(n_714), .Y(n_799) );
INVx1_ASAP7_75t_L g896 ( .A(n_714), .Y(n_896) );
BUFx3_ASAP7_75t_L g1184 ( .A(n_714), .Y(n_1184) );
AND2x4_ASAP7_75t_L g742 ( .A(n_715), .B(n_731), .Y(n_742) );
AND2x2_ASAP7_75t_L g753 ( .A(n_715), .B(n_720), .Y(n_753) );
AND2x2_ASAP7_75t_L g840 ( .A(n_715), .B(n_731), .Y(n_840) );
AND2x2_ASAP7_75t_L g942 ( .A(n_715), .B(n_720), .Y(n_942) );
BUFx8_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
BUFx6f_ASAP7_75t_L g805 ( .A(n_719), .Y(n_805) );
AND2x4_ASAP7_75t_L g722 ( .A(n_720), .B(n_723), .Y(n_722) );
BUFx3_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
BUFx12f_ASAP7_75t_L g806 ( .A(n_722), .Y(n_806) );
BUFx6f_ASAP7_75t_L g880 ( .A(n_722), .Y(n_880) );
BUFx6f_ASAP7_75t_L g964 ( .A(n_722), .Y(n_964) );
BUFx6f_ASAP7_75t_L g1283 ( .A(n_722), .Y(n_1283) );
NOR3xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_738), .C(n_748), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B1(n_732), .B2(n_733), .Y(n_725) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g822 ( .A(n_729), .Y(n_822) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
BUFx6f_ASAP7_75t_L g905 ( .A(n_730), .Y(n_905) );
BUFx3_ASAP7_75t_L g955 ( .A(n_730), .Y(n_955) );
BUFx3_ASAP7_75t_L g1003 ( .A(n_730), .Y(n_1003) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx3_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
BUFx6f_ASAP7_75t_L g918 ( .A(n_736), .Y(n_918) );
INVx1_ASAP7_75t_L g1032 ( .A(n_736), .Y(n_1032) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
BUFx3_ASAP7_75t_L g812 ( .A(n_737), .Y(n_812) );
BUFx6f_ASAP7_75t_L g875 ( .A(n_737), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .B1(n_743), .B2(n_744), .Y(n_738) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
BUFx3_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
BUFx6f_ASAP7_75t_L g815 ( .A(n_742), .Y(n_815) );
BUFx8_ASAP7_75t_SL g871 ( .A(n_742), .Y(n_871) );
INVx2_ASAP7_75t_L g910 ( .A(n_742), .Y(n_910) );
BUFx6f_ASAP7_75t_L g951 ( .A(n_742), .Y(n_951) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
BUFx3_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx3_ASAP7_75t_L g982 ( .A(n_746), .Y(n_982) );
BUFx6f_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx3_ASAP7_75t_L g873 ( .A(n_747), .Y(n_873) );
BUFx6f_ASAP7_75t_L g911 ( .A(n_747), .Y(n_911) );
OAI21xp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B(n_754), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx3_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g914 ( .A(n_752), .Y(n_914) );
INVx2_ASAP7_75t_L g959 ( .A(n_752), .Y(n_959) );
INVx2_ASAP7_75t_L g1067 ( .A(n_752), .Y(n_1067) );
INVx2_ASAP7_75t_L g1148 ( .A(n_752), .Y(n_1148) );
INVx2_ASAP7_75t_L g1338 ( .A(n_752), .Y(n_1338) );
INVx3_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g820 ( .A(n_753), .Y(n_820) );
BUFx3_ASAP7_75t_L g832 ( .A(n_753), .Y(n_832) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx4_ASAP7_75t_L g813 ( .A(n_756), .Y(n_813) );
INVx2_ASAP7_75t_L g916 ( .A(n_756), .Y(n_916) );
INVx3_ASAP7_75t_L g1005 ( .A(n_756), .Y(n_1005) );
INVx2_ASAP7_75t_L g1065 ( .A(n_756), .Y(n_1065) );
OAI21xp5_ASAP7_75t_L g1266 ( .A1(n_756), .A2(n_1267), .B(n_1268), .Y(n_1266) );
INVx5_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
BUFx2_ASAP7_75t_L g953 ( .A(n_757), .Y(n_953) );
BUFx4f_ASAP7_75t_L g988 ( .A(n_757), .Y(n_988) );
BUFx2_ASAP7_75t_L g1210 ( .A(n_757), .Y(n_1210) );
AND2x4_ASAP7_75t_L g757 ( .A(n_758), .B(n_762), .Y(n_757) );
AND2x2_ASAP7_75t_L g838 ( .A(n_758), .B(n_762), .Y(n_838) );
AND2x4_ASAP7_75t_L g867 ( .A(n_758), .B(n_762), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVx1_ASAP7_75t_L g769 ( .A(n_760), .Y(n_769) );
INVx4_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g906 ( .A(n_766), .B(n_907), .Y(n_906) );
NOR2xp33_ASAP7_75t_L g956 ( .A(n_766), .B(n_957), .Y(n_956) );
NOR2xp33_ASAP7_75t_L g1016 ( .A(n_766), .B(n_1017), .Y(n_1016) );
NOR2xp33_ASAP7_75t_L g1125 ( .A(n_766), .B(n_1126), .Y(n_1125) );
NOR2xp33_ASAP7_75t_L g1249 ( .A(n_766), .B(n_1250), .Y(n_1249) );
NOR2xp33_ASAP7_75t_L g1339 ( .A(n_766), .B(n_1340), .Y(n_1339) );
INVx3_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx4_ASAP7_75t_L g843 ( .A(n_767), .Y(n_843) );
INVx3_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
BUFx6f_ASAP7_75t_L g826 ( .A(n_768), .Y(n_826) );
INVxp33_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
BUFx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
BUFx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_783), .Y(n_782) );
NAND3xp33_ASAP7_75t_SL g785 ( .A(n_786), .B(n_788), .C(n_972), .Y(n_785) );
INVx1_ASAP7_75t_L g1192 ( .A(n_786), .Y(n_1192) );
INVx2_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
OAI32xp33_ASAP7_75t_L g1191 ( .A1(n_788), .A2(n_972), .A3(n_1192), .B1(n_1193), .B2(n_1349), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1344 ( .A1(n_788), .A2(n_789), .B1(n_972), .B2(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_791), .B1(n_857), .B2(n_971), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
XOR2x2_ASAP7_75t_L g792 ( .A(n_793), .B(n_828), .Y(n_792) );
INVx1_ASAP7_75t_L g827 ( .A(n_795), .Y(n_827) );
NAND4xp75_ASAP7_75t_L g795 ( .A(n_796), .B(n_803), .C(n_810), .D(n_816), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_797), .B(n_800), .Y(n_796) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_807), .Y(n_803) );
BUFx3_ASAP7_75t_L g1324 ( .A(n_805), .Y(n_1324) );
BUFx2_ASAP7_75t_SL g1320 ( .A(n_808), .Y(n_1320) );
AND2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_814), .Y(n_810) );
BUFx2_ASAP7_75t_L g1331 ( .A(n_812), .Y(n_1331) );
INVx2_ASAP7_75t_L g1042 ( .A(n_813), .Y(n_1042) );
BUFx3_ASAP7_75t_L g1333 ( .A(n_815), .Y(n_1333) );
AND2x2_ASAP7_75t_L g816 ( .A(n_817), .B(n_821), .Y(n_816) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g863 ( .A(n_819), .Y(n_863) );
INVx2_ASAP7_75t_L g1288 ( .A(n_819), .Y(n_1288) );
BUFx6f_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx2_ASAP7_75t_L g1300 ( .A(n_820), .Y(n_1300) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
NOR2xp33_ASAP7_75t_L g944 ( .A(n_825), .B(n_945), .Y(n_944) );
NOR2xp33_ASAP7_75t_L g1212 ( .A(n_825), .B(n_1213), .Y(n_1212) );
NOR2xp33_ASAP7_75t_L g1228 ( .A(n_825), .B(n_1229), .Y(n_1228) );
BUFx6f_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_SL g1045 ( .A(n_826), .Y(n_1045) );
BUFx6f_ASAP7_75t_L g1153 ( .A(n_826), .Y(n_1153) );
INVx1_ASAP7_75t_L g1292 ( .A(n_826), .Y(n_1292) );
OR2x2_ASAP7_75t_L g829 ( .A(n_830), .B(n_844), .Y(n_829) );
NAND4xp25_ASAP7_75t_L g830 ( .A(n_831), .B(n_833), .C(n_836), .D(n_839), .Y(n_830) );
INVx2_ASAP7_75t_L g1039 ( .A(n_832), .Y(n_1039) );
INVx1_ASAP7_75t_L g1106 ( .A(n_832), .Y(n_1106) );
BUFx3_ASAP7_75t_L g1265 ( .A(n_832), .Y(n_1265) );
INVx2_ASAP7_75t_L g938 ( .A(n_835), .Y(n_938) );
INVx1_ASAP7_75t_L g936 ( .A(n_837), .Y(n_936) );
INVx2_ASAP7_75t_L g1133 ( .A(n_837), .Y(n_1133) );
HB1xp67_ASAP7_75t_L g943 ( .A(n_840), .Y(n_943) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
INVx4_ASAP7_75t_L g869 ( .A(n_843), .Y(n_869) );
NOR2xp33_ASAP7_75t_L g1068 ( .A(n_843), .B(n_1069), .Y(n_1068) );
NOR2xp33_ASAP7_75t_L g1074 ( .A(n_843), .B(n_1075), .Y(n_1074) );
INVx1_ASAP7_75t_L g1108 ( .A(n_843), .Y(n_1108) );
NOR2xp33_ASAP7_75t_L g1304 ( .A(n_843), .B(n_1305), .Y(n_1304) );
NAND4xp25_ASAP7_75t_L g844 ( .A(n_845), .B(n_848), .C(n_851), .D(n_854), .Y(n_844) );
INVx2_ASAP7_75t_L g933 ( .A(n_852), .Y(n_933) );
INVx2_ASAP7_75t_L g971 ( .A(n_857), .Y(n_971) );
OAI22x1_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_885), .B1(n_886), .B2(n_969), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_L g970 ( .A(n_859), .Y(n_970) );
OR2x2_ASAP7_75t_L g860 ( .A(n_861), .B(n_876), .Y(n_860) );
NAND3xp33_ASAP7_75t_L g861 ( .A(n_862), .B(n_870), .C(n_874), .Y(n_861) );
OAI21xp33_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_866), .B(n_868), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g1128 ( .A1(n_866), .A2(n_1129), .B1(n_1131), .B2(n_1133), .Y(n_1128) );
INVx4_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx2_ASAP7_75t_L g998 ( .A(n_869), .Y(n_998) );
INVx1_ASAP7_75t_L g1014 ( .A(n_871), .Y(n_1014) );
INVx3_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx2_ASAP7_75t_L g1034 ( .A(n_873), .Y(n_1034) );
INVx2_ASAP7_75t_L g1334 ( .A(n_873), .Y(n_1334) );
INVx3_ASAP7_75t_L g980 ( .A(n_875), .Y(n_980) );
NAND4xp25_ASAP7_75t_L g876 ( .A(n_877), .B(n_879), .C(n_881), .D(n_883), .Y(n_876) );
BUFx3_ASAP7_75t_L g1327 ( .A(n_882), .Y(n_1327) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
XNOR2x1_ASAP7_75t_L g886 ( .A(n_887), .B(n_919), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
XNOR2x1_ASAP7_75t_L g888 ( .A(n_889), .B(n_890), .Y(n_888) );
NOR2x1_ASAP7_75t_L g890 ( .A(n_891), .B(n_901), .Y(n_890) );
NAND4xp25_ASAP7_75t_L g891 ( .A(n_892), .B(n_897), .C(n_899), .D(n_900), .Y(n_891) );
BUFx6f_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx2_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
NAND3xp33_ASAP7_75t_L g901 ( .A(n_902), .B(n_912), .C(n_915), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_904), .B(n_908), .Y(n_903) );
INVx4_ASAP7_75t_L g986 ( .A(n_905), .Y(n_986) );
INVx3_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g1271 ( .A(n_910), .Y(n_1271) );
BUFx3_ASAP7_75t_L g1101 ( .A(n_911), .Y(n_1101) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx2_ASAP7_75t_L g1103 ( .A(n_918), .Y(n_1103) );
HB1xp67_ASAP7_75t_L g1176 ( .A(n_918), .Y(n_1176) );
OAI22x1_ASAP7_75t_L g919 ( .A1(n_920), .A2(n_946), .B1(n_947), .B2(n_968), .Y(n_919) );
INVx2_ASAP7_75t_L g968 ( .A(n_920), .Y(n_968) );
NAND4xp75_ASAP7_75t_L g921 ( .A(n_922), .B(n_927), .C(n_930), .D(n_940), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_923), .B(n_925), .Y(n_922) );
BUFx2_ASAP7_75t_SL g1321 ( .A(n_924), .Y(n_1321) );
BUFx3_ASAP7_75t_L g1181 ( .A(n_926), .Y(n_1181) );
AND2x2_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .Y(n_927) );
NOR2xp33_ASAP7_75t_L g930 ( .A(n_931), .B(n_935), .Y(n_930) );
OAI21xp33_ASAP7_75t_L g931 ( .A1(n_932), .A2(n_933), .B(n_934), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_936), .A2(n_937), .B1(n_938), .B2(n_939), .Y(n_935) );
HB1xp67_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
INVx2_ASAP7_75t_L g1227 ( .A(n_942), .Y(n_1227) );
INVx2_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
NOR2x1_ASAP7_75t_L g948 ( .A(n_949), .B(n_960), .Y(n_948) );
NAND4xp25_ASAP7_75t_L g949 ( .A(n_950), .B(n_952), .C(n_954), .D(n_958), .Y(n_949) );
BUFx3_ASAP7_75t_L g1100 ( .A(n_951), .Y(n_1100) );
INVx2_ASAP7_75t_L g1171 ( .A(n_951), .Y(n_1171) );
BUFx2_ASAP7_75t_L g1330 ( .A(n_955), .Y(n_1330) );
NAND4xp25_ASAP7_75t_SL g960 ( .A(n_961), .B(n_965), .C(n_966), .D(n_967), .Y(n_960) );
BUFx6f_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
BUFx4f_ASAP7_75t_L g1157 ( .A(n_963), .Y(n_1157) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVxp67_ASAP7_75t_SL g1345 ( .A(n_972), .Y(n_1345) );
XOR2xp5_ASAP7_75t_L g972 ( .A(n_973), .B(n_1093), .Y(n_972) );
AO22x2_ASAP7_75t_L g973 ( .A1(n_974), .A2(n_1047), .B1(n_1090), .B2(n_1092), .Y(n_973) );
INVx1_ASAP7_75t_L g1092 ( .A(n_974), .Y(n_1092) );
AOI22xp5_ASAP7_75t_L g974 ( .A1(n_975), .A2(n_1019), .B1(n_1020), .B2(n_1046), .Y(n_974) );
INVx1_ASAP7_75t_L g1046 ( .A(n_975), .Y(n_1046) );
XNOR2xp5_ASAP7_75t_L g975 ( .A(n_976), .B(n_999), .Y(n_975) );
NAND4xp75_ASAP7_75t_L g977 ( .A(n_978), .B(n_989), .C(n_992), .D(n_995), .Y(n_977) );
NOR2xp67_ASAP7_75t_L g978 ( .A(n_979), .B(n_984), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_980), .A2(n_981), .B1(n_982), .B2(n_983), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g1169 ( .A1(n_982), .A2(n_1170), .B1(n_1171), .B2(n_1172), .Y(n_1169) );
OAI21xp5_ASAP7_75t_L g984 ( .A1(n_985), .A2(n_986), .B(n_987), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g1173 ( .A1(n_986), .A2(n_1174), .B1(n_1175), .B2(n_1176), .Y(n_1173) );
AND2x2_ASAP7_75t_L g989 ( .A(n_990), .B(n_991), .Y(n_989) );
AND2x2_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
NOR2xp33_ASAP7_75t_L g996 ( .A(n_997), .B(n_998), .Y(n_996) );
INVx1_ASAP7_75t_L g1086 ( .A(n_999), .Y(n_1086) );
HB1xp67_ASAP7_75t_L g1088 ( .A(n_999), .Y(n_1088) );
XOR2x2_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1018), .Y(n_999) );
NOR4xp75_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1006), .C(n_1009), .D(n_1012), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1004), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1008), .Y(n_1006) );
NAND2xp5_ASAP7_75t_SL g1009 ( .A(n_1010), .B(n_1011), .Y(n_1009) );
OAI21x1_ASAP7_75t_SL g1012 ( .A1(n_1013), .A2(n_1014), .B(n_1015), .Y(n_1012) );
INVx2_ASAP7_75t_SL g1019 ( .A(n_1020), .Y(n_1019) );
NAND4xp75_ASAP7_75t_SL g1021 ( .A(n_1022), .B(n_1026), .C(n_1030), .D(n_1035), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1025), .Y(n_1022) );
BUFx3_ASAP7_75t_L g1114 ( .A(n_1024), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1028), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1033), .Y(n_1030) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx2_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_1041), .A2(n_1042), .B1(n_1043), .B2(n_1044), .Y(n_1040) );
INVx2_ASAP7_75t_SL g1044 ( .A(n_1045), .Y(n_1044) );
OAI21xp5_ASAP7_75t_L g1047 ( .A1(n_1048), .A2(n_1085), .B(n_1087), .Y(n_1047) );
AOI22x1_ASAP7_75t_SL g1090 ( .A1(n_1048), .A2(n_1086), .B1(n_1088), .B2(n_1091), .Y(n_1090) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
INVx2_ASAP7_75t_L g1089 ( .A(n_1049), .Y(n_1089) );
AO22x2_ASAP7_75t_L g1049 ( .A1(n_1050), .A2(n_1051), .B1(n_1071), .B2(n_1084), .Y(n_1049) );
INVx2_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
INVx2_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
NAND4xp75_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1058), .C(n_1062), .D(n_1066), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1056), .Y(n_1054) );
BUFx2_ASAP7_75t_L g1165 ( .A(n_1057), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1060), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1064), .Y(n_1062) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1071), .Y(n_1084) );
NAND3x1_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1076), .C(n_1079), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1078), .Y(n_1076) );
AND4x1_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1081), .C(n_1082), .D(n_1083), .Y(n_1079) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1089), .Y(n_1087) );
INVx2_ASAP7_75t_L g1091 ( .A(n_1089), .Y(n_1091) );
AO22x2_ASAP7_75t_L g1093 ( .A1(n_1094), .A2(n_1095), .B1(n_1118), .B2(n_1190), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
BUFx2_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
XOR2x2_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1117), .Y(n_1096) );
NOR2x1_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1109), .Y(n_1097) );
NAND4xp25_ASAP7_75t_L g1098 ( .A(n_1099), .B(n_1102), .C(n_1104), .D(n_1107), .Y(n_1098) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1105), .Y(n_1188) );
INVx2_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
NAND4xp25_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1112), .C(n_1115), .D(n_1116), .Y(n_1109) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1118), .Y(n_1190) );
AO22x2_ASAP7_75t_L g1118 ( .A1(n_1119), .A2(n_1120), .B1(n_1160), .B2(n_1161), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
XOR2xp5_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1142), .Y(n_1120) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1122), .Y(n_1141) );
NOR2x1_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1135), .Y(n_1122) );
NAND3xp33_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1127), .C(n_1134), .Y(n_1123) );
CKINVDCx16_ASAP7_75t_R g1129 ( .A(n_1130), .Y(n_1129) );
CKINVDCx9p33_ASAP7_75t_R g1131 ( .A(n_1132), .Y(n_1131) );
NAND4xp25_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1137), .C(n_1138), .D(n_1139), .Y(n_1135) );
XNOR2xp5_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1144), .Y(n_1142) );
NOR2xp67_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1154), .Y(n_1144) );
NAND4xp25_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1147), .C(n_1149), .D(n_1150), .Y(n_1145) );
NOR2xp33_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1153), .Y(n_1151) );
INVx2_ASAP7_75t_L g1269 ( .A(n_1153), .Y(n_1269) );
NAND4xp25_ASAP7_75t_SL g1154 ( .A(n_1155), .B(n_1156), .C(n_1158), .D(n_1159), .Y(n_1154) );
INVx2_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
NAND4xp75_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1168), .C(n_1177), .D(n_1185), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1166), .Y(n_1163) );
NOR2x1_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1173), .Y(n_1168) );
OA21x2_ASAP7_75t_L g1223 ( .A1(n_1171), .A2(n_1224), .B(n_1225), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1182), .Y(n_1177) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
BUFx2_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
OAI21xp33_ASAP7_75t_L g1186 ( .A1(n_1187), .A2(n_1188), .B(n_1189), .Y(n_1186) );
INVxp67_ASAP7_75t_SL g1347 ( .A(n_1193), .Y(n_1347) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
OAI22xp33_ASAP7_75t_L g1194 ( .A1(n_1195), .A2(n_1275), .B1(n_1342), .B2(n_1343), .Y(n_1194) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1195), .Y(n_1342) );
XNOR2xp5_ASAP7_75t_L g1195 ( .A(n_1196), .B(n_1254), .Y(n_1195) );
AO22x2_ASAP7_75t_L g1196 ( .A1(n_1197), .A2(n_1236), .B1(n_1252), .B2(n_1253), .Y(n_1196) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1197), .Y(n_1253) );
XNOR2x1_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1217), .Y(n_1197) );
OAI22x1_ASAP7_75t_L g1198 ( .A1(n_1199), .A2(n_1206), .B1(n_1215), .B2(n_1216), .Y(n_1198) );
HB1xp67_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
NOR2xp33_ASAP7_75t_L g1215 ( .A(n_1200), .B(n_1207), .Y(n_1215) );
NAND4xp25_ASAP7_75t_L g1200 ( .A(n_1201), .B(n_1202), .C(n_1204), .D(n_1205), .Y(n_1200) );
NAND4xp25_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1209), .C(n_1211), .D(n_1214), .Y(n_1207) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1217), .Y(n_1274) );
NAND4xp75_ASAP7_75t_L g1218 ( .A(n_1219), .B(n_1223), .C(n_1230), .D(n_1233), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1220), .B(n_1221), .Y(n_1219) );
INVx2_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1232), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1234), .B(n_1235), .Y(n_1233) );
BUFx3_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1237), .Y(n_1252) );
XNOR2x1_ASAP7_75t_L g1294 ( .A(n_1237), .B(n_1295), .Y(n_1294) );
XNOR2x1_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1251), .Y(n_1237) );
NAND4xp75_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1242), .C(n_1245), .D(n_1248), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1241), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1244), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1246), .B(n_1247), .Y(n_1245) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
XNOR2xp5_ASAP7_75t_L g1255 ( .A(n_1256), .B(n_1274), .Y(n_1255) );
XNOR2x1_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1273), .Y(n_1256) );
OR2x2_ASAP7_75t_L g1257 ( .A(n_1258), .B(n_1263), .Y(n_1257) );
NAND4xp25_ASAP7_75t_SL g1258 ( .A(n_1259), .B(n_1260), .C(n_1261), .D(n_1262), .Y(n_1258) );
NAND3xp33_ASAP7_75t_L g1263 ( .A(n_1264), .B(n_1270), .C(n_1272), .Y(n_1263) );
INVxp67_ASAP7_75t_SL g1343 ( .A(n_1275), .Y(n_1343) );
AOI21xp5_ASAP7_75t_L g1275 ( .A1(n_1276), .A2(n_1313), .B(n_1341), .Y(n_1275) );
INVx2_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1277), .B(n_1314), .Y(n_1341) );
OA22x2_ASAP7_75t_L g1277 ( .A1(n_1278), .A2(n_1294), .B1(n_1311), .B2(n_1312), .Y(n_1277) );
INVx1_ASAP7_75t_SL g1311 ( .A(n_1278), .Y(n_1311) );
XOR2x2_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1293), .Y(n_1278) );
NOR2x1_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1286), .Y(n_1279) );
NAND4xp25_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1282), .C(n_1284), .D(n_1285), .Y(n_1280) );
HB1xp67_ASAP7_75t_L g1325 ( .A(n_1283), .Y(n_1325) );
NAND4xp25_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1289), .C(n_1290), .D(n_1291), .Y(n_1286) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1294), .Y(n_1312) );
XNOR2x1_ASAP7_75t_L g1295 ( .A(n_1296), .B(n_1297), .Y(n_1295) );
OR2x2_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1306), .Y(n_1297) );
NAND4xp25_ASAP7_75t_L g1298 ( .A(n_1299), .B(n_1301), .C(n_1302), .D(n_1303), .Y(n_1298) );
NAND4xp25_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1308), .C(n_1309), .D(n_1310), .Y(n_1306) );
INVx2_ASAP7_75t_SL g1313 ( .A(n_1314), .Y(n_1313) );
NAND4xp75_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1322), .C(n_1328), .D(n_1335), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1319), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1326), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1332), .Y(n_1328) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
endmodule