module fake_jpeg_25097_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVxp67_ASAP7_75t_SL g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_22),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_21),
.B(n_15),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_30),
.Y(n_35)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_27),
.C(n_22),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_23),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_29),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_24),
.A2(n_19),
.B1(n_14),
.B2(n_20),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_30),
.B1(n_24),
.B2(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_51),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_47),
.B(n_50),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

CKINVDCx10_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_24),
.B1(n_27),
.B2(n_23),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_27),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_57),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_41),
.Y(n_56)
);

FAx1_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_59),
.CI(n_16),
.CON(n_71),
.SN(n_71)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_36),
.Y(n_57)
);

AOI32xp33_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_34),
.A3(n_35),
.B1(n_13),
.B2(n_17),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_42),
.C(n_35),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_32),
.C(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_42),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_67),
.C(n_63),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_45),
.B(n_44),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_68),
.B(n_71),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_43),
.B1(n_48),
.B2(n_46),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_48),
.B1(n_20),
.B2(n_13),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_72),
.B(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_74),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_55),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_72),
.C(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_78),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_60),
.B(n_55),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_69),
.B(n_1),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_60),
.B1(n_16),
.B2(n_12),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_70),
.B1(n_74),
.B2(n_65),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_12),
.C(n_18),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_86),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_84),
.B(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_88),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_87),
.Y(n_94)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_93),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_0),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_95),
.B(n_7),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_79),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_97),
.B(n_1),
.Y(n_100)
);

AO21x2_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_80),
.B(n_3),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_97),
.A2(n_92),
.B(n_5),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_98),
.A2(n_100),
.B(n_4),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_8),
.B1(n_9),
.B2(n_4),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_102),
.C(n_9),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_4),
.Y(n_104)
);


endmodule