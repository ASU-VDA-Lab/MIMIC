module fake_netlist_1_3433_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_1), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_10), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_2), .B(n_7), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_14), .B(n_0), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_11), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_13), .B(n_0), .Y(n_18) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_17), .B(n_16), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_11), .B(n_15), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_19), .B(n_12), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_15), .Y(n_22) );
AOI22xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_20), .B1(n_12), .B2(n_11), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_21), .B(n_20), .Y(n_24) );
OAI22xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_22), .B1(n_1), .B2(n_2), .Y(n_25) );
AND2x2_ASAP7_75t_SL g26 ( .A(n_23), .B(n_0), .Y(n_26) );
O2A1O1Ixp33_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_1), .B(n_2), .C(n_3), .Y(n_27) );
AOI22xp33_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
NOR3xp33_ASAP7_75t_L g30 ( .A(n_28), .B(n_26), .C(n_5), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
OAI21xp5_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_9), .B(n_6), .Y(n_32) );
AOI22xp33_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_4), .B1(n_7), .B2(n_8), .Y(n_33) );
AOI22x1_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_31), .B1(n_8), .B2(n_9), .Y(n_34) );
endmodule