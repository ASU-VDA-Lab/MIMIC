module fake_netlist_1_1322_n_24 (n_3, n_1, n_2, n_0, n_24);
input n_3;
input n_1;
input n_2;
input n_0;
output n_24;
wire n_20;
wire n_5;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
wire n_6;
wire n_4;
wire n_7;
CKINVDCx5p33_ASAP7_75t_R g4 ( .A(n_2), .Y(n_4) );
CKINVDCx5p33_ASAP7_75t_R g5 ( .A(n_2), .Y(n_5) );
INVx2_ASAP7_75t_L g6 ( .A(n_1), .Y(n_6) );
CKINVDCx5p33_ASAP7_75t_R g7 ( .A(n_0), .Y(n_7) );
INVx4_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
OAI21x1_ASAP7_75t_L g9 ( .A1(n_6), .A2(n_0), .B(n_1), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_4), .B(n_0), .Y(n_10) );
AOI21xp5_ASAP7_75t_L g11 ( .A1(n_6), .A2(n_5), .B(n_3), .Y(n_11) );
AND2x4_ASAP7_75t_L g12 ( .A(n_8), .B(n_3), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_8), .B(n_10), .Y(n_13) );
BUFx2_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_13), .B(n_11), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_15), .B(n_12), .Y(n_18) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_17), .B(n_16), .Y(n_19) );
NOR3xp33_ASAP7_75t_L g20 ( .A(n_18), .B(n_12), .C(n_16), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_19), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_18), .Y(n_22) );
NOR2x1p5_ASAP7_75t_L g23 ( .A(n_21), .B(n_12), .Y(n_23) );
AOI22xp5_ASAP7_75t_SL g24 ( .A1(n_23), .A2(n_22), .B1(n_21), .B2(n_7), .Y(n_24) );
endmodule