module real_aes_7187_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_713, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_713;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g457 ( .A1(n_0), .A2(n_195), .B(n_458), .C(n_461), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_1), .B(n_452), .Y(n_462) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
INVx1_ASAP7_75t_L g230 ( .A(n_3), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_4), .B(n_147), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_5), .A2(n_447), .B(n_535), .Y(n_534) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_6), .A2(n_170), .B(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_7), .A2(n_36), .B1(n_140), .B2(n_164), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_8), .B(n_170), .Y(n_242) );
AND2x6_ASAP7_75t_L g155 ( .A(n_9), .B(n_156), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_10), .A2(n_155), .B(n_438), .C(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_11), .B(n_37), .Y(n_114) );
INVx1_ASAP7_75t_L g705 ( .A(n_11), .Y(n_705) );
INVx1_ASAP7_75t_L g136 ( .A(n_12), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_13), .B(n_145), .Y(n_178) );
INVx1_ASAP7_75t_L g222 ( .A(n_14), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_15), .B(n_147), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_16), .B(n_171), .Y(n_209) );
AO32x2_ASAP7_75t_L g192 ( .A1(n_17), .A2(n_169), .A3(n_170), .B1(n_193), .B2(n_197), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_18), .B(n_140), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_19), .B(n_171), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_20), .A2(n_52), .B1(n_140), .B2(n_164), .Y(n_196) );
AOI22xp33_ASAP7_75t_SL g167 ( .A1(n_21), .A2(n_79), .B1(n_140), .B2(n_145), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_22), .B(n_140), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_23), .A2(n_169), .B(n_438), .C(n_485), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_24), .A2(n_169), .B(n_438), .C(n_500), .Y(n_499) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_25), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_26), .B(n_132), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_27), .A2(n_117), .B1(n_118), .B2(n_119), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_27), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_28), .A2(n_447), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_29), .B(n_132), .Y(n_157) );
INVx2_ASAP7_75t_L g142 ( .A(n_30), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_31), .A2(n_444), .B(n_470), .C(n_471), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_32), .B(n_140), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_33), .B(n_132), .Y(n_185) );
OAI22xp5_ASAP7_75t_SL g697 ( .A1(n_34), .A2(n_41), .B1(n_428), .B2(n_698), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_34), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_35), .B(n_180), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_37), .B(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_38), .B(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_39), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_40), .B(n_147), .Y(n_523) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_41), .A2(n_123), .B1(n_428), .B2(n_429), .Y(n_122) );
INVx1_ASAP7_75t_L g428 ( .A(n_41), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_42), .B(n_447), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_43), .A2(n_444), .B(n_470), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_44), .B(n_140), .Y(n_237) );
INVx1_ASAP7_75t_L g459 ( .A(n_45), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g163 ( .A1(n_46), .A2(n_88), .B1(n_164), .B2(n_165), .Y(n_163) );
INVx1_ASAP7_75t_L g522 ( .A(n_47), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_48), .B(n_140), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_49), .B(n_140), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_50), .B(n_447), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_51), .B(n_228), .Y(n_241) );
AOI22xp33_ASAP7_75t_SL g213 ( .A1(n_53), .A2(n_57), .B1(n_140), .B2(n_145), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_54), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_55), .B(n_140), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_56), .B(n_140), .Y(n_250) );
INVx1_ASAP7_75t_L g156 ( .A(n_58), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_59), .B(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_60), .B(n_452), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_61), .A2(n_225), .B(n_228), .C(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_62), .B(n_140), .Y(n_231) );
INVx1_ASAP7_75t_L g135 ( .A(n_63), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_64), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_65), .B(n_147), .Y(n_475) );
AO32x2_ASAP7_75t_L g161 ( .A1(n_66), .A2(n_162), .A3(n_168), .B1(n_169), .B2(n_170), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_67), .B(n_148), .Y(n_512) );
INVx1_ASAP7_75t_L g249 ( .A(n_68), .Y(n_249) );
INVx1_ASAP7_75t_L g143 ( .A(n_69), .Y(n_143) );
CKINVDCx16_ASAP7_75t_R g455 ( .A(n_70), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_71), .B(n_474), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g437 ( .A1(n_72), .A2(n_438), .B(n_440), .C(n_444), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_73), .B(n_145), .Y(n_144) );
CKINVDCx16_ASAP7_75t_R g536 ( .A(n_74), .Y(n_536) );
INVx1_ASAP7_75t_L g710 ( .A(n_75), .Y(n_710) );
AOI22xp33_ASAP7_75t_SL g100 ( .A1(n_76), .A2(n_101), .B1(n_700), .B2(n_711), .Y(n_100) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_77), .B(n_473), .Y(n_487) );
AOI22xp5_ASAP7_75t_SL g115 ( .A1(n_78), .A2(n_111), .B1(n_116), .B2(n_690), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_80), .B(n_164), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_81), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_82), .B(n_145), .Y(n_152) );
INVx2_ASAP7_75t_L g133 ( .A(n_83), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_84), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_85), .B(n_166), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_86), .B(n_145), .Y(n_238) );
OR2x2_ASAP7_75t_L g110 ( .A(n_87), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g121 ( .A(n_87), .Y(n_121) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_89), .A2(n_99), .B1(n_145), .B2(n_146), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_90), .B(n_447), .Y(n_468) );
INVx1_ASAP7_75t_L g472 ( .A(n_91), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_92), .Y(n_107) );
INVxp67_ASAP7_75t_L g539 ( .A(n_93), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_94), .B(n_145), .Y(n_247) );
INVx1_ASAP7_75t_L g441 ( .A(n_95), .Y(n_441) );
INVx1_ASAP7_75t_L g508 ( .A(n_96), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_97), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g524 ( .A(n_98), .B(n_132), .Y(n_524) );
AOI22x1_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_105), .B1(n_115), .B2(n_693), .Y(n_101) );
NOR2xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_106), .A2(n_694), .B(n_699), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_110), .Y(n_699) );
NOR2x2_ASAP7_75t_L g692 ( .A(n_111), .B(n_121), .Y(n_692) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
NAND3xp33_ASAP7_75t_SL g707 ( .A(n_113), .B(n_121), .C(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AO22x2_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_122), .B1(n_430), .B2(n_689), .Y(n_120) );
INVx1_ASAP7_75t_L g689 ( .A(n_121), .Y(n_689) );
INVx1_ASAP7_75t_L g429 ( .A(n_123), .Y(n_429) );
OAI22xp5_ASAP7_75t_SL g695 ( .A1(n_123), .A2(n_429), .B1(n_696), .B2(n_697), .Y(n_695) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_349), .Y(n_123) );
NAND3xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_298), .C(n_340), .Y(n_124) );
AOI211xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_203), .B(n_252), .C(n_274), .Y(n_125) );
OAI211xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_158), .B(n_186), .C(n_198), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_128), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g361 ( .A(n_128), .B(n_278), .Y(n_361) );
BUFx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g263 ( .A(n_129), .B(n_189), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_129), .B(n_174), .Y(n_380) );
INVx1_ASAP7_75t_L g398 ( .A(n_129), .Y(n_398) );
AND2x2_ASAP7_75t_L g407 ( .A(n_129), .B(n_295), .Y(n_407) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OR2x2_ASAP7_75t_L g290 ( .A(n_130), .B(n_174), .Y(n_290) );
AND2x2_ASAP7_75t_L g348 ( .A(n_130), .B(n_295), .Y(n_348) );
INVx1_ASAP7_75t_L g392 ( .A(n_130), .Y(n_392) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OR2x2_ASAP7_75t_L g269 ( .A(n_131), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g277 ( .A(n_131), .Y(n_277) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_131), .Y(n_317) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_137), .B(n_157), .Y(n_131) );
INVx2_ASAP7_75t_L g168 ( .A(n_132), .Y(n_168) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_132), .A2(n_175), .B(n_185), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_132), .A2(n_468), .B(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g491 ( .A(n_132), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_132), .A2(n_519), .B(n_520), .Y(n_518) );
AND2x2_ASAP7_75t_SL g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_L g171 ( .A(n_133), .B(n_134), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
OAI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_150), .B(n_155), .Y(n_137) );
O2A1O1Ixp5_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_143), .B(n_144), .C(n_147), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_140), .Y(n_443) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g164 ( .A(n_141), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_141), .Y(n_165) );
AND2x6_ASAP7_75t_L g438 ( .A(n_141), .B(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g146 ( .A(n_142), .Y(n_146) );
INVx1_ASAP7_75t_L g229 ( .A(n_142), .Y(n_229) );
INVx2_ASAP7_75t_L g223 ( .A(n_145), .Y(n_223) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g195 ( .A(n_147), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_147), .A2(n_237), .B(n_238), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_147), .A2(n_246), .B(n_247), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_147), .B(n_539), .Y(n_538) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
OAI22xp5_ASAP7_75t_SL g162 ( .A1(n_148), .A2(n_163), .B1(n_166), .B2(n_167), .Y(n_162) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_149), .Y(n_154) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_149), .Y(n_166) );
INVx1_ASAP7_75t_L g180 ( .A(n_149), .Y(n_180) );
INVx1_ASAP7_75t_L g439 ( .A(n_149), .Y(n_439) );
AND2x2_ASAP7_75t_L g448 ( .A(n_149), .B(n_229), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_153), .Y(n_150) );
INVx1_ASAP7_75t_L g225 ( .A(n_153), .Y(n_225) );
INVx4_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g474 ( .A(n_154), .Y(n_474) );
BUFx3_ASAP7_75t_L g169 ( .A(n_155), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g175 ( .A1(n_155), .A2(n_176), .B(n_181), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_155), .A2(n_221), .B(n_226), .Y(n_220) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_155), .A2(n_236), .B(n_239), .Y(n_235) );
INVx4_ASAP7_75t_SL g445 ( .A(n_155), .Y(n_445) );
AND2x4_ASAP7_75t_L g447 ( .A(n_155), .B(n_448), .Y(n_447) );
NAND2x1p5_ASAP7_75t_L g509 ( .A(n_155), .B(n_448), .Y(n_509) );
INVxp67_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_172), .Y(n_159) );
AND2x2_ASAP7_75t_L g256 ( .A(n_160), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g289 ( .A(n_160), .Y(n_289) );
OR2x2_ASAP7_75t_L g415 ( .A(n_160), .B(n_416), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_160), .B(n_174), .Y(n_419) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g189 ( .A(n_161), .Y(n_189) );
INVx1_ASAP7_75t_L g201 ( .A(n_161), .Y(n_201) );
AND2x2_ASAP7_75t_L g278 ( .A(n_161), .B(n_191), .Y(n_278) );
AND2x2_ASAP7_75t_L g318 ( .A(n_161), .B(n_192), .Y(n_318) );
INVx2_ASAP7_75t_L g461 ( .A(n_165), .Y(n_461) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_165), .Y(n_476) );
INVx2_ASAP7_75t_L g184 ( .A(n_166), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_166), .A2(n_194), .B1(n_195), .B2(n_196), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_166), .A2(n_195), .B1(n_212), .B2(n_213), .Y(n_211) );
INVx4_ASAP7_75t_L g460 ( .A(n_166), .Y(n_460) );
INVx1_ASAP7_75t_L g488 ( .A(n_168), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g210 ( .A(n_169), .B(n_211), .C(n_214), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g244 ( .A1(n_169), .A2(n_245), .B(n_248), .Y(n_244) );
INVx4_ASAP7_75t_L g214 ( .A(n_170), .Y(n_214) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_170), .A2(n_235), .B(n_242), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_170), .A2(n_498), .B(n_499), .Y(n_497) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_170), .Y(n_533) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g197 ( .A(n_171), .Y(n_197) );
INVxp67_ASAP7_75t_L g360 ( .A(n_172), .Y(n_360) );
AND2x4_ASAP7_75t_L g385 ( .A(n_172), .B(n_278), .Y(n_385) );
BUFx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_SL g276 ( .A(n_173), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g190 ( .A(n_174), .B(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g264 ( .A(n_174), .B(n_192), .Y(n_264) );
INVx1_ASAP7_75t_L g270 ( .A(n_174), .Y(n_270) );
INVx2_ASAP7_75t_L g296 ( .A(n_174), .Y(n_296) );
AND2x2_ASAP7_75t_L g312 ( .A(n_174), .B(n_313), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_179), .Y(n_176) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_184), .Y(n_181) );
O2A1O1Ixp5_ASAP7_75t_L g248 ( .A1(n_184), .A2(n_227), .B(n_249), .C(n_250), .Y(n_248) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_187), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_190), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
BUFx2_ASAP7_75t_L g267 ( .A(n_189), .Y(n_267) );
AND2x2_ASAP7_75t_L g375 ( .A(n_189), .B(n_191), .Y(n_375) );
AND2x2_ASAP7_75t_L g292 ( .A(n_190), .B(n_277), .Y(n_292) );
AND2x2_ASAP7_75t_L g391 ( .A(n_190), .B(n_392), .Y(n_391) );
NOR2xp67_ASAP7_75t_L g313 ( .A(n_191), .B(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g416 ( .A(n_191), .B(n_277), .Y(n_416) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
BUFx2_ASAP7_75t_L g202 ( .A(n_192), .Y(n_202) );
AND2x2_ASAP7_75t_L g295 ( .A(n_192), .B(n_296), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_195), .A2(n_227), .B(n_230), .C(n_231), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_195), .A2(n_240), .B(n_241), .Y(n_239) );
INVx2_ASAP7_75t_L g219 ( .A(n_197), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_197), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_202), .Y(n_199) );
AND2x2_ASAP7_75t_L g341 ( .A(n_200), .B(n_276), .Y(n_341) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_201), .B(n_277), .Y(n_326) );
INVx2_ASAP7_75t_L g325 ( .A(n_202), .Y(n_325) );
OAI222xp33_ASAP7_75t_L g329 ( .A1(n_202), .A2(n_269), .B1(n_330), .B2(n_332), .C1(n_333), .C2(n_336), .Y(n_329) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_215), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g254 ( .A(n_207), .Y(n_254) );
OR2x2_ASAP7_75t_L g365 ( .A(n_207), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx3_ASAP7_75t_L g287 ( .A(n_208), .Y(n_287) );
NOR2x1_ASAP7_75t_L g338 ( .A(n_208), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g344 ( .A(n_208), .B(n_258), .Y(n_344) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
INVx1_ASAP7_75t_L g305 ( .A(n_209), .Y(n_305) );
AO21x1_ASAP7_75t_L g304 ( .A1(n_211), .A2(n_214), .B(n_305), .Y(n_304) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_214), .A2(n_436), .B(n_449), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_214), .B(n_450), .Y(n_449) );
INVx3_ASAP7_75t_L g452 ( .A(n_214), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_214), .B(n_478), .Y(n_477) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_214), .A2(n_507), .B(n_514), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_215), .A2(n_308), .B1(n_347), .B2(n_348), .Y(n_346) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_233), .Y(n_215) );
INVx3_ASAP7_75t_L g280 ( .A(n_216), .Y(n_280) );
OR2x2_ASAP7_75t_L g413 ( .A(n_216), .B(n_289), .Y(n_413) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g286 ( .A(n_217), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g302 ( .A(n_217), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g310 ( .A(n_217), .B(n_258), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_217), .B(n_234), .Y(n_366) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g257 ( .A(n_218), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g261 ( .A(n_218), .B(n_234), .Y(n_261) );
AND2x2_ASAP7_75t_L g337 ( .A(n_218), .B(n_284), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_218), .B(n_243), .Y(n_377) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_232), .Y(n_218) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_219), .A2(n_244), .B(n_251), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_224), .C(n_225), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_223), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_223), .A2(n_512), .B(n_513), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_L g440 ( .A1(n_225), .A2(n_441), .B(n_442), .C(n_443), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_227), .A2(n_486), .B(n_487), .Y(n_485) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_233), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g293 ( .A(n_233), .B(n_254), .Y(n_293) );
AND2x2_ASAP7_75t_L g297 ( .A(n_233), .B(n_287), .Y(n_297) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_243), .Y(n_233) );
INVx3_ASAP7_75t_L g258 ( .A(n_234), .Y(n_258) );
AND2x2_ASAP7_75t_L g283 ( .A(n_234), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g418 ( .A(n_234), .B(n_401), .Y(n_418) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_243), .Y(n_272) );
INVx2_ASAP7_75t_L g284 ( .A(n_243), .Y(n_284) );
AND2x2_ASAP7_75t_L g328 ( .A(n_243), .B(n_304), .Y(n_328) );
INVx1_ASAP7_75t_L g371 ( .A(n_243), .Y(n_371) );
OR2x2_ASAP7_75t_L g402 ( .A(n_243), .B(n_304), .Y(n_402) );
AND2x2_ASAP7_75t_L g422 ( .A(n_243), .B(n_258), .Y(n_422) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_255), .B(n_259), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g260 ( .A(n_254), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_254), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g379 ( .A(n_256), .Y(n_379) );
INVx2_ASAP7_75t_SL g273 ( .A(n_257), .Y(n_273) );
AND2x2_ASAP7_75t_L g393 ( .A(n_257), .B(n_287), .Y(n_393) );
INVx2_ASAP7_75t_L g339 ( .A(n_258), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_258), .B(n_371), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_262), .B1(n_265), .B2(n_271), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_261), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_SL g427 ( .A(n_261), .Y(n_427) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g352 ( .A(n_263), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_263), .B(n_295), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_264), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g368 ( .A(n_264), .B(n_317), .Y(n_368) );
INVx2_ASAP7_75t_L g424 ( .A(n_264), .Y(n_424) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
AND2x2_ASAP7_75t_L g294 ( .A(n_267), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_267), .B(n_312), .Y(n_345) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_269), .B(n_289), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g406 ( .A(n_272), .Y(n_406) );
O2A1O1Ixp33_ASAP7_75t_SL g356 ( .A1(n_273), .A2(n_357), .B(n_359), .C(n_362), .Y(n_356) );
OR2x2_ASAP7_75t_L g383 ( .A(n_273), .B(n_287), .Y(n_383) );
OAI221xp5_ASAP7_75t_SL g274 ( .A1(n_275), .A2(n_279), .B1(n_281), .B2(n_288), .C(n_291), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_276), .B(n_278), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_276), .B(n_325), .Y(n_332) );
AND2x2_ASAP7_75t_L g374 ( .A(n_276), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g410 ( .A(n_276), .Y(n_410) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_277), .Y(n_301) );
INVx1_ASAP7_75t_L g314 ( .A(n_277), .Y(n_314) );
NOR2xp67_ASAP7_75t_L g334 ( .A(n_280), .B(n_335), .Y(n_334) );
INVxp67_ASAP7_75t_L g388 ( .A(n_280), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_280), .B(n_328), .Y(n_404) );
INVx2_ASAP7_75t_L g390 ( .A(n_281), .Y(n_390) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_285), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g331 ( .A(n_283), .B(n_302), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_L g340 ( .A1(n_283), .A2(n_299), .B(n_341), .C(n_342), .Y(n_340) );
AND2x2_ASAP7_75t_L g309 ( .A(n_284), .B(n_304), .Y(n_309) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_288), .B(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
OR2x2_ASAP7_75t_L g357 ( .A(n_289), .B(n_358), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_293), .B1(n_294), .B2(n_297), .Y(n_291) );
INVx1_ASAP7_75t_L g411 ( .A(n_293), .Y(n_411) );
INVx1_ASAP7_75t_L g358 ( .A(n_295), .Y(n_358) );
INVx1_ASAP7_75t_L g409 ( .A(n_297), .Y(n_409) );
AOI211xp5_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_302), .B(n_306), .C(n_329), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g321 ( .A(n_301), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g372 ( .A(n_302), .Y(n_372) );
AND2x2_ASAP7_75t_L g421 ( .A(n_302), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OAI21xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_311), .B(n_319), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx2_ASAP7_75t_L g335 ( .A(n_309), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_309), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g327 ( .A(n_310), .B(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g403 ( .A(n_310), .Y(n_403) );
OAI32xp33_ASAP7_75t_L g414 ( .A1(n_310), .A2(n_362), .A3(n_369), .B1(n_410), .B2(n_415), .Y(n_414) );
NOR2xp33_ASAP7_75t_SL g311 ( .A(n_312), .B(n_315), .Y(n_311) );
INVx1_ASAP7_75t_SL g382 ( .A(n_312), .Y(n_382) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_SL g322 ( .A(n_318), .Y(n_322) );
OAI21xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_323), .B(n_327), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_321), .A2(n_369), .B1(n_395), .B2(n_397), .Y(n_394) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_325), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g362 ( .A(n_328), .Y(n_362) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2x1p5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g355 ( .A(n_339), .Y(n_355) );
OAI21xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_345), .B(n_346), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_348), .A2(n_390), .B1(n_391), .B2(n_393), .C(n_394), .Y(n_389) );
NAND5xp2_ASAP7_75t_L g349 ( .A(n_350), .B(n_373), .C(n_389), .D(n_399), .E(n_417), .Y(n_349) );
AOI211xp5_ASAP7_75t_SL g350 ( .A1(n_351), .A2(n_353), .B(n_356), .C(n_363), .Y(n_350) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g420 ( .A(n_357), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
OAI22xp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B1(n_367), .B2(n_369), .Y(n_363) );
INVx1_ASAP7_75t_SL g396 ( .A(n_366), .Y(n_396) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI322xp33_ASAP7_75t_L g378 ( .A1(n_369), .A2(n_379), .A3(n_380), .B1(n_381), .B2(n_382), .C1(n_383), .C2(n_384), .Y(n_378) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
INVx1_ASAP7_75t_L g381 ( .A(n_371), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_371), .B(n_396), .Y(n_395) );
AOI211xp5_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_376), .B(n_378), .C(n_386), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI22xp33_ASAP7_75t_L g408 ( .A1(n_382), .A2(n_409), .B1(n_410), .B2(n_411), .Y(n_408) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g425 ( .A(n_392), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_407), .B1(n_408), .B2(n_412), .C(n_414), .Y(n_399) );
OAI211xp5_ASAP7_75t_SL g400 ( .A1(n_401), .A2(n_403), .B(n_404), .C(n_405), .Y(n_400) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g426 ( .A(n_402), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_420), .B2(n_421), .C(n_423), .Y(n_417) );
AOI21xp33_ASAP7_75t_SL g423 ( .A1(n_424), .A2(n_425), .B(n_426), .Y(n_423) );
NAND2x1p5_ASAP7_75t_L g430 ( .A(n_431), .B(n_632), .Y(n_430) );
AND4x1_ASAP7_75t_L g431 ( .A(n_432), .B(n_572), .C(n_587), .D(n_612), .Y(n_431) );
NOR2xp33_ASAP7_75t_SL g432 ( .A(n_433), .B(n_545), .Y(n_432) );
OAI21xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_463), .B(n_525), .Y(n_433) );
AND2x2_ASAP7_75t_L g575 ( .A(n_434), .B(n_480), .Y(n_575) );
AND2x2_ASAP7_75t_L g588 ( .A(n_434), .B(n_479), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_434), .B(n_464), .Y(n_638) );
INVx1_ASAP7_75t_L g642 ( .A(n_434), .Y(n_642) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_451), .Y(n_434) );
INVx2_ASAP7_75t_L g559 ( .A(n_435), .Y(n_559) );
BUFx2_ASAP7_75t_L g586 ( .A(n_435), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_446), .Y(n_436) );
INVx5_ASAP7_75t_L g456 ( .A(n_438), .Y(n_456) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
O2A1O1Ixp33_ASAP7_75t_SL g454 ( .A1(n_445), .A2(n_455), .B(n_456), .C(n_457), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_445), .A2(n_456), .B(n_536), .C(n_537), .Y(n_535) );
BUFx2_ASAP7_75t_L g483 ( .A(n_447), .Y(n_483) );
AND2x2_ASAP7_75t_L g526 ( .A(n_451), .B(n_480), .Y(n_526) );
INVx2_ASAP7_75t_L g542 ( .A(n_451), .Y(n_542) );
AND2x2_ASAP7_75t_L g551 ( .A(n_451), .B(n_479), .Y(n_551) );
AND2x2_ASAP7_75t_L g630 ( .A(n_451), .B(n_559), .Y(n_630) );
OA21x2_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B(n_462), .Y(n_451) );
INVx2_ASAP7_75t_L g470 ( .A(n_456), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_492), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_464), .B(n_557), .Y(n_595) );
INVx1_ASAP7_75t_L g683 ( .A(n_464), .Y(n_683) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_479), .Y(n_464) );
AND2x2_ASAP7_75t_L g541 ( .A(n_465), .B(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g555 ( .A(n_465), .B(n_556), .Y(n_555) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_465), .Y(n_584) );
OR2x2_ASAP7_75t_L g616 ( .A(n_465), .B(n_558), .Y(n_616) );
AND2x2_ASAP7_75t_L g624 ( .A(n_465), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g657 ( .A(n_465), .B(n_626), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_465), .B(n_526), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_465), .B(n_586), .Y(n_682) );
AND2x2_ASAP7_75t_L g688 ( .A(n_465), .B(n_575), .Y(n_688) );
INVx5_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g548 ( .A(n_466), .Y(n_548) );
AND2x2_ASAP7_75t_L g578 ( .A(n_466), .B(n_558), .Y(n_578) );
AND2x2_ASAP7_75t_L g611 ( .A(n_466), .B(n_571), .Y(n_611) );
AND2x2_ASAP7_75t_L g631 ( .A(n_466), .B(n_480), .Y(n_631) );
AND2x2_ASAP7_75t_L g665 ( .A(n_466), .B(n_531), .Y(n_665) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_477), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B(n_475), .C(n_476), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_473), .A2(n_476), .B(n_522), .C(n_523), .Y(n_521) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x4_ASAP7_75t_L g571 ( .A(n_479), .B(n_542), .Y(n_571) );
AND2x2_ASAP7_75t_L g582 ( .A(n_479), .B(n_578), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_479), .B(n_558), .Y(n_621) );
INVx2_ASAP7_75t_L g636 ( .A(n_479), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_479), .B(n_570), .Y(n_659) );
AND2x2_ASAP7_75t_L g678 ( .A(n_479), .B(n_630), .Y(n_678) );
INVx5_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_480), .Y(n_577) );
AND2x2_ASAP7_75t_L g585 ( .A(n_480), .B(n_586), .Y(n_585) );
AND2x4_ASAP7_75t_L g626 ( .A(n_480), .B(n_542), .Y(n_626) );
OR2x6_ASAP7_75t_L g480 ( .A(n_481), .B(n_489), .Y(n_480) );
AOI21xp5_ASAP7_75t_SL g481 ( .A1(n_482), .A2(n_484), .B(n_488), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .Y(n_493) );
AND2x2_ASAP7_75t_L g549 ( .A(n_494), .B(n_532), .Y(n_549) );
INVx1_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_495), .B(n_506), .Y(n_529) );
OR2x2_ASAP7_75t_L g562 ( .A(n_495), .B(n_532), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_495), .B(n_532), .Y(n_567) );
AND2x2_ASAP7_75t_L g594 ( .A(n_495), .B(n_531), .Y(n_594) );
AND2x2_ASAP7_75t_L g646 ( .A(n_495), .B(n_505), .Y(n_646) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_496), .B(n_516), .Y(n_554) );
AND2x2_ASAP7_75t_L g590 ( .A(n_496), .B(n_506), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_503), .B(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g580 ( .A(n_504), .B(n_562), .Y(n_580) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_516), .Y(n_504) );
OAI322xp33_ASAP7_75t_L g545 ( .A1(n_505), .A2(n_546), .A3(n_550), .B1(n_552), .B2(n_555), .C1(n_560), .C2(n_568), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_505), .B(n_531), .Y(n_553) );
OR2x2_ASAP7_75t_L g563 ( .A(n_505), .B(n_517), .Y(n_563) );
AND2x2_ASAP7_75t_L g565 ( .A(n_505), .B(n_517), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_505), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_505), .B(n_532), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_505), .B(n_661), .Y(n_660) );
INVx5_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_506), .B(n_549), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B(n_510), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_516), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g543 ( .A(n_516), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_516), .B(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g605 ( .A(n_516), .B(n_532), .Y(n_605) );
AOI211xp5_ASAP7_75t_SL g633 ( .A1(n_516), .A2(n_634), .B(n_637), .C(n_649), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_516), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g671 ( .A(n_516), .B(n_646), .Y(n_671) );
INVx5_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g599 ( .A(n_517), .B(n_532), .Y(n_599) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_517), .Y(n_608) );
AND2x2_ASAP7_75t_L g648 ( .A(n_517), .B(n_646), .Y(n_648) );
AND2x2_ASAP7_75t_SL g679 ( .A(n_517), .B(n_549), .Y(n_679) );
AND2x2_ASAP7_75t_L g686 ( .A(n_517), .B(n_645), .Y(n_686) );
OR2x6_ASAP7_75t_L g517 ( .A(n_518), .B(n_524), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B1(n_541), .B2(n_543), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_526), .B(n_548), .Y(n_596) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g544 ( .A(n_529), .Y(n_544) );
OR2x2_ASAP7_75t_L g604 ( .A(n_529), .B(n_605), .Y(n_604) );
OAI221xp5_ASAP7_75t_SL g652 ( .A1(n_529), .A2(n_653), .B1(n_655), .B2(n_656), .C(n_658), .Y(n_652) );
INVx2_ASAP7_75t_L g591 ( .A(n_530), .Y(n_591) );
AND2x2_ASAP7_75t_L g564 ( .A(n_531), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g654 ( .A(n_531), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_531), .B(n_646), .Y(n_667) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVxp67_ASAP7_75t_L g609 ( .A(n_532), .Y(n_609) );
AND2x2_ASAP7_75t_L g645 ( .A(n_532), .B(n_646), .Y(n_645) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B(n_540), .Y(n_532) );
AND2x2_ASAP7_75t_L g647 ( .A(n_541), .B(n_586), .Y(n_647) );
AND2x2_ASAP7_75t_L g557 ( .A(n_542), .B(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_542), .B(n_615), .Y(n_614) );
NOR2xp33_ASAP7_75t_SL g628 ( .A(n_544), .B(n_591), .Y(n_628) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g634 ( .A(n_547), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
OR2x2_ASAP7_75t_L g620 ( .A(n_548), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g685 ( .A(n_548), .B(n_630), .Y(n_685) );
INVx2_ASAP7_75t_L g618 ( .A(n_549), .Y(n_618) );
NAND4xp25_ASAP7_75t_SL g681 ( .A(n_550), .B(n_682), .C(n_683), .D(n_684), .Y(n_681) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_551), .B(n_615), .Y(n_650) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_SL g687 ( .A(n_554), .Y(n_687) );
O2A1O1Ixp33_ASAP7_75t_SL g649 ( .A1(n_555), .A2(n_618), .B(n_622), .C(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g644 ( .A(n_557), .B(n_636), .Y(n_644) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_558), .Y(n_570) );
INVx1_ASAP7_75t_L g625 ( .A(n_558), .Y(n_625) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_559), .Y(n_602) );
AOI211xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_563), .B(n_564), .C(n_566), .Y(n_560) );
AND2x2_ASAP7_75t_L g581 ( .A(n_561), .B(n_565), .Y(n_581) );
OAI322xp33_ASAP7_75t_SL g619 ( .A1(n_561), .A2(n_620), .A3(n_622), .B1(n_623), .B2(n_627), .C1(n_628), .C2(n_629), .Y(n_619) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g641 ( .A(n_563), .B(n_567), .Y(n_641) );
INVx1_ASAP7_75t_L g622 ( .A(n_565), .Y(n_622) );
INVx1_ASAP7_75t_SL g640 ( .A(n_567), .Y(n_640) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
AOI222xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_579), .B1(n_581), .B2(n_582), .C1(n_583), .C2(n_713), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_574), .B(n_576), .Y(n_573) );
OAI322xp33_ASAP7_75t_L g662 ( .A1(n_574), .A2(n_636), .A3(n_641), .B1(n_663), .B2(n_664), .C1(n_666), .C2(n_667), .Y(n_662) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_575), .A2(n_589), .B1(n_613), .B2(n_617), .C(n_619), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
OAI222xp33_ASAP7_75t_L g592 ( .A1(n_580), .A2(n_593), .B1(n_595), .B2(n_596), .C1(n_597), .C2(n_600), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_582), .A2(n_589), .B1(n_659), .B2(n_660), .Y(n_658) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
AOI211xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B(n_592), .C(n_603), .Y(n_587) );
O2A1O1Ixp33_ASAP7_75t_L g668 ( .A1(n_589), .A2(n_626), .B(n_669), .C(n_672), .Y(n_668) );
AND2x4_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AND2x2_ASAP7_75t_L g598 ( .A(n_590), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_SL g661 ( .A(n_594), .Y(n_661) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_601), .B(n_626), .Y(n_655) );
BUFx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI21xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_606), .B(n_610), .Y(n_603) );
OAI221xp5_ASAP7_75t_SL g672 ( .A1(n_604), .A2(n_673), .B1(n_674), .B2(n_675), .C(n_676), .Y(n_672) );
INVxp33_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_608), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_615), .B(n_626), .Y(n_666) );
INVx2_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
AND2x2_ASAP7_75t_L g677 ( .A(n_630), .B(n_636), .Y(n_677) );
AND4x1_ASAP7_75t_L g632 ( .A(n_633), .B(n_651), .C(n_668), .D(n_680), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI221xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_639), .B1(n_641), .B2(n_642), .C(n_643), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B1(n_647), .B2(n_648), .Y(n_643) );
INVx1_ASAP7_75t_L g673 ( .A(n_644), .Y(n_673) );
INVx1_ASAP7_75t_SL g663 ( .A(n_648), .Y(n_663) );
NOR2xp33_ASAP7_75t_SL g651 ( .A(n_652), .B(n_662), .Y(n_651) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_664), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_671), .A2(n_677), .B1(n_678), .B2(n_679), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_686), .B1(n_687), .B2(n_688), .Y(n_680) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx3_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
CKINVDCx16_ASAP7_75t_R g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g711 ( .A(n_702), .Y(n_711) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_706), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
CKINVDCx14_ASAP7_75t_R g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
endmodule