module fake_jpeg_4006_n_143 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx16f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx11_ASAP7_75t_SL g13 ( 
.A(n_4),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx8_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_22),
.B(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx12_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_21),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_29),
.B1(n_14),
.B2(n_20),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_45),
.B1(n_49),
.B2(n_51),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_14),
.B1(n_20),
.B2(n_29),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_14),
.B1(n_20),
.B2(n_27),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_48),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_32),
.B(n_19),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_30),
.A2(n_26),
.B1(n_25),
.B2(n_27),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_31),
.Y(n_57)
);

AOI22x1_ASAP7_75t_L g51 ( 
.A1(n_31),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_50),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_27),
.B1(n_26),
.B2(n_39),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_52),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_58),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_36),
.B1(n_18),
.B2(n_17),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_24),
.C(n_23),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_51),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_63),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_50),
.B(n_51),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_65),
.B1(n_69),
.B2(n_74),
.Y(n_79)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_51),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_67),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_70),
.B(n_71),
.Y(n_78)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_73),
.B(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_43),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_64),
.C(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_72),
.B(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_80),
.Y(n_98)
);

AOI221xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_73),
.B1(n_72),
.B2(n_58),
.C(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_84),
.Y(n_89)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_59),
.B1(n_56),
.B2(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_75),
.C(n_61),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_95),
.C(n_86),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_92),
.B1(n_96),
.B2(n_91),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_66),
.B1(n_45),
.B2(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_46),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_15),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_41),
.A3(n_33),
.B1(n_49),
.B2(n_19),
.C1(n_23),
.C2(n_21),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_84),
.Y(n_106)
);

AND2x4_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_24),
.Y(n_95)
);

AO32x1_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_15),
.A3(n_36),
.B1(n_28),
.B2(n_21),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_96),
.B(n_42),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_102),
.B1(n_104),
.B2(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_105),
.C(n_10),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_109),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_23),
.C(n_62),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_108),
.C(n_97),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_62),
.C(n_42),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_101),
.A2(n_97),
.B(n_95),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_115),
.B(n_102),
.C(n_15),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_113),
.C(n_116),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_62),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_12),
.B1(n_10),
.B2(n_17),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_107),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_110),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_124),
.B(n_119),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_112),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_123),
.C(n_125),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_28),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_121),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_12),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_126),
.A2(n_127),
.B(n_129),
.Y(n_132)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_16),
.A3(n_12),
.B1(n_18),
.B2(n_17),
.C1(n_4),
.C2(n_6),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_6),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_120),
.A2(n_16),
.B(n_18),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_6),
.B(n_9),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_133),
.B(n_134),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_132),
.Y(n_139)
);

OAI21x1_ASAP7_75t_SL g136 ( 
.A1(n_131),
.A2(n_3),
.B(n_7),
.Y(n_136)
);

AOI31xp33_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_3),
.A3(n_7),
.B(n_8),
.Y(n_137)
);

OAI321xp33_ASAP7_75t_L g140 ( 
.A1(n_137),
.A2(n_139),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_1),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_140),
.A2(n_141),
.B1(n_0),
.B2(n_15),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_8),
.C(n_9),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_0),
.Y(n_143)
);


endmodule