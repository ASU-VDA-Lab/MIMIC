module fake_netlist_5_122_n_1784 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_408, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_397, n_111, n_155, n_43, n_116, n_22, n_423, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_417, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_325, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_422, n_72, n_104, n_41, n_415, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_430, n_313, n_88, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_239, n_420, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_441, n_312, n_429, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_425, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_437, n_66, n_177, n_60, n_403, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_409, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_391, n_434, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_52, n_278, n_110, n_1784);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_408;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_397;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_417;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_422;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_239;
input n_420;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_441;
input n_312;
input n_429;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_425;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_409;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_391;
input n_434;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1784;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_920;
wire n_1289;
wire n_1517;
wire n_1669;
wire n_976;
wire n_1449;
wire n_1566;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1556;
wire n_1384;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_464;
wire n_1582;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_647;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_1038;
wire n_520;
wire n_1369;
wire n_1660;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_1194;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_677;
wire n_1333;
wire n_1121;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1163;
wire n_906;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1591;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1562;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_450;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_824;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_815;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_1519;
wire n_950;
wire n_1553;
wire n_1346;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1305;
wire n_873;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_507;
wire n_1560;
wire n_1605;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_1307;
wire n_988;
wire n_814;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1149;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_1638;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1411;
wire n_622;
wire n_1577;
wire n_1087;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_1086;
wire n_796;
wire n_1619;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_585;
wire n_1739;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_575;
wire n_480;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1642;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_313),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_243),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_113),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_328),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_207),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_430),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_427),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_327),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_62),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_237),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_3),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_246),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_356),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_347),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_121),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_33),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_134),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_215),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_191),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_226),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_21),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_238),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_245),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_154),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_6),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_270),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_116),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_19),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_429),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_110),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_47),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_16),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_422),
.Y(n_479)
);

BUFx4f_ASAP7_75t_SL g480 ( 
.A(n_319),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_48),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_208),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_176),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_434),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_350),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_209),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_310),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_69),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_411),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_113),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_386),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_433),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_281),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_446),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_261),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_37),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_406),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_54),
.Y(n_498)
);

INVxp33_ASAP7_75t_L g499 ( 
.A(n_212),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_314),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_289),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_138),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_53),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_210),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_230),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_219),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_102),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_267),
.Y(n_508)
);

BUFx10_ASAP7_75t_L g509 ( 
.A(n_194),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_165),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_83),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_143),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_234),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_318),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_378),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_277),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_21),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_432),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_11),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_188),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_200),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_117),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_44),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_425),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_54),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_178),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_216),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_244),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_385),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_346),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_444),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_235),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_320),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_441),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_89),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_391),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_92),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_63),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_345),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_90),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_16),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_428),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_129),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_280),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_8),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g546 ( 
.A(n_423),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_64),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_85),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_338),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_96),
.Y(n_550)
);

CKINVDCx16_ASAP7_75t_R g551 ( 
.A(n_46),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_201),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_442),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_20),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_424),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_150),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_362),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_410),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_436),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_291),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_288),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_374),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_324),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_431),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_155),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_413),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_418),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_123),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_240),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_248),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_110),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_37),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_46),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_273),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_298),
.Y(n_575)
);

CKINVDCx16_ASAP7_75t_R g576 ( 
.A(n_44),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_124),
.Y(n_577)
);

BUFx10_ASAP7_75t_L g578 ( 
.A(n_242),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_268),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_184),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_340),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_315),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_89),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_365),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_11),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_198),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_20),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_8),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_232),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_185),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_58),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_335),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_387),
.Y(n_593)
);

CKINVDCx16_ASAP7_75t_R g594 ( 
.A(n_22),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_256),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_421),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_70),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_321),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_73),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_426),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_239),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_199),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_332),
.Y(n_603)
);

BUFx10_ASAP7_75t_L g604 ( 
.A(n_330),
.Y(n_604)
);

CKINVDCx11_ASAP7_75t_R g605 ( 
.A(n_375),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_260),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_296),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_241),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_122),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_133),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_148),
.Y(n_611)
);

CKINVDCx14_ASAP7_75t_R g612 ( 
.A(n_55),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_250),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_228),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_272),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_153),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_25),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_128),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_155),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_285),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_351),
.Y(n_621)
);

BUFx10_ASAP7_75t_L g622 ( 
.A(n_304),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_0),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_6),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_0),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_618),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_512),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_618),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_454),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_467),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_502),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_535),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_459),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_538),
.Y(n_634)
);

INVxp67_ASAP7_75t_SL g635 ( 
.A(n_512),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_540),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_503),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_541),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_597),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_447),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_599),
.Y(n_641)
);

INVxp67_ASAP7_75t_SL g642 ( 
.A(n_572),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_483),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_619),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_505),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_524),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_572),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_539),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_460),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_544),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_544),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_596),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_457),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_596),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_549),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_450),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_511),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_509),
.Y(n_658)
);

INVxp67_ASAP7_75t_SL g659 ( 
.A(n_537),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_451),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_452),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_520),
.Y(n_662)
);

CKINVDCx16_ASAP7_75t_R g663 ( 
.A(n_551),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_449),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_448),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_456),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_509),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_520),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_465),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_477),
.Y(n_670)
);

BUFx2_ASAP7_75t_SL g671 ( 
.A(n_598),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_466),
.Y(n_672)
);

CKINVDCx16_ASAP7_75t_R g673 ( 
.A(n_576),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_509),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_520),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_487),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_458),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_559),
.Y(n_678)
);

INVxp67_ASAP7_75t_SL g679 ( 
.A(n_609),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_493),
.Y(n_680)
);

CKINVDCx16_ASAP7_75t_R g681 ( 
.A(n_594),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_464),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_497),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_578),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_468),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_471),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_563),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_578),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_564),
.Y(n_689)
);

INVxp33_ASAP7_75t_SL g690 ( 
.A(n_455),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_611),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_550),
.Y(n_692)
);

CKINVDCx16_ASAP7_75t_R g693 ( 
.A(n_612),
.Y(n_693)
);

CKINVDCx16_ASAP7_75t_R g694 ( 
.A(n_612),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_567),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_515),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_520),
.Y(n_697)
);

INVxp67_ASAP7_75t_SL g698 ( 
.A(n_453),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_521),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_472),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_527),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_453),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_531),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_532),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_533),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_475),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_542),
.Y(n_707)
);

INVxp67_ASAP7_75t_SL g708 ( 
.A(n_469),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_479),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_552),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_553),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_668),
.Y(n_712)
);

INVx5_ASAP7_75t_L g713 ( 
.A(n_662),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_671),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_662),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_675),
.Y(n_716)
);

OA21x2_ASAP7_75t_L g717 ( 
.A1(n_697),
.A2(n_489),
.B(n_469),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_662),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_640),
.B(n_613),
.Y(n_719)
);

AOI22x1_ASAP7_75t_SL g720 ( 
.A1(n_629),
.A2(n_571),
.B1(n_470),
.B2(n_517),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_658),
.B(n_534),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_658),
.B(n_546),
.Y(n_722)
);

OA21x2_ASAP7_75t_L g723 ( 
.A1(n_698),
.A2(n_603),
.B(n_489),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_702),
.Y(n_724)
);

OAI21x1_ASAP7_75t_L g725 ( 
.A1(n_704),
.A2(n_699),
.B(n_696),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_662),
.Y(n_726)
);

OA21x2_ASAP7_75t_L g727 ( 
.A1(n_698),
.A2(n_560),
.B(n_555),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_647),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_691),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_665),
.B(n_566),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_SL g731 ( 
.A1(n_692),
.A2(n_571),
.B1(n_470),
.B2(n_598),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_692),
.A2(n_653),
.B1(n_694),
.B2(n_693),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_684),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_677),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_636),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_682),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_685),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_638),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_654),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_708),
.B(n_690),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_667),
.B(n_688),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_654),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_667),
.B(n_570),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_627),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_700),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_630),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_656),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_708),
.B(n_637),
.Y(n_748)
);

AND2x2_ASAP7_75t_SL g749 ( 
.A(n_663),
.B(n_581),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_673),
.A2(n_608),
.B1(n_569),
.B2(n_462),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_660),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_631),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_706),
.B(n_593),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_627),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_661),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_691),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_666),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_635),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_669),
.Y(n_759)
);

OAI21x1_ASAP7_75t_L g760 ( 
.A1(n_672),
.A2(n_606),
.B(n_602),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_632),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_637),
.A2(n_499),
.B1(n_463),
.B2(n_473),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_688),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_676),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_680),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_734),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_712),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_725),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_733),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_712),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_736),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_736),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_714),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_716),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_714),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_746),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_745),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_746),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_737),
.Y(n_779)
);

INVx8_ASAP7_75t_L g780 ( 
.A(n_721),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_746),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_752),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_737),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_739),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_763),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_741),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_740),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_750),
.Y(n_788)
);

CKINVDCx16_ASAP7_75t_R g789 ( 
.A(n_732),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_716),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_752),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_752),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_740),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_720),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_R g795 ( 
.A(n_739),
.B(n_709),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_741),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_719),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_715),
.Y(n_798)
);

CKINVDCx16_ASAP7_75t_R g799 ( 
.A(n_721),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_749),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_729),
.B(n_681),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_R g802 ( 
.A(n_742),
.B(n_633),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_749),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_730),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_761),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_761),
.Y(n_806)
);

CKINVDCx16_ASAP7_75t_R g807 ( 
.A(n_731),
.Y(n_807)
);

INVxp67_ASAP7_75t_L g808 ( 
.A(n_748),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_753),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_742),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_744),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_724),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_R g813 ( 
.A(n_754),
.B(n_643),
.Y(n_813)
);

AND3x1_ASAP7_75t_L g814 ( 
.A(n_748),
.B(n_674),
.C(n_628),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_747),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_747),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_758),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_751),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_762),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_722),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_722),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_743),
.Y(n_822)
);

INVxp67_ASAP7_75t_SL g823 ( 
.A(n_715),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_729),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_755),
.Y(n_825)
);

NOR2xp67_ASAP7_75t_L g826 ( 
.A(n_756),
.B(n_664),
.Y(n_826)
);

BUFx8_ASAP7_75t_L g827 ( 
.A(n_743),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_756),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_715),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_735),
.Y(n_830)
);

AO21x2_ASAP7_75t_L g831 ( 
.A1(n_760),
.A2(n_620),
.B(n_683),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_735),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_804),
.A2(n_608),
.B1(n_646),
.B2(n_645),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_809),
.B(n_686),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_766),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_828),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_784),
.B(n_755),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_786),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_767),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_810),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_808),
.B(n_723),
.Y(n_841)
);

AND2x2_ASAP7_75t_SL g842 ( 
.A(n_807),
.B(n_648),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_769),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_816),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_826),
.B(n_657),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_811),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_771),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_768),
.A2(n_727),
.B1(n_723),
.B2(n_657),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_830),
.Y(n_849)
);

INVx4_ASAP7_75t_L g850 ( 
.A(n_832),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_770),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_787),
.B(n_659),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_824),
.Y(n_853)
);

INVx4_ASAP7_75t_L g854 ( 
.A(n_780),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_797),
.B(n_536),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_784),
.B(n_727),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_817),
.B(n_655),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_793),
.B(n_678),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_818),
.Y(n_859)
);

INVx4_ASAP7_75t_L g860 ( 
.A(n_780),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_780),
.Y(n_861)
);

AND2x6_ASAP7_75t_L g862 ( 
.A(n_801),
.B(n_626),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_785),
.B(n_687),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_776),
.B(n_727),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_796),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_825),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_820),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_774),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_778),
.B(n_765),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_790),
.Y(n_870)
);

XOR2xp5_ASAP7_75t_L g871 ( 
.A(n_788),
.B(n_689),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_798),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_827),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_812),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_799),
.B(n_659),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_773),
.B(n_679),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_781),
.B(n_757),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_831),
.A2(n_499),
.B1(n_717),
.B2(n_679),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_782),
.B(n_759),
.Y(n_879)
);

INVx5_ASAP7_75t_L g880 ( 
.A(n_829),
.Y(n_880)
);

OR2x6_ASAP7_75t_L g881 ( 
.A(n_827),
.B(n_651),
.Y(n_881)
);

INVx5_ASAP7_75t_L g882 ( 
.A(n_829),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_822),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_821),
.B(n_695),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_791),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_802),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_775),
.B(n_777),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_792),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_779),
.B(n_605),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_805),
.B(n_806),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_783),
.B(n_605),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_813),
.Y(n_892)
);

OR2x6_ASAP7_75t_SL g893 ( 
.A(n_772),
.B(n_461),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_819),
.B(n_565),
.Y(n_894)
);

AO22x2_ASAP7_75t_L g895 ( 
.A1(n_789),
.A2(n_800),
.B1(n_803),
.B2(n_814),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_823),
.B(n_474),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_795),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_802),
.B(n_476),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_794),
.B(n_649),
.Y(n_899)
);

BUFx10_ASAP7_75t_L g900 ( 
.A(n_766),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_780),
.Y(n_901)
);

BUFx10_ASAP7_75t_L g902 ( 
.A(n_766),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_828),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_828),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_830),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_826),
.B(n_670),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_815),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_766),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_766),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_815),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_786),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_780),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_766),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_767),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_780),
.Y(n_915)
);

INVx4_ASAP7_75t_L g916 ( 
.A(n_830),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_767),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_826),
.Y(n_918)
);

AND2x6_ASAP7_75t_L g919 ( 
.A(n_768),
.B(n_650),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_766),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_815),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_824),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_766),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_804),
.B(n_478),
.Y(n_924)
);

AND2x6_ASAP7_75t_L g925 ( 
.A(n_768),
.B(n_652),
.Y(n_925)
);

INVx8_ASAP7_75t_L g926 ( 
.A(n_780),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_784),
.B(n_764),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_837),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_843),
.Y(n_929)
);

NOR3xp33_ASAP7_75t_L g930 ( 
.A(n_894),
.B(n_670),
.C(n_639),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_835),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_837),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_927),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_927),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_862),
.A2(n_482),
.B1(n_485),
.B2(n_484),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_834),
.B(n_481),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_875),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_868),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_SL g939 ( 
.A1(n_871),
.A2(n_545),
.B1(n_568),
.B2(n_523),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_870),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_851),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_844),
.Y(n_942)
);

AO22x2_ASAP7_75t_L g943 ( 
.A1(n_852),
.A2(n_642),
.B1(n_703),
.B2(n_701),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_859),
.Y(n_944)
);

AND2x6_ASAP7_75t_L g945 ( 
.A(n_897),
.B(n_705),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_866),
.Y(n_946)
);

OAI22xp33_ASAP7_75t_SL g947 ( 
.A1(n_855),
.A2(n_490),
.B1(n_496),
.B2(n_488),
.Y(n_947)
);

AO22x2_ASAP7_75t_L g948 ( 
.A1(n_857),
.A2(n_710),
.B1(n_711),
.B2(n_707),
.Y(n_948)
);

NAND2x1p5_ASAP7_75t_L g949 ( 
.A(n_901),
.B(n_728),
.Y(n_949)
);

NAND2x1p5_ASAP7_75t_L g950 ( 
.A(n_901),
.B(n_738),
.Y(n_950)
);

NAND3xp33_ASAP7_75t_L g951 ( 
.A(n_924),
.B(n_507),
.C(n_498),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_907),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_912),
.B(n_634),
.Y(n_953)
);

INVxp67_ASAP7_75t_L g954 ( 
.A(n_906),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_910),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_846),
.B(n_519),
.Y(n_956)
);

BUFx8_ASAP7_75t_L g957 ( 
.A(n_922),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_841),
.B(n_738),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_876),
.Y(n_959)
);

OAI221xp5_ASAP7_75t_L g960 ( 
.A1(n_918),
.A2(n_543),
.B1(n_547),
.B2(n_525),
.C(n_522),
.Y(n_960)
);

AO22x2_ASAP7_75t_L g961 ( 
.A1(n_853),
.A2(n_644),
.B1(n_641),
.B2(n_12),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_858),
.B(n_548),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_921),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_914),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_SL g965 ( 
.A(n_908),
.B(n_578),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_879),
.Y(n_966)
);

NAND2x1p5_ASAP7_75t_L g967 ( 
.A(n_912),
.B(n_915),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_879),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_869),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_917),
.Y(n_970)
);

OR2x2_ASAP7_75t_SL g971 ( 
.A(n_903),
.B(n_604),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_909),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_856),
.A2(n_604),
.B1(n_622),
.B2(n_480),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_833),
.B(n_554),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_877),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_896),
.A2(n_491),
.B(n_492),
.C(n_486),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_912),
.B(n_715),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_892),
.B(n_556),
.Y(n_978)
);

NAND2x1p5_ASAP7_75t_L g979 ( 
.A(n_915),
.B(n_718),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_SL g980 ( 
.A(n_913),
.B(n_604),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_836),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_848),
.B(n_494),
.Y(n_982)
);

NAND2x1p5_ASAP7_75t_L g983 ( 
.A(n_915),
.B(n_718),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_849),
.B(n_495),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_904),
.B(n_573),
.Y(n_985)
);

AO22x2_ASAP7_75t_L g986 ( 
.A1(n_884),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_849),
.B(n_577),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_911),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_838),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_878),
.B(n_888),
.Y(n_990)
);

OAI221xp5_ASAP7_75t_L g991 ( 
.A1(n_898),
.A2(n_587),
.B1(n_588),
.B2(n_585),
.C(n_583),
.Y(n_991)
);

CKINVDCx20_ASAP7_75t_R g992 ( 
.A(n_920),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_883),
.Y(n_993)
);

OR2x6_ASAP7_75t_L g994 ( 
.A(n_926),
.B(n_718),
.Y(n_994)
);

INVx8_ASAP7_75t_L g995 ( 
.A(n_926),
.Y(n_995)
);

INVxp67_ASAP7_75t_L g996 ( 
.A(n_887),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_854),
.B(n_164),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_923),
.Y(n_998)
);

NAND2x1p5_ASAP7_75t_L g999 ( 
.A(n_854),
.B(n_860),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_874),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_860),
.B(n_861),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_850),
.B(n_166),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_850),
.B(n_591),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_883),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_883),
.Y(n_1005)
);

NAND3x1_ASAP7_75t_L g1006 ( 
.A(n_863),
.B(n_622),
.C(n_610),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_905),
.B(n_500),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_905),
.B(n_501),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_890),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_862),
.B(n_504),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_916),
.B(n_167),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_885),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_873),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_872),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_872),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_886),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_899),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_865),
.Y(n_1018)
);

OAI221xp5_ASAP7_75t_L g1019 ( 
.A1(n_889),
.A2(n_623),
.B1(n_624),
.B2(n_617),
.C(n_616),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_864),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_895),
.A2(n_919),
.B1(n_925),
.B2(n_840),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_891),
.B(n_625),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_880),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_880),
.Y(n_1024)
);

INVxp67_ASAP7_75t_L g1025 ( 
.A(n_867),
.Y(n_1025)
);

NAND2x1p5_ASAP7_75t_L g1026 ( 
.A(n_880),
.B(n_882),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_847),
.B(n_506),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_882),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_881),
.B(n_168),
.Y(n_1029)
);

OAI221xp5_ASAP7_75t_L g1030 ( 
.A1(n_881),
.A2(n_513),
.B1(n_514),
.B2(n_510),
.C(n_508),
.Y(n_1030)
);

INVx1_ASAP7_75t_SL g1031 ( 
.A(n_900),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_900),
.B(n_516),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_919),
.B(n_518),
.Y(n_1033)
);

NAND2x1p5_ASAP7_75t_L g1034 ( 
.A(n_882),
.B(n_718),
.Y(n_1034)
);

NAND2x1p5_ASAP7_75t_L g1035 ( 
.A(n_842),
.B(n_726),
.Y(n_1035)
);

NAND2x1p5_ASAP7_75t_L g1036 ( 
.A(n_902),
.B(n_726),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_902),
.B(n_622),
.Y(n_1037)
);

AO22x2_ASAP7_75t_L g1038 ( 
.A1(n_895),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_925),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_893),
.B(n_526),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_925),
.Y(n_1041)
);

NAND2x1p5_ASAP7_75t_L g1042 ( 
.A(n_925),
.B(n_726),
.Y(n_1042)
);

BUFx8_ASAP7_75t_L g1043 ( 
.A(n_922),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_843),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_843),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_894),
.B(n_528),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_837),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_837),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_894),
.B(n_529),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_843),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_845),
.B(n_530),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_837),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_839),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_843),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_901),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_901),
.B(n_169),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_894),
.B(n_557),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_894),
.A2(n_561),
.B1(n_562),
.B2(n_558),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_837),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_837),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_901),
.B(n_170),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_839),
.Y(n_1062)
);

INVxp67_ASAP7_75t_L g1063 ( 
.A(n_875),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1020),
.A2(n_575),
.B(n_574),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1049),
.B(n_579),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_1055),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_959),
.B(n_580),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_990),
.A2(n_584),
.B(n_582),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_982),
.A2(n_713),
.B(n_589),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1057),
.B(n_954),
.Y(n_1070)
);

BUFx12f_ASAP7_75t_L g1071 ( 
.A(n_957),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_969),
.B(n_586),
.Y(n_1072)
);

AOI22x1_ASAP7_75t_L g1073 ( 
.A1(n_1039),
.A2(n_592),
.B1(n_595),
.B2(n_590),
.Y(n_1073)
);

INVxp67_ASAP7_75t_L g1074 ( 
.A(n_1050),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_975),
.B(n_600),
.Y(n_1075)
);

NOR2xp67_ASAP7_75t_L g1076 ( 
.A(n_931),
.B(n_601),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1051),
.B(n_607),
.Y(n_1077)
);

INVx11_ASAP7_75t_L g1078 ( 
.A(n_1043),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_937),
.B(n_614),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_1001),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_962),
.B(n_615),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_1044),
.B(n_621),
.Y(n_1082)
);

BUFx8_ASAP7_75t_L g1083 ( 
.A(n_988),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_974),
.A2(n_9),
.B(n_5),
.C(n_7),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_942),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1022),
.A2(n_713),
.B1(n_172),
.B2(n_173),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1041),
.A2(n_174),
.B(n_171),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_1055),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1033),
.A2(n_177),
.B(n_175),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_929),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_941),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_991),
.A2(n_14),
.B(n_10),
.C(n_13),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1010),
.A2(n_180),
.B(n_179),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_1045),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_947),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_1095)
);

INVxp67_ASAP7_75t_L g1096 ( 
.A(n_989),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1021),
.A2(n_182),
.B1(n_183),
.B2(n_181),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1063),
.B(n_15),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_1054),
.B(n_928),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_SL g1100 ( 
.A1(n_976),
.A2(n_187),
.B(n_189),
.C(n_186),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_944),
.B(n_17),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_946),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_952),
.B(n_17),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_SL g1104 ( 
.A(n_965),
.B(n_18),
.C(n_19),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_955),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_993),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_963),
.B(n_18),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_932),
.B(n_22),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_1014),
.Y(n_1109)
);

OR2x6_ASAP7_75t_L g1110 ( 
.A(n_995),
.B(n_23),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_933),
.A2(n_192),
.B1(n_193),
.B2(n_190),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_1017),
.B(n_24),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_938),
.A2(n_196),
.B(n_195),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_1004),
.B(n_197),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_L g1115 ( 
.A(n_936),
.B(n_25),
.C(n_26),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_995),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_966),
.A2(n_968),
.B(n_997),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_997),
.A2(n_203),
.B(n_202),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_934),
.A2(n_205),
.B1(n_206),
.B2(n_204),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_972),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1047),
.B(n_1048),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1052),
.B(n_26),
.Y(n_1122)
);

AO21x2_ASAP7_75t_L g1123 ( 
.A1(n_940),
.A2(n_213),
.B(n_211),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_996),
.B(n_27),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_964),
.Y(n_1125)
);

O2A1O1Ixp33_ASAP7_75t_SL g1126 ( 
.A1(n_1015),
.A2(n_217),
.B(n_218),
.C(n_214),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_930),
.B(n_28),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1059),
.B(n_1060),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_1016),
.B(n_29),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_978),
.B(n_29),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_998),
.B(n_220),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_992),
.Y(n_1132)
);

BUFx12f_ASAP7_75t_L g1133 ( 
.A(n_1013),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_1002),
.B(n_1011),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_1002),
.B(n_221),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_945),
.B(n_30),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_945),
.B(n_30),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1027),
.B(n_31),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_970),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1009),
.A2(n_223),
.B1(n_224),
.B2(n_222),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_985),
.B(n_31),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_1005),
.B(n_225),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1019),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_999),
.A2(n_229),
.B(n_227),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1000),
.A2(n_233),
.B1(n_236),
.B2(n_231),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_1013),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_945),
.B(n_32),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_1018),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_981),
.B(n_34),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_987),
.B(n_35),
.Y(n_1150)
);

NAND3xp33_ASAP7_75t_L g1151 ( 
.A(n_1058),
.B(n_35),
.C(n_36),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1003),
.A2(n_39),
.B(n_36),
.C(n_38),
.Y(n_1152)
);

BUFx4f_ASAP7_75t_L g1153 ( 
.A(n_967),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_1031),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1053),
.A2(n_1062),
.B(n_1042),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_956),
.B(n_38),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_943),
.B(n_39),
.Y(n_1157)
);

NOR2xp67_ASAP7_75t_L g1158 ( 
.A(n_1025),
.B(n_247),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_953),
.B(n_249),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1056),
.A2(n_252),
.B(n_251),
.Y(n_1160)
);

OR2x6_ASAP7_75t_SL g1161 ( 
.A(n_951),
.B(n_40),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_1035),
.B(n_40),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_943),
.B(n_41),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_948),
.A2(n_960),
.B1(n_1012),
.B2(n_1038),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1061),
.A2(n_254),
.B(n_253),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1023),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1061),
.A2(n_257),
.B(n_255),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1024),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_973),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1028),
.Y(n_1170)
);

INVx6_ASAP7_75t_L g1171 ( 
.A(n_953),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1011),
.A2(n_935),
.B1(n_949),
.B2(n_948),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1032),
.B(n_1037),
.Y(n_1173)
);

NOR3xp33_ASAP7_75t_L g1174 ( 
.A(n_939),
.B(n_1030),
.C(n_1040),
.Y(n_1174)
);

AO21x1_ASAP7_75t_L g1175 ( 
.A1(n_984),
.A2(n_42),
.B(n_43),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_950),
.A2(n_259),
.B(n_258),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1007),
.A2(n_48),
.B(n_45),
.C(n_47),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_1008),
.B(n_45),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1026),
.A2(n_263),
.B(n_262),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_980),
.B(n_1036),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_994),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_986),
.B(n_49),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_961),
.B(n_50),
.Y(n_1183)
);

NAND3xp33_ASAP7_75t_L g1184 ( 
.A(n_1029),
.B(n_51),
.C(n_52),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_977),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_979),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1038),
.B(n_51),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_961),
.B(n_52),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_983),
.B(n_53),
.Y(n_1189)
);

AND2x2_ASAP7_75t_SL g1190 ( 
.A(n_971),
.B(n_55),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_994),
.B(n_56),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1034),
.A2(n_265),
.B(n_264),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1006),
.B(n_57),
.Y(n_1193)
);

AOI21xp33_ASAP7_75t_L g1194 ( 
.A1(n_1046),
.A2(n_57),
.B(n_58),
.Y(n_1194)
);

INVxp67_ASAP7_75t_L g1195 ( 
.A(n_1050),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_959),
.B(n_59),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1046),
.B(n_59),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1046),
.B(n_60),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_959),
.B(n_60),
.Y(n_1199)
);

AOI21x1_ASAP7_75t_L g1200 ( 
.A1(n_958),
.A2(n_269),
.B(n_266),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1046),
.A2(n_63),
.B(n_61),
.C(n_62),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1050),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_959),
.B(n_61),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1085),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1173),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1102),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_1154),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1070),
.B(n_65),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1074),
.B(n_66),
.Y(n_1209)
);

INVx4_ASAP7_75t_L g1210 ( 
.A(n_1133),
.Y(n_1210)
);

NOR2x1_ASAP7_75t_L g1211 ( 
.A(n_1132),
.B(n_271),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1105),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1066),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1138),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1202),
.B(n_71),
.Y(n_1215)
);

INVxp67_ASAP7_75t_L g1216 ( 
.A(n_1094),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1134),
.B(n_72),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1072),
.B(n_72),
.Y(n_1218)
);

OA22x2_ASAP7_75t_L g1219 ( 
.A1(n_1183),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1195),
.B(n_75),
.Y(n_1220)
);

OA22x2_ASAP7_75t_L g1221 ( 
.A1(n_1110),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1156),
.B(n_76),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1075),
.B(n_77),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1066),
.Y(n_1224)
);

INVxp67_ASAP7_75t_L g1225 ( 
.A(n_1106),
.Y(n_1225)
);

OAI21xp33_ASAP7_75t_L g1226 ( 
.A1(n_1197),
.A2(n_78),
.B(n_79),
.Y(n_1226)
);

BUFx12f_ASAP7_75t_L g1227 ( 
.A(n_1071),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1096),
.B(n_80),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_1120),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1081),
.B(n_80),
.Y(n_1230)
);

NOR3xp33_ASAP7_75t_SL g1231 ( 
.A(n_1104),
.B(n_81),
.C(n_82),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1198),
.B(n_81),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1116),
.B(n_445),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1150),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_1234)
);

AOI21xp33_ASAP7_75t_L g1235 ( 
.A1(n_1065),
.A2(n_85),
.B(n_86),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1117),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1083),
.Y(n_1237)
);

NAND2xp33_ASAP7_75t_L g1238 ( 
.A(n_1130),
.B(n_274),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1077),
.A2(n_276),
.B(n_275),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1090),
.B(n_91),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1164),
.B(n_91),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1083),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1141),
.B(n_92),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1172),
.A2(n_279),
.B(n_278),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1153),
.B(n_93),
.Y(n_1245)
);

NOR3xp33_ASAP7_75t_L g1246 ( 
.A(n_1174),
.B(n_94),
.C(n_95),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1113),
.A2(n_96),
.B(n_94),
.C(n_95),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1153),
.B(n_97),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1146),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1151),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1095),
.A2(n_100),
.B(n_98),
.C(n_99),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1116),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_1148),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1155),
.A2(n_283),
.B(n_282),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1088),
.B(n_1076),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1101),
.B(n_101),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1069),
.A2(n_286),
.B(n_284),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1135),
.A2(n_1087),
.B(n_1089),
.Y(n_1258)
);

OAI21xp33_ASAP7_75t_SL g1259 ( 
.A1(n_1103),
.A2(n_103),
.B(n_104),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1080),
.Y(n_1260)
);

AO21x1_ASAP7_75t_L g1261 ( 
.A1(n_1097),
.A2(n_105),
.B(n_106),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1088),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1194),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1171),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_1264)
);

O2A1O1Ixp33_ASAP7_75t_SL g1265 ( 
.A1(n_1169),
.A2(n_339),
.B(n_440),
.C(n_439),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1171),
.B(n_108),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1116),
.B(n_287),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1180),
.B(n_109),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1107),
.B(n_111),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1196),
.B(n_111),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1199),
.B(n_112),
.Y(n_1271)
);

AO22x1_ASAP7_75t_L g1272 ( 
.A1(n_1159),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1064),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_SL g1274 ( 
.A(n_1190),
.B(n_290),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1159),
.B(n_117),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1114),
.B(n_118),
.Y(n_1276)
);

NOR3xp33_ASAP7_75t_SL g1277 ( 
.A(n_1193),
.B(n_118),
.C(n_119),
.Y(n_1277)
);

OR2x6_ASAP7_75t_SL g1278 ( 
.A(n_1184),
.B(n_119),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1109),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1203),
.B(n_120),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1091),
.B(n_120),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1078),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1127),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1166),
.B(n_292),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1067),
.B(n_124),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1092),
.A2(n_1143),
.B(n_1068),
.C(n_1160),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1079),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1093),
.A2(n_294),
.B(n_293),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1114),
.B(n_125),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1124),
.B(n_126),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1142),
.B(n_295),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1165),
.A2(n_128),
.B(n_129),
.C(n_130),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1167),
.A2(n_130),
.B(n_131),
.C(n_132),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_R g1294 ( 
.A(n_1109),
.B(n_297),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1125),
.B(n_131),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1158),
.B(n_133),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1098),
.B(n_134),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1168),
.B(n_135),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1084),
.A2(n_135),
.B(n_136),
.C(n_137),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1118),
.A2(n_300),
.B(n_299),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1139),
.B(n_136),
.Y(n_1301)
);

NAND2xp33_ASAP7_75t_SL g1302 ( 
.A(n_1178),
.B(n_137),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1112),
.B(n_1161),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1099),
.B(n_139),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1108),
.B(n_140),
.Y(n_1305)
);

A2O1A1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1115),
.A2(n_141),
.B(n_142),
.C(n_143),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1170),
.B(n_141),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1181),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_SL g1309 ( 
.A1(n_1177),
.A2(n_370),
.B(n_438),
.C(n_437),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1122),
.B(n_142),
.Y(n_1310)
);

OAI21xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1121),
.A2(n_144),
.B(n_145),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1185),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1162),
.Y(n_1313)
);

CKINVDCx12_ASAP7_75t_R g1314 ( 
.A(n_1110),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1186),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1200),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1149),
.B(n_1128),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1201),
.A2(n_144),
.B(n_145),
.C(n_146),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1082),
.B(n_146),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1157),
.B(n_147),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1163),
.B(n_1182),
.Y(n_1321)
);

NAND2x1_ASAP7_75t_L g1322 ( 
.A(n_1144),
.B(n_301),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1123),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1129),
.B(n_147),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1187),
.B(n_148),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1189),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1175),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1191),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1086),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1188),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1152),
.B(n_149),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1131),
.Y(n_1332)
);

BUFx8_ASAP7_75t_L g1333 ( 
.A(n_1136),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1137),
.B(n_151),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1147),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1123),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1111),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1119),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1179),
.B(n_156),
.Y(n_1339)
);

NOR2x1_ASAP7_75t_R g1340 ( 
.A(n_1073),
.B(n_302),
.Y(n_1340)
);

BUFx12f_ASAP7_75t_L g1341 ( 
.A(n_1100),
.Y(n_1341)
);

NOR3xp33_ASAP7_75t_SL g1342 ( 
.A(n_1140),
.B(n_157),
.C(n_158),
.Y(n_1342)
);

INVx11_ASAP7_75t_L g1343 ( 
.A(n_1192),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1145),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1176),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1252),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1249),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1204),
.Y(n_1348)
);

INVx5_ASAP7_75t_L g1349 ( 
.A(n_1213),
.Y(n_1349)
);

CKINVDCx16_ASAP7_75t_R g1350 ( 
.A(n_1229),
.Y(n_1350)
);

BUFx4f_ASAP7_75t_L g1351 ( 
.A(n_1227),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1212),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1207),
.Y(n_1353)
);

BUFx12f_ASAP7_75t_L g1354 ( 
.A(n_1282),
.Y(n_1354)
);

INVx4_ASAP7_75t_L g1355 ( 
.A(n_1213),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1213),
.Y(n_1356)
);

BUFx12f_ASAP7_75t_L g1357 ( 
.A(n_1210),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1262),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1206),
.Y(n_1359)
);

BUFx12f_ASAP7_75t_L g1360 ( 
.A(n_1210),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1313),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1216),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1253),
.Y(n_1363)
);

INVxp67_ASAP7_75t_SL g1364 ( 
.A(n_1279),
.Y(n_1364)
);

INVx5_ASAP7_75t_L g1365 ( 
.A(n_1224),
.Y(n_1365)
);

CKINVDCx6p67_ASAP7_75t_R g1366 ( 
.A(n_1237),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1308),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1224),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1333),
.Y(n_1369)
);

BUFx12f_ASAP7_75t_L g1370 ( 
.A(n_1242),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1333),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1224),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1330),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1312),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1312),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1315),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1315),
.B(n_303),
.Y(n_1377)
);

INVxp67_ASAP7_75t_SL g1378 ( 
.A(n_1225),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_1314),
.Y(n_1379)
);

INVx3_ASAP7_75t_SL g1380 ( 
.A(n_1255),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1328),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1332),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1321),
.B(n_1126),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1233),
.Y(n_1384)
);

CKINVDCx6p67_ASAP7_75t_R g1385 ( 
.A(n_1278),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1297),
.B(n_159),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1317),
.B(n_159),
.Y(n_1387)
);

INVx1_ASAP7_75t_SL g1388 ( 
.A(n_1326),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1281),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1267),
.Y(n_1390)
);

OR2x6_ASAP7_75t_L g1391 ( 
.A(n_1291),
.B(n_305),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1295),
.Y(n_1392)
);

INVxp67_ASAP7_75t_SL g1393 ( 
.A(n_1260),
.Y(n_1393)
);

INVx3_ASAP7_75t_SL g1394 ( 
.A(n_1332),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1332),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1324),
.B(n_160),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1303),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1284),
.Y(n_1398)
);

INVx5_ASAP7_75t_L g1399 ( 
.A(n_1260),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1327),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1266),
.Y(n_1401)
);

INVx6_ASAP7_75t_SL g1402 ( 
.A(n_1221),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1209),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1302),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1301),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_SL g1406 ( 
.A(n_1345),
.Y(n_1406)
);

INVx5_ASAP7_75t_L g1407 ( 
.A(n_1341),
.Y(n_1407)
);

NAND2x1p5_ASAP7_75t_L g1408 ( 
.A(n_1211),
.B(n_306),
.Y(n_1408)
);

BUFx12f_ASAP7_75t_L g1409 ( 
.A(n_1339),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1325),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1294),
.Y(n_1411)
);

NAND2x1p5_ASAP7_75t_L g1412 ( 
.A(n_1322),
.B(n_307),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1208),
.B(n_160),
.Y(n_1413)
);

INVx4_ASAP7_75t_L g1414 ( 
.A(n_1343),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_1220),
.Y(n_1415)
);

CKINVDCx6p67_ASAP7_75t_R g1416 ( 
.A(n_1245),
.Y(n_1416)
);

INVxp67_ASAP7_75t_SL g1417 ( 
.A(n_1217),
.Y(n_1417)
);

INVx5_ASAP7_75t_SL g1418 ( 
.A(n_1344),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1316),
.Y(n_1419)
);

BUFx12f_ASAP7_75t_L g1420 ( 
.A(n_1337),
.Y(n_1420)
);

BUFx2_ASAP7_75t_SL g1421 ( 
.A(n_1219),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1275),
.B(n_308),
.Y(n_1422)
);

INVx4_ASAP7_75t_L g1423 ( 
.A(n_1316),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1228),
.Y(n_1424)
);

INVx8_ASAP7_75t_L g1425 ( 
.A(n_1323),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1268),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1320),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1230),
.B(n_161),
.Y(n_1428)
);

BUFx4_ASAP7_75t_SL g1429 ( 
.A(n_1336),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1243),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1246),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_1431)
);

BUFx4f_ASAP7_75t_SL g1432 ( 
.A(n_1215),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1311),
.Y(n_1433)
);

INVx3_ASAP7_75t_L g1434 ( 
.A(n_1218),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1277),
.Y(n_1435)
);

BUFx2_ASAP7_75t_SL g1436 ( 
.A(n_1296),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1304),
.Y(n_1437)
);

CKINVDCx11_ASAP7_75t_R g1438 ( 
.A(n_1335),
.Y(n_1438)
);

INVx3_ASAP7_75t_SL g1439 ( 
.A(n_1240),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1232),
.B(n_162),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1276),
.Y(n_1441)
);

NAND3xp33_ASAP7_75t_L g1442 ( 
.A(n_1290),
.B(n_163),
.C(n_309),
.Y(n_1442)
);

NAND2x1p5_ASAP7_75t_L g1443 ( 
.A(n_1289),
.B(n_311),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1248),
.Y(n_1444)
);

INVx3_ASAP7_75t_SL g1445 ( 
.A(n_1222),
.Y(n_1445)
);

BUFx12f_ASAP7_75t_L g1446 ( 
.A(n_1272),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1338),
.Y(n_1447)
);

INVx5_ASAP7_75t_L g1448 ( 
.A(n_1340),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1286),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1298),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1223),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1285),
.Y(n_1452)
);

INVxp67_ASAP7_75t_L g1453 ( 
.A(n_1307),
.Y(n_1453)
);

BUFx12f_ASAP7_75t_L g1454 ( 
.A(n_1259),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1274),
.A2(n_312),
.B1(n_316),
.B2(n_317),
.Y(n_1455)
);

BUFx8_ASAP7_75t_SL g1456 ( 
.A(n_1270),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_SL g1457 ( 
.A1(n_1329),
.A2(n_322),
.B1(n_323),
.B2(n_325),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1319),
.Y(n_1458)
);

BUFx8_ASAP7_75t_L g1459 ( 
.A(n_1231),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1271),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1241),
.B(n_443),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_1280),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1334),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1305),
.Y(n_1464)
);

OR2x6_ASAP7_75t_L g1465 ( 
.A(n_1244),
.B(n_326),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1310),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1256),
.Y(n_1467)
);

NAND2x1_ASAP7_75t_L g1468 ( 
.A(n_1258),
.B(n_435),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1438),
.A2(n_1273),
.B1(n_1235),
.B2(n_1226),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1361),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1347),
.Y(n_1471)
);

NAND2x1p5_ASAP7_75t_L g1472 ( 
.A(n_1349),
.B(n_1254),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1449),
.A2(n_1261),
.B1(n_1263),
.B2(n_1250),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1468),
.A2(n_1257),
.B(n_1288),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1350),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1452),
.A2(n_1331),
.B1(n_1214),
.B2(n_1283),
.Y(n_1476)
);

O2A1O1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1428),
.A2(n_1247),
.B(n_1251),
.C(n_1234),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1361),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1410),
.B(n_1269),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1458),
.A2(n_1205),
.B1(n_1236),
.B2(n_1287),
.Y(n_1480)
);

NOR2xp67_ASAP7_75t_L g1481 ( 
.A(n_1414),
.B(n_1239),
.Y(n_1481)
);

BUFx12f_ASAP7_75t_L g1482 ( 
.A(n_1354),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1363),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1369),
.Y(n_1484)
);

INVx6_ASAP7_75t_L g1485 ( 
.A(n_1357),
.Y(n_1485)
);

NAND2x1p5_ASAP7_75t_L g1486 ( 
.A(n_1349),
.B(n_1300),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1381),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1367),
.Y(n_1488)
);

A2O1A1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1422),
.A2(n_1299),
.B(n_1318),
.C(n_1342),
.Y(n_1489)
);

OAI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1442),
.A2(n_1293),
.B(n_1292),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1348),
.Y(n_1491)
);

INVx4_ASAP7_75t_SL g1492 ( 
.A(n_1380),
.Y(n_1492)
);

AOI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1404),
.A2(n_1238),
.B1(n_1264),
.B2(n_1306),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1426),
.B(n_329),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1352),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1419),
.A2(n_1265),
.B(n_1309),
.Y(n_1496)
);

INVxp67_ASAP7_75t_SL g1497 ( 
.A(n_1364),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1398),
.B(n_331),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1400),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1400),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1412),
.A2(n_333),
.B(n_334),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1359),
.Y(n_1502)
);

NAND2x1p5_ASAP7_75t_L g1503 ( 
.A(n_1349),
.B(n_336),
.Y(n_1503)
);

INVx3_ASAP7_75t_SL g1504 ( 
.A(n_1366),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1383),
.A2(n_337),
.B(n_341),
.Y(n_1505)
);

BUFx2_ASAP7_75t_SL g1506 ( 
.A(n_1407),
.Y(n_1506)
);

AOI222xp33_ASAP7_75t_L g1507 ( 
.A1(n_1440),
.A2(n_342),
.B1(n_343),
.B2(n_344),
.C1(n_348),
.C2(n_349),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1425),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1374),
.Y(n_1509)
);

BUFx12f_ASAP7_75t_L g1510 ( 
.A(n_1360),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1408),
.A2(n_352),
.B(n_353),
.Y(n_1511)
);

CKINVDCx20_ASAP7_75t_R g1512 ( 
.A(n_1371),
.Y(n_1512)
);

CKINVDCx11_ASAP7_75t_R g1513 ( 
.A(n_1379),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1425),
.Y(n_1514)
);

INVx4_ASAP7_75t_SL g1515 ( 
.A(n_1394),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1346),
.Y(n_1516)
);

AO31x2_ASAP7_75t_L g1517 ( 
.A1(n_1423),
.A2(n_354),
.A3(n_355),
.B(n_357),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1465),
.A2(n_358),
.B(n_359),
.Y(n_1518)
);

OA21x2_ASAP7_75t_L g1519 ( 
.A1(n_1433),
.A2(n_360),
.B(n_361),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1399),
.Y(n_1520)
);

BUFx8_ASAP7_75t_L g1521 ( 
.A(n_1370),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1465),
.A2(n_363),
.B(n_364),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1406),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1460),
.B(n_366),
.Y(n_1524)
);

BUFx12f_ASAP7_75t_L g1525 ( 
.A(n_1373),
.Y(n_1525)
);

OR2x6_ASAP7_75t_L g1526 ( 
.A(n_1391),
.B(n_367),
.Y(n_1526)
);

NAND3xp33_ASAP7_75t_L g1527 ( 
.A(n_1431),
.B(n_368),
.C(n_369),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1446),
.A2(n_371),
.B1(n_372),
.B2(n_373),
.Y(n_1528)
);

AO21x2_ASAP7_75t_L g1529 ( 
.A1(n_1417),
.A2(n_376),
.B(n_377),
.Y(n_1529)
);

AOI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1451),
.A2(n_379),
.B1(n_380),
.B2(n_381),
.Y(n_1530)
);

AO21x2_ASAP7_75t_L g1531 ( 
.A1(n_1389),
.A2(n_382),
.B(n_383),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1358),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1462),
.B(n_384),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_1356),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1453),
.A2(n_388),
.B(n_389),
.Y(n_1535)
);

OR2x6_ASAP7_75t_L g1536 ( 
.A(n_1391),
.B(n_390),
.Y(n_1536)
);

AO21x2_ASAP7_75t_L g1537 ( 
.A1(n_1392),
.A2(n_392),
.B(n_393),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1433),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1410),
.B(n_394),
.Y(n_1539)
);

O2A1O1Ixp33_ASAP7_75t_L g1540 ( 
.A1(n_1413),
.A2(n_395),
.B(n_396),
.C(n_397),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_SL g1541 ( 
.A1(n_1421),
.A2(n_398),
.B1(n_399),
.B2(n_400),
.Y(n_1541)
);

AOI21xp33_ASAP7_75t_L g1542 ( 
.A1(n_1434),
.A2(n_401),
.B(n_402),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1502),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1469),
.A2(n_1437),
.B1(n_1385),
.B2(n_1421),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1523),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1499),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1499),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_SL g1548 ( 
.A1(n_1490),
.A2(n_1454),
.B1(n_1436),
.B2(n_1420),
.Y(n_1548)
);

AO21x1_ASAP7_75t_L g1549 ( 
.A1(n_1477),
.A2(n_1387),
.B(n_1405),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1479),
.B(n_1397),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1500),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1476),
.A2(n_1480),
.B1(n_1489),
.B2(n_1493),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1538),
.B(n_1427),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1488),
.B(n_1467),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1500),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1538),
.B(n_1430),
.Y(n_1556)
);

INVx4_ASAP7_75t_SL g1557 ( 
.A(n_1517),
.Y(n_1557)
);

AO21x1_ASAP7_75t_SL g1558 ( 
.A1(n_1535),
.A2(n_1461),
.B(n_1429),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1470),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1474),
.A2(n_1443),
.B(n_1393),
.Y(n_1560)
);

BUFx12f_ASAP7_75t_L g1561 ( 
.A(n_1513),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1491),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1497),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1495),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_SL g1565 ( 
.A1(n_1519),
.A2(n_1436),
.B1(n_1463),
.B2(n_1459),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1523),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1485),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1473),
.A2(n_1450),
.B1(n_1445),
.B2(n_1459),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1478),
.Y(n_1569)
);

INVx2_ASAP7_75t_SL g1570 ( 
.A(n_1520),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1508),
.B(n_1395),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1519),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1496),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1487),
.Y(n_1574)
);

AOI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1507),
.A2(n_1435),
.B1(n_1416),
.B2(n_1409),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1559),
.B(n_1471),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1569),
.B(n_1508),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1552),
.A2(n_1527),
.B1(n_1536),
.B2(n_1526),
.Y(n_1578)
);

AOI221xp5_ASAP7_75t_L g1579 ( 
.A1(n_1549),
.A2(n_1464),
.B1(n_1466),
.B2(n_1396),
.C(n_1494),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1569),
.B(n_1388),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1546),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1546),
.Y(n_1582)
);

INVxp33_ASAP7_75t_SL g1583 ( 
.A(n_1574),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1570),
.B(n_1514),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1545),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1554),
.B(n_1532),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1563),
.B(n_1447),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1550),
.B(n_1475),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1545),
.B(n_1367),
.Y(n_1589)
);

INVx8_ASAP7_75t_L g1590 ( 
.A(n_1561),
.Y(n_1590)
);

OAI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1575),
.A2(n_1540),
.B(n_1518),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1543),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1561),
.Y(n_1593)
);

AO21x2_ASAP7_75t_L g1594 ( 
.A1(n_1572),
.A2(n_1481),
.B(n_1537),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1566),
.Y(n_1595)
);

BUFx10_ASAP7_75t_L g1596 ( 
.A(n_1567),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_R g1597 ( 
.A(n_1566),
.B(n_1484),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1547),
.B(n_1464),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1562),
.Y(n_1599)
);

NAND2xp33_ASAP7_75t_R g1600 ( 
.A(n_1571),
.B(n_1526),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1553),
.B(n_1492),
.Y(n_1601)
);

NAND2xp33_ASAP7_75t_R g1602 ( 
.A(n_1571),
.B(n_1556),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1547),
.B(n_1466),
.Y(n_1603)
);

NAND2xp33_ASAP7_75t_R g1604 ( 
.A(n_1571),
.B(n_1536),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1543),
.Y(n_1605)
);

OAI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1565),
.A2(n_1522),
.B(n_1530),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1592),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1605),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1605),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1581),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1582),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1576),
.B(n_1551),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1577),
.B(n_1551),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1577),
.B(n_1555),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1580),
.B(n_1562),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1585),
.B(n_1557),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1599),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1593),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1598),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1587),
.B(n_1564),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1584),
.Y(n_1621)
);

OAI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1595),
.A2(n_1573),
.B(n_1560),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1607),
.Y(n_1623)
);

AO21x2_ASAP7_75t_L g1624 ( 
.A1(n_1608),
.A2(n_1594),
.B(n_1597),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1618),
.B(n_1485),
.Y(n_1625)
);

OAI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1619),
.A2(n_1602),
.B1(n_1591),
.B2(n_1600),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1618),
.B(n_1590),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1607),
.Y(n_1628)
);

OAI32xp33_ASAP7_75t_L g1629 ( 
.A1(n_1615),
.A2(n_1604),
.A3(n_1578),
.B1(n_1544),
.B2(n_1583),
.Y(n_1629)
);

AO21x2_ASAP7_75t_L g1630 ( 
.A1(n_1622),
.A2(n_1609),
.B(n_1608),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1623),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1624),
.B(n_1613),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1630),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1628),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1630),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1627),
.Y(n_1636)
);

AND2x4_ASAP7_75t_SL g1637 ( 
.A(n_1632),
.B(n_1596),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1636),
.B(n_1613),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1631),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1636),
.B(n_1626),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1634),
.B(n_1619),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1635),
.B(n_1614),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1633),
.B(n_1614),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1633),
.B(n_1612),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1636),
.B(n_1612),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1634),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1638),
.B(n_1610),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1639),
.Y(n_1648)
);

INVxp67_ASAP7_75t_SL g1649 ( 
.A(n_1640),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1637),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1639),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1641),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1646),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1643),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1645),
.B(n_1625),
.Y(n_1655)
);

OR2x6_ASAP7_75t_L g1656 ( 
.A(n_1644),
.B(n_1590),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1642),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1655),
.B(n_1596),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1650),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1655),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1649),
.B(n_1603),
.Y(n_1661)
);

OA21x2_ASAP7_75t_L g1662 ( 
.A1(n_1648),
.A2(n_1606),
.B(n_1622),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1651),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1654),
.B(n_1620),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1657),
.Y(n_1665)
);

NOR2xp67_ASAP7_75t_L g1666 ( 
.A(n_1659),
.B(n_1652),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1660),
.B(n_1653),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1661),
.B(n_1647),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1665),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1666),
.A2(n_1658),
.B1(n_1656),
.B2(n_1657),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1669),
.Y(n_1671)
);

NAND3xp33_ASAP7_75t_L g1672 ( 
.A(n_1667),
.B(n_1665),
.C(n_1663),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1668),
.Y(n_1673)
);

NAND2x1p5_ASAP7_75t_L g1674 ( 
.A(n_1673),
.B(n_1351),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1672),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1670),
.B(n_1656),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1671),
.B(n_1664),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1673),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1678),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1677),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1675),
.B(n_1662),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1676),
.B(n_1662),
.Y(n_1682)
);

OAI21xp5_ASAP7_75t_SL g1683 ( 
.A1(n_1674),
.A2(n_1528),
.B(n_1353),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1674),
.Y(n_1684)
);

NAND2x1_ASAP7_75t_L g1685 ( 
.A(n_1676),
.B(n_1483),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1678),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1678),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1676),
.B(n_1504),
.Y(n_1688)
);

NAND4xp25_ASAP7_75t_SL g1689 ( 
.A(n_1681),
.B(n_1512),
.C(n_1579),
.D(n_1568),
.Y(n_1689)
);

NAND3xp33_ASAP7_75t_L g1690 ( 
.A(n_1679),
.B(n_1521),
.C(n_1524),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1688),
.B(n_1525),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1682),
.B(n_1588),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1686),
.B(n_1586),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1684),
.B(n_1482),
.Y(n_1694)
);

OAI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1683),
.A2(n_1407),
.B1(n_1510),
.B2(n_1448),
.Y(n_1695)
);

OAI21xp33_ASAP7_75t_L g1696 ( 
.A1(n_1680),
.A2(n_1629),
.B(n_1568),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1687),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_1685),
.Y(n_1698)
);

NAND3xp33_ASAP7_75t_L g1699 ( 
.A(n_1683),
.B(n_1521),
.C(n_1533),
.Y(n_1699)
);

NOR3x1_ASAP7_75t_L g1700 ( 
.A(n_1685),
.B(n_1378),
.C(n_1411),
.Y(n_1700)
);

AOI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1694),
.A2(n_1506),
.B1(n_1492),
.B2(n_1415),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_L g1702 ( 
.A(n_1697),
.B(n_1386),
.C(n_1455),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1698),
.Y(n_1703)
);

AOI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1696),
.A2(n_1629),
.B1(n_1424),
.B2(n_1403),
.C(n_1362),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1689),
.A2(n_1691),
.B1(n_1692),
.B2(n_1690),
.Y(n_1705)
);

AOI221xp5_ASAP7_75t_L g1706 ( 
.A1(n_1695),
.A2(n_1516),
.B1(n_1401),
.B2(n_1544),
.C(n_1439),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1693),
.B(n_1700),
.Y(n_1707)
);

OAI21xp33_ASAP7_75t_L g1708 ( 
.A1(n_1699),
.A2(n_1601),
.B(n_1548),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1694),
.A2(n_1515),
.B1(n_1432),
.B2(n_1407),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1692),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1692),
.B(n_1456),
.Y(n_1711)
);

OAI21xp5_ASAP7_75t_SL g1712 ( 
.A1(n_1694),
.A2(n_1541),
.B(n_1503),
.Y(n_1712)
);

NAND4xp75_ASAP7_75t_L g1713 ( 
.A(n_1710),
.B(n_1539),
.C(n_1542),
.D(n_1515),
.Y(n_1713)
);

AOI221xp5_ASAP7_75t_L g1714 ( 
.A1(n_1703),
.A2(n_1444),
.B1(n_1611),
.B2(n_1498),
.C(n_1441),
.Y(n_1714)
);

AOI211xp5_ASAP7_75t_L g1715 ( 
.A1(n_1707),
.A2(n_1498),
.B(n_1377),
.C(n_1444),
.Y(n_1715)
);

NOR3xp33_ASAP7_75t_L g1716 ( 
.A(n_1711),
.B(n_1377),
.C(n_1382),
.Y(n_1716)
);

NOR3xp33_ASAP7_75t_L g1717 ( 
.A(n_1705),
.B(n_1355),
.C(n_1457),
.Y(n_1717)
);

AOI211xp5_ASAP7_75t_L g1718 ( 
.A1(n_1701),
.A2(n_1441),
.B(n_1374),
.C(n_1376),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_R g1719 ( 
.A(n_1709),
.B(n_403),
.Y(n_1719)
);

AO22x2_ASAP7_75t_L g1720 ( 
.A1(n_1702),
.A2(n_1557),
.B1(n_1509),
.B2(n_1611),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1708),
.A2(n_1448),
.B(n_1529),
.Y(n_1721)
);

XNOR2xp5_ASAP7_75t_L g1722 ( 
.A(n_1706),
.B(n_1384),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1704),
.B(n_1589),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1723),
.Y(n_1724)
);

A2O1A1Ixp33_ASAP7_75t_L g1725 ( 
.A1(n_1721),
.A2(n_1712),
.B(n_1616),
.C(n_1448),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1717),
.B(n_1715),
.Y(n_1726)
);

NAND2x2_ASAP7_75t_L g1727 ( 
.A(n_1719),
.B(n_1390),
.Y(n_1727)
);

AND3x4_ASAP7_75t_L g1728 ( 
.A(n_1716),
.B(n_1616),
.C(n_1584),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1718),
.B(n_1418),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1720),
.Y(n_1730)
);

AOI21xp33_ASAP7_75t_SL g1731 ( 
.A1(n_1722),
.A2(n_404),
.B(n_405),
.Y(n_1731)
);

AOI22x1_ASAP7_75t_L g1732 ( 
.A1(n_1720),
.A2(n_1713),
.B1(n_1714),
.B2(n_1368),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1723),
.B(n_1375),
.Y(n_1733)
);

NOR2x1_ASAP7_75t_L g1734 ( 
.A(n_1713),
.B(n_1537),
.Y(n_1734)
);

NOR3x1_ASAP7_75t_L g1735 ( 
.A(n_1724),
.B(n_1729),
.C(n_1730),
.Y(n_1735)
);

NAND2x1p5_ASAP7_75t_L g1736 ( 
.A(n_1734),
.B(n_1732),
.Y(n_1736)
);

NOR2x1_ASAP7_75t_L g1737 ( 
.A(n_1725),
.B(n_1531),
.Y(n_1737)
);

NAND5xp2_ASAP7_75t_L g1738 ( 
.A(n_1726),
.B(n_1402),
.C(n_1486),
.D(n_1472),
.E(n_1558),
.Y(n_1738)
);

XNOR2x1_ASAP7_75t_L g1739 ( 
.A(n_1728),
.B(n_407),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1731),
.B(n_1418),
.Y(n_1740)
);

NAND2x1p5_ASAP7_75t_L g1741 ( 
.A(n_1733),
.B(n_1727),
.Y(n_1741)
);

NOR2xp67_ASAP7_75t_L g1742 ( 
.A(n_1731),
.B(n_408),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1724),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1743),
.Y(n_1744)
);

CKINVDCx16_ASAP7_75t_R g1745 ( 
.A(n_1740),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_1735),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_1736),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1739),
.B(n_1617),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1742),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1741),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1738),
.Y(n_1751)
);

AOI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1746),
.A2(n_1737),
.B1(n_1616),
.B2(n_1621),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1747),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1744),
.A2(n_1365),
.B1(n_1402),
.B2(n_1621),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1751),
.A2(n_1365),
.B1(n_1621),
.B2(n_1534),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1747),
.Y(n_1756)
);

XNOR2xp5_ASAP7_75t_L g1757 ( 
.A(n_1750),
.B(n_409),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1749),
.B(n_1376),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1753),
.B(n_1745),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1756),
.B(n_1748),
.Y(n_1760)
);

XNOR2xp5_ASAP7_75t_L g1761 ( 
.A(n_1757),
.B(n_412),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1758),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1752),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1754),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1761),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1759),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1760),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1763),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1762),
.Y(n_1769)
);

CKINVDCx20_ASAP7_75t_R g1770 ( 
.A(n_1764),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1768),
.A2(n_1755),
.B(n_1511),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1767),
.Y(n_1772)
);

XOR2xp5_ASAP7_75t_L g1773 ( 
.A(n_1770),
.B(n_414),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1769),
.Y(n_1774)
);

NOR2xp67_ASAP7_75t_L g1775 ( 
.A(n_1772),
.B(n_1766),
.Y(n_1775)
);

OAI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1774),
.A2(n_1765),
.B1(n_1365),
.B2(n_1372),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1773),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1777),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1775),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1779),
.A2(n_1776),
.B1(n_1771),
.B2(n_1368),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_SL g1781 ( 
.A1(n_1780),
.A2(n_1778),
.B1(n_1356),
.B2(n_1372),
.Y(n_1781)
);

AO21x2_ASAP7_75t_L g1782 ( 
.A1(n_1781),
.A2(n_1501),
.B(n_1505),
.Y(n_1782)
);

AOI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1782),
.A2(n_415),
.B(n_416),
.Y(n_1783)
);

AOI211xp5_ASAP7_75t_L g1784 ( 
.A1(n_1783),
.A2(n_417),
.B(n_419),
.C(n_420),
.Y(n_1784)
);


endmodule