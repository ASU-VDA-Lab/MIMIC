module fake_jpeg_9404_n_45 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_45);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_45;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_29),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_21),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_24),
.C(n_2),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_32),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_12),
.B1(n_17),
.B2(n_16),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_33),
.A2(n_37),
.B(n_10),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_1),
.B(n_2),
.Y(n_41)
);

AND2x6_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_6),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_41),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_39),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_38),
.C(n_35),
.Y(n_44)
);

AOI31xp33_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_36),
.A3(n_3),
.B(n_34),
.Y(n_45)
);


endmodule