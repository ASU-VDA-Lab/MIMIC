module fake_netlist_6_452_n_1080 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1080);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1080;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_1008;
wire n_760;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_758;
wire n_720;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_870;
wire n_904;
wire n_366;
wire n_709;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_984;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_964;
wire n_802;
wire n_982;
wire n_831;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_409;
wire n_345;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_427;
wire n_288;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_187),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_53),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_123),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_186),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_101),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_73),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_48),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_160),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_32),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_66),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_40),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_12),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_181),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_15),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_188),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_85),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_80),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_65),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_42),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_170),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_139),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_6),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_93),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_71),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_44),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_89),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_45),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_6),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_17),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_72),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_154),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_84),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_142),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_167),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_57),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_39),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_163),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_159),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_156),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_68),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_147),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_29),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_105),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_106),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_49),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_109),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_179),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_5),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_77),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_75),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_102),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_117),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_64),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_140),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_150),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_121),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_118),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_183),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_189),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_17),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_114),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_35),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_108),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_7),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_208),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_211),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_205),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_263),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_194),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_196),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_200),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_237),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_201),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_223),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g274 ( 
.A(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_202),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_203),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_197),
.Y(n_277)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_254),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_197),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_213),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g281 ( 
.A(n_257),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_207),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_195),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_214),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_204),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_225),
.Y(n_286)
);

INVxp33_ASAP7_75t_SL g287 ( 
.A(n_259),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_229),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_210),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_206),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_209),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_207),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_230),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_215),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_236),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_216),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_238),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_239),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_251),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_252),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_217),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_220),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_225),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_255),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_260),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_259),
.Y(n_306)
);

INVxp33_ASAP7_75t_SL g307 ( 
.A(n_227),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_261),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_233),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_233),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_241),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_223),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_223),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_312),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_262),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_273),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_285),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_268),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_273),
.Y(n_319)
);

NOR2x1_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_223),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_290),
.B(n_218),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_306),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_266),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_269),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_306),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_291),
.B(n_219),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_270),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_272),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_275),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_276),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_264),
.Y(n_334)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_282),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_280),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_284),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_288),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_294),
.B(n_221),
.Y(n_339)
);

NOR2x1_ASAP7_75t_L g340 ( 
.A(n_282),
.B(n_240),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_264),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_293),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_222),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_289),
.Y(n_344)
);

NOR2x1_ASAP7_75t_L g345 ( 
.A(n_295),
.B(n_240),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_297),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_298),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_301),
.B(n_224),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_299),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_300),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_274),
.B(n_278),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_281),
.B(n_231),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_292),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_304),
.B(n_232),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_265),
.A2(n_247),
.B1(n_226),
.B2(n_245),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_305),
.B(n_226),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_311),
.A2(n_212),
.B1(n_228),
.B2(n_244),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_289),
.B(n_240),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_302),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_302),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_307),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_307),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_311),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_271),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_287),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_287),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_277),
.B(n_240),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_317),
.Y(n_369)
);

BUFx6f_ASAP7_75t_SL g370 ( 
.A(n_368),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_317),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_353),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_324),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_353),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_335),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_330),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_334),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_341),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_344),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_234),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_315),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_330),
.Y(n_383)
);

NAND2xp33_ASAP7_75t_R g384 ( 
.A(n_368),
.B(n_0),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_361),
.B(n_277),
.Y(n_385)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_316),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_323),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_319),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_333),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_329),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_339),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_340),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_333),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_325),
.Y(n_394)
);

CKINVDCx6p67_ASAP7_75t_R g395 ( 
.A(n_364),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_325),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_326),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_343),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_326),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_316),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_348),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_316),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_368),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_361),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_360),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_316),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_332),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_318),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_360),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_332),
.Y(n_411)
);

NOR2x1p5_ASAP7_75t_L g412 ( 
.A(n_365),
.B(n_198),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_324),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_328),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_332),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_318),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_328),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_350),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_350),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_362),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_316),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_350),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_366),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_362),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_350),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_354),
.B(n_351),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_359),
.B(n_242),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_350),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_322),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_362),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_318),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_331),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_362),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_357),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_R g435 ( 
.A(n_363),
.B(n_367),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_322),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_357),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_368),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_365),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_331),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_331),
.Y(n_441)
);

NOR2x1p5_ASAP7_75t_L g442 ( 
.A(n_404),
.B(n_367),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_377),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_363),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_405),
.B(n_359),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_377),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_359),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_382),
.B(n_352),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_385),
.B(n_356),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_376),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_441),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g452 ( 
.A(n_381),
.B(n_431),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_410),
.B(n_438),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_388),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_373),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_409),
.B(n_416),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_409),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_441),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g459 ( 
.A(n_434),
.B(n_355),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_388),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_387),
.B(n_279),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_390),
.B(n_279),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_416),
.B(n_349),
.Y(n_463)
);

NAND3x1_ASAP7_75t_L g464 ( 
.A(n_437),
.B(n_340),
.C(n_356),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_428),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_428),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_391),
.A2(n_349),
.B1(n_248),
.B2(n_256),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_429),
.Y(n_468)
);

CKINVDCx8_ASAP7_75t_R g469 ( 
.A(n_369),
.Y(n_469)
);

NOR3xp33_ASAP7_75t_L g470 ( 
.A(n_413),
.B(n_336),
.C(n_327),
.Y(n_470)
);

BUFx4f_ASAP7_75t_L g471 ( 
.A(n_381),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_403),
.A2(n_349),
.B1(n_322),
.B2(n_337),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_428),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_383),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_398),
.B(n_335),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_428),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_429),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_417),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_401),
.B(n_335),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_436),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_412),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_414),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_436),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_389),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_393),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_381),
.B(n_335),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_420),
.B(n_286),
.Y(n_488)
);

AND2x2_ASAP7_75t_SL g489 ( 
.A(n_384),
.B(n_286),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_396),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_424),
.B(n_335),
.Y(n_491)
);

AND2x6_ASAP7_75t_L g492 ( 
.A(n_432),
.B(n_345),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_397),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_440),
.B(n_335),
.Y(n_494)
);

AND2x2_ASAP7_75t_SL g495 ( 
.A(n_384),
.B(n_303),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_399),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_402),
.Y(n_497)
);

INVx6_ASAP7_75t_L g498 ( 
.A(n_400),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_371),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_435),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_430),
.B(n_303),
.Y(n_501)
);

INVx4_ASAP7_75t_SL g502 ( 
.A(n_370),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_402),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_407),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_392),
.B(n_322),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_433),
.B(n_198),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_427),
.B(n_327),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_406),
.B(n_337),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_439),
.B(n_199),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_408),
.B(n_336),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_435),
.B(n_199),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_400),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_411),
.A2(n_337),
.B1(n_347),
.B2(n_346),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_372),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_374),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_400),
.Y(n_516)
);

OR2x6_ASAP7_75t_L g517 ( 
.A(n_395),
.B(n_338),
.Y(n_517)
);

OR2x6_ASAP7_75t_L g518 ( 
.A(n_370),
.B(n_338),
.Y(n_518)
);

AND2x6_ASAP7_75t_L g519 ( 
.A(n_407),
.B(n_345),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_378),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_379),
.B(n_342),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_421),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_380),
.B(n_207),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_457),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_521),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_447),
.B(n_448),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_455),
.Y(n_527)
);

AO22x2_ASAP7_75t_L g528 ( 
.A1(n_459),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_444),
.B(n_423),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_477),
.Y(n_530)
);

INVxp67_ASAP7_75t_SL g531 ( 
.A(n_451),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_477),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_480),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_423),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_480),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_456),
.B(n_342),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_457),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_460),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_460),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_507),
.A2(n_425),
.B1(n_422),
.B2(n_419),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_484),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_484),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_449),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_486),
.B(n_458),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_485),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_485),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_489),
.A2(n_235),
.B1(n_258),
.B2(n_246),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_490),
.Y(n_548)
);

AO22x2_ASAP7_75t_L g549 ( 
.A1(n_495),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_490),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_L g551 ( 
.A(n_452),
.B(n_492),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_496),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_456),
.B(n_346),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_496),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_478),
.B(n_347),
.Y(n_555)
);

AND2x6_ASAP7_75t_L g556 ( 
.A(n_453),
.B(n_421),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_457),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_445),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_509),
.B(n_418),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_449),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_482),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_450),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_474),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_493),
.B(n_235),
.Y(n_564)
);

NAND2x1p5_ASAP7_75t_L g565 ( 
.A(n_471),
.B(n_415),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_520),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_514),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_510),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_486),
.B(n_358),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_463),
.Y(n_570)
);

NOR2xp67_ASAP7_75t_L g571 ( 
.A(n_515),
.B(n_467),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_468),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_510),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_483),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_461),
.A2(n_258),
.B1(n_249),
.B2(n_253),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_462),
.B(n_243),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_508),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_499),
.B(n_321),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_503),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_503),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_463),
.Y(n_581)
);

OAI221xp5_ASAP7_75t_L g582 ( 
.A1(n_472),
.A2(n_314),
.B1(n_320),
.B2(n_5),
.C(n_7),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_458),
.B(n_314),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_443),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_535),
.Y(n_585)
);

A2O1A1Ixp33_ASAP7_75t_L g586 ( 
.A1(n_526),
.A2(n_507),
.B(n_488),
.C(n_501),
.Y(n_586)
);

NAND2x1_ASAP7_75t_L g587 ( 
.A(n_530),
.B(n_465),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_559),
.B(n_493),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_549),
.A2(n_493),
.B1(n_470),
.B2(n_452),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_577),
.A2(n_464),
.B(n_505),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_544),
.A2(n_476),
.B(n_465),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_529),
.B(n_525),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_525),
.B(n_469),
.Y(n_593)
);

O2A1O1Ixp5_ASAP7_75t_L g594 ( 
.A1(n_576),
.A2(n_479),
.B(n_487),
.C(n_491),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_532),
.Y(n_595)
);

A2O1A1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_558),
.A2(n_481),
.B(n_451),
.C(n_511),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_527),
.B(n_442),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_SL g598 ( 
.A(n_582),
.B(n_523),
.Y(n_598)
);

OAI21x1_ASAP7_75t_L g599 ( 
.A1(n_565),
.A2(n_569),
.B(n_579),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_541),
.B(n_475),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_567),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_542),
.B(n_506),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_544),
.A2(n_476),
.B(n_473),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_533),
.Y(n_604)
);

O2A1O1Ixp33_ASAP7_75t_L g605 ( 
.A1(n_558),
.A2(n_454),
.B(n_446),
.C(n_518),
.Y(n_605)
);

A2O1A1Ixp33_ASAP7_75t_L g606 ( 
.A1(n_545),
.A2(n_522),
.B(n_497),
.C(n_504),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_570),
.A2(n_452),
.B1(n_492),
.B2(n_494),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_551),
.A2(n_473),
.B(n_466),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_528),
.A2(n_518),
.B1(n_513),
.B2(n_517),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_583),
.A2(n_466),
.B(n_512),
.Y(n_610)
);

O2A1O1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_582),
.A2(n_497),
.B(n_504),
.C(n_516),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_549),
.A2(n_492),
.B1(n_519),
.B2(n_494),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_569),
.A2(n_531),
.B(n_540),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_546),
.B(n_519),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_570),
.A2(n_375),
.B(n_386),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_568),
.A2(n_375),
.B(n_386),
.Y(n_616)
);

AND2x4_ASAP7_75t_SL g617 ( 
.A(n_524),
.B(n_517),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_548),
.B(n_519),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_550),
.B(n_552),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g620 ( 
.A1(n_554),
.A2(n_519),
.B(n_320),
.Y(n_620)
);

O2A1O1Ixp5_ASAP7_75t_L g621 ( 
.A1(n_564),
.A2(n_498),
.B(n_502),
.C(n_386),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_573),
.A2(n_539),
.B(n_538),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_571),
.A2(n_498),
.B1(n_502),
.B2(n_386),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_524),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_580),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_572),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_536),
.A2(n_34),
.B(n_33),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_536),
.A2(n_37),
.B(n_36),
.Y(n_628)
);

BUFx4f_ASAP7_75t_L g629 ( 
.A(n_524),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_578),
.B(n_3),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_553),
.A2(n_41),
.B(n_38),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_574),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_562),
.Y(n_633)
);

AND2x2_ASAP7_75t_SL g634 ( 
.A(n_534),
.B(n_4),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_563),
.B(n_8),
.Y(n_635)
);

AO21x1_ASAP7_75t_L g636 ( 
.A1(n_565),
.A2(n_8),
.B(n_9),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_561),
.B(n_9),
.Y(n_637)
);

NOR2xp67_ASAP7_75t_L g638 ( 
.A(n_566),
.B(n_561),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_584),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_592),
.B(n_581),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_588),
.A2(n_553),
.B(n_537),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_613),
.A2(n_557),
.B(n_537),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_586),
.B(n_566),
.Y(n_643)
);

NAND2x1p5_ASAP7_75t_L g644 ( 
.A(n_629),
.B(n_537),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_593),
.B(n_555),
.Y(n_645)
);

A2O1A1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_598),
.A2(n_560),
.B(n_543),
.C(n_557),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_598),
.B(n_556),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_591),
.A2(n_557),
.B(n_560),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_SL g649 ( 
.A1(n_634),
.A2(n_547),
.B1(n_549),
.B2(n_528),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_633),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_602),
.B(n_575),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_603),
.A2(n_528),
.B(n_556),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_585),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_638),
.B(n_556),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_597),
.B(n_556),
.Y(n_655)
);

A2O1A1Ixp33_ASAP7_75t_L g656 ( 
.A1(n_590),
.A2(n_605),
.B(n_596),
.C(n_594),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_630),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_629),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_601),
.B(n_10),
.Y(n_659)
);

NOR2x1_ASAP7_75t_R g660 ( 
.A(n_624),
.B(n_43),
.Y(n_660)
);

OR2x6_ASAP7_75t_SL g661 ( 
.A(n_609),
.B(n_11),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_609),
.B(n_13),
.Y(n_662)
);

A2O1A1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_590),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_619),
.B(n_14),
.Y(n_664)
);

OA22x2_ASAP7_75t_L g665 ( 
.A1(n_617),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_600),
.B(n_16),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_595),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_624),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_624),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_632),
.B(n_193),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_626),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_604),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_625),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_639),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_635),
.B(n_18),
.Y(n_675)
);

O2A1O1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_637),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_618),
.B(n_20),
.Y(n_677)
);

AOI21x1_ASAP7_75t_L g678 ( 
.A1(n_610),
.A2(n_192),
.B(n_113),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_614),
.B(n_21),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_622),
.B(n_22),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_589),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_614),
.B(n_23),
.Y(n_682)
);

BUFx12f_ASAP7_75t_L g683 ( 
.A(n_636),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_606),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_623),
.B(n_612),
.Y(n_685)
);

NOR3xp33_ASAP7_75t_SL g686 ( 
.A(n_627),
.B(n_24),
.C(n_25),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_607),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_599),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_587),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_611),
.A2(n_119),
.B(n_191),
.Y(n_690)
);

BUFx4f_ASAP7_75t_L g691 ( 
.A(n_621),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_620),
.B(n_26),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_608),
.A2(n_116),
.B(n_190),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_628),
.Y(n_694)
);

INVxp67_ASAP7_75t_SL g695 ( 
.A(n_672),
.Y(n_695)
);

INVxp67_ASAP7_75t_SL g696 ( 
.A(n_640),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_669),
.Y(n_697)
);

CKINVDCx6p67_ASAP7_75t_R g698 ( 
.A(n_658),
.Y(n_698)
);

NAND2x1p5_ASAP7_75t_L g699 ( 
.A(n_658),
.B(n_631),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_669),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_674),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_649),
.A2(n_620),
.B1(n_616),
.B2(n_615),
.Y(n_702)
);

INVxp67_ASAP7_75t_SL g703 ( 
.A(n_671),
.Y(n_703)
);

NAND2x1p5_ASAP7_75t_L g704 ( 
.A(n_669),
.B(n_46),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_667),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_645),
.B(n_27),
.Y(n_706)
);

INVx6_ASAP7_75t_L g707 ( 
.A(n_671),
.Y(n_707)
);

INVx5_ASAP7_75t_L g708 ( 
.A(n_668),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_668),
.Y(n_709)
);

BUFx4f_ASAP7_75t_SL g710 ( 
.A(n_671),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_659),
.Y(n_711)
);

INVx8_ASAP7_75t_L g712 ( 
.A(n_670),
.Y(n_712)
);

NAND2x1p5_ASAP7_75t_L g713 ( 
.A(n_654),
.B(n_47),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_644),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_650),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_653),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_651),
.B(n_28),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_643),
.B(n_28),
.Y(n_718)
);

BUFx8_ASAP7_75t_L g719 ( 
.A(n_692),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_655),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_670),
.Y(n_721)
);

INVx8_ASAP7_75t_L g722 ( 
.A(n_683),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_689),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_673),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_646),
.B(n_29),
.Y(n_725)
);

NAND2x1p5_ASAP7_75t_L g726 ( 
.A(n_689),
.B(n_50),
.Y(n_726)
);

INVx5_ASAP7_75t_SL g727 ( 
.A(n_660),
.Y(n_727)
);

BUFx2_ASAP7_75t_SL g728 ( 
.A(n_665),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_661),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_686),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_691),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_666),
.B(n_30),
.Y(n_732)
);

BUFx6f_ASAP7_75t_SL g733 ( 
.A(n_694),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_691),
.Y(n_734)
);

BUFx6f_ASAP7_75t_SL g735 ( 
.A(n_684),
.Y(n_735)
);

CKINVDCx11_ASAP7_75t_R g736 ( 
.A(n_688),
.Y(n_736)
);

INVx2_ASAP7_75t_R g737 ( 
.A(n_656),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_647),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_682),
.Y(n_739)
);

BUFx8_ASAP7_75t_SL g740 ( 
.A(n_675),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_680),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_679),
.B(n_30),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_678),
.Y(n_743)
);

BUFx8_ASAP7_75t_L g744 ( 
.A(n_676),
.Y(n_744)
);

NAND2x1p5_ASAP7_75t_L g745 ( 
.A(n_641),
.B(n_51),
.Y(n_745)
);

NAND2x1p5_ASAP7_75t_L g746 ( 
.A(n_685),
.B(n_52),
.Y(n_746)
);

INVx6_ASAP7_75t_SL g747 ( 
.A(n_663),
.Y(n_747)
);

NAND2x1p5_ASAP7_75t_L g748 ( 
.A(n_662),
.B(n_54),
.Y(n_748)
);

INVx8_ASAP7_75t_L g749 ( 
.A(n_648),
.Y(n_749)
);

INVxp67_ASAP7_75t_SL g750 ( 
.A(n_642),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_664),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_677),
.B(n_31),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_652),
.Y(n_753)
);

NAND2x1p5_ASAP7_75t_L g754 ( 
.A(n_681),
.B(n_55),
.Y(n_754)
);

NAND2x1p5_ASAP7_75t_L g755 ( 
.A(n_687),
.B(n_56),
.Y(n_755)
);

NAND2x1p5_ASAP7_75t_L g756 ( 
.A(n_693),
.B(n_58),
.Y(n_756)
);

OR2x6_ASAP7_75t_L g757 ( 
.A(n_690),
.B(n_59),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_657),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_640),
.Y(n_759)
);

INVx5_ASAP7_75t_SL g760 ( 
.A(n_669),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_711),
.B(n_60),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_753),
.Y(n_762)
);

INVx5_ASAP7_75t_L g763 ( 
.A(n_731),
.Y(n_763)
);

AO32x2_ASAP7_75t_L g764 ( 
.A1(n_737),
.A2(n_31),
.A3(n_32),
.B1(n_61),
.B2(n_62),
.Y(n_764)
);

OA21x2_ASAP7_75t_L g765 ( 
.A1(n_743),
.A2(n_63),
.B(n_67),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_715),
.Y(n_766)
);

OA21x2_ASAP7_75t_L g767 ( 
.A1(n_743),
.A2(n_69),
.B(n_70),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_716),
.Y(n_768)
);

BUFx10_ASAP7_75t_L g769 ( 
.A(n_735),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_753),
.Y(n_770)
);

NAND2x1p5_ASAP7_75t_L g771 ( 
.A(n_708),
.B(n_74),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_716),
.Y(n_772)
);

NOR3xp33_ASAP7_75t_L g773 ( 
.A(n_717),
.B(n_76),
.C(n_78),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_742),
.B(n_79),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_705),
.Y(n_775)
);

OAI222xp33_ASAP7_75t_L g776 ( 
.A1(n_758),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.C1(n_86),
.C2(n_87),
.Y(n_776)
);

O2A1O1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_706),
.A2(n_88),
.B(n_90),
.C(n_91),
.Y(n_777)
);

OAI21x1_ASAP7_75t_L g778 ( 
.A1(n_750),
.A2(n_92),
.B(n_94),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_739),
.A2(n_95),
.B(n_96),
.C(n_97),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_699),
.A2(n_98),
.B(n_99),
.Y(n_780)
);

OAI21x1_ASAP7_75t_L g781 ( 
.A1(n_756),
.A2(n_702),
.B(n_745),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_725),
.A2(n_100),
.B(n_103),
.C(n_104),
.Y(n_782)
);

AOI221x1_ASAP7_75t_L g783 ( 
.A1(n_741),
.A2(n_107),
.B1(n_110),
.B2(n_111),
.C(n_112),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_707),
.Y(n_784)
);

OAI21x1_ASAP7_75t_L g785 ( 
.A1(n_741),
.A2(n_115),
.B(n_120),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_733),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_695),
.Y(n_787)
);

CKINVDCx11_ASAP7_75t_R g788 ( 
.A(n_736),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_696),
.B(n_759),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_721),
.B(n_703),
.Y(n_790)
);

OA21x2_ASAP7_75t_L g791 ( 
.A1(n_718),
.A2(n_122),
.B(n_124),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_721),
.B(n_125),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_720),
.B(n_126),
.Y(n_793)
);

OAI21x1_ASAP7_75t_L g794 ( 
.A1(n_746),
.A2(n_127),
.B(n_128),
.Y(n_794)
);

AO32x2_ASAP7_75t_L g795 ( 
.A1(n_697),
.A2(n_129),
.A3(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_730),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_796)
);

OAI21x1_ASAP7_75t_L g797 ( 
.A1(n_723),
.A2(n_136),
.B(n_137),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_724),
.Y(n_798)
);

OAI21x1_ASAP7_75t_SL g799 ( 
.A1(n_718),
.A2(n_138),
.B(n_141),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_738),
.Y(n_800)
);

NOR2xp67_ASAP7_75t_L g801 ( 
.A(n_751),
.B(n_143),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_707),
.Y(n_802)
);

INVx5_ASAP7_75t_L g803 ( 
.A(n_731),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_712),
.A2(n_144),
.B(n_145),
.C(n_146),
.Y(n_804)
);

OAI21x1_ASAP7_75t_L g805 ( 
.A1(n_723),
.A2(n_148),
.B(n_149),
.Y(n_805)
);

OAI21x1_ASAP7_75t_L g806 ( 
.A1(n_713),
.A2(n_151),
.B(n_152),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_726),
.A2(n_153),
.B(n_155),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_738),
.Y(n_808)
);

BUFx8_ASAP7_75t_L g809 ( 
.A(n_735),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_738),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_731),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_759),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_740),
.B(n_157),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_700),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_749),
.A2(n_158),
.B(n_161),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_733),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_728),
.B(n_162),
.Y(n_817)
);

OAI21x1_ASAP7_75t_L g818 ( 
.A1(n_704),
.A2(n_164),
.B(n_166),
.Y(n_818)
);

NAND2x1p5_ASAP7_75t_L g819 ( 
.A(n_708),
.B(n_168),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_762),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_762),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_766),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_787),
.B(n_732),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_770),
.B(n_752),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_770),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_812),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_814),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_769),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_769),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_768),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_772),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_789),
.Y(n_832)
);

BUFx12f_ASAP7_75t_L g833 ( 
.A(n_788),
.Y(n_833)
);

CKINVDCx6p67_ASAP7_75t_R g834 ( 
.A(n_763),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_775),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_800),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_786),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_809),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_786),
.Y(n_839)
);

NOR2xp67_ASAP7_75t_L g840 ( 
.A(n_816),
.B(n_734),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_765),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_810),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_809),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_798),
.Y(n_844)
);

OA21x2_ASAP7_75t_L g845 ( 
.A1(n_783),
.A2(n_701),
.B(n_747),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_764),
.Y(n_846)
);

BUFx2_ASAP7_75t_SL g847 ( 
.A(n_816),
.Y(n_847)
);

AO21x1_ASAP7_75t_SL g848 ( 
.A1(n_776),
.A2(n_744),
.B(n_747),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_773),
.A2(n_744),
.B1(n_754),
.B2(n_755),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_808),
.Y(n_850)
);

AO21x2_ASAP7_75t_L g851 ( 
.A1(n_781),
.A2(n_749),
.B(n_757),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_765),
.Y(n_852)
);

BUFx2_ASAP7_75t_L g853 ( 
.A(n_790),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_764),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_802),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_764),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_767),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_767),
.Y(n_858)
);

AOI21x1_ASAP7_75t_L g859 ( 
.A1(n_778),
.A2(n_757),
.B(n_734),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_791),
.Y(n_860)
);

INVx5_ASAP7_75t_L g861 ( 
.A(n_763),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_791),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_795),
.Y(n_863)
);

NAND2x1p5_ASAP7_75t_L g864 ( 
.A(n_763),
.B(n_734),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_795),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_795),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_785),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_837),
.Y(n_868)
);

INVxp33_ASAP7_75t_SL g869 ( 
.A(n_843),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_835),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_820),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_822),
.B(n_821),
.Y(n_872)
);

OAI22xp33_ASAP7_75t_L g873 ( 
.A1(n_845),
.A2(n_729),
.B1(n_817),
.B2(n_722),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_R g874 ( 
.A(n_843),
.B(n_811),
.Y(n_874)
);

NAND2xp33_ASAP7_75t_R g875 ( 
.A(n_853),
.B(n_813),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_821),
.B(n_811),
.Y(n_876)
);

AND2x2_ASAP7_75t_SL g877 ( 
.A(n_866),
.B(n_792),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_825),
.B(n_774),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_820),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_833),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_826),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_832),
.B(n_719),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_853),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_825),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_848),
.A2(n_719),
.B1(n_728),
.B2(n_799),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_836),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_830),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_824),
.B(n_793),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_849),
.A2(n_777),
.B(n_779),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_R g890 ( 
.A(n_838),
.B(n_710),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_824),
.B(n_701),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_835),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_828),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_844),
.B(n_722),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_R g895 ( 
.A(n_833),
.B(n_698),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_R g896 ( 
.A(n_834),
.B(n_803),
.Y(n_896)
);

INVx6_ASAP7_75t_L g897 ( 
.A(n_861),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_827),
.B(n_761),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_836),
.Y(n_899)
);

NOR2x1p5_ASAP7_75t_L g900 ( 
.A(n_880),
.B(n_828),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_881),
.B(n_860),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_879),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_879),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_886),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_883),
.B(n_837),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_868),
.B(n_839),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_886),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_883),
.B(n_839),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_886),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_899),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_884),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_899),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_884),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_868),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_870),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_875),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_876),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_872),
.B(n_846),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_870),
.B(n_860),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_887),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_872),
.B(n_892),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_887),
.Y(n_922)
);

AO21x2_ASAP7_75t_L g923 ( 
.A1(n_911),
.A2(n_862),
.B(n_858),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_902),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_916),
.A2(n_889),
.B1(n_873),
.B2(n_885),
.Y(n_925)
);

OAI21xp33_ASAP7_75t_L g926 ( 
.A1(n_901),
.A2(n_888),
.B(n_878),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_SL g927 ( 
.A1(n_905),
.A2(n_845),
.B1(n_863),
.B2(n_866),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_901),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_904),
.Y(n_929)
);

CKINVDCx6p67_ASAP7_75t_R g930 ( 
.A(n_906),
.Y(n_930)
);

AO21x2_ASAP7_75t_L g931 ( 
.A1(n_911),
.A2(n_862),
.B(n_841),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_914),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_904),
.Y(n_933)
);

NOR2x1_ASAP7_75t_SL g934 ( 
.A(n_905),
.B(n_847),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_902),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_917),
.B(n_877),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_909),
.B(n_893),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_921),
.B(n_878),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_907),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_930),
.B(n_908),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_924),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_924),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_925),
.B(n_921),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_SL g944 ( 
.A1(n_927),
.A2(n_815),
.B(n_869),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_930),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_936),
.A2(n_900),
.B1(n_863),
.B2(n_846),
.Y(n_946)
);

AO21x2_ASAP7_75t_L g947 ( 
.A1(n_934),
.A2(n_913),
.B(n_903),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_935),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_923),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_926),
.B(n_908),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_940),
.B(n_945),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_943),
.B(n_932),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_940),
.B(n_934),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_941),
.Y(n_954)
);

OR2x6_ASAP7_75t_L g955 ( 
.A(n_944),
.B(n_828),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_947),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_942),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_945),
.B(n_936),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_952),
.B(n_950),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_954),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_954),
.Y(n_961)
);

OR2x2_ASAP7_75t_L g962 ( 
.A(n_958),
.B(n_948),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_955),
.A2(n_951),
.B1(n_953),
.B2(n_946),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_957),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_955),
.B(n_938),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_960),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_963),
.A2(n_953),
.B1(n_880),
.B2(n_957),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_962),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_961),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_964),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_965),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_959),
.B(n_937),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_962),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_960),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_960),
.Y(n_975)
);

NAND3xp33_ASAP7_75t_L g976 ( 
.A(n_960),
.B(n_956),
.C(n_949),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_972),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_968),
.B(n_869),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_968),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_971),
.B(n_895),
.Y(n_980)
);

NAND2x1p5_ASAP7_75t_L g981 ( 
.A(n_973),
.B(n_828),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_966),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_969),
.Y(n_983)
);

NAND2x1_ASAP7_75t_SL g984 ( 
.A(n_970),
.B(n_928),
.Y(n_984)
);

OAI21xp33_ASAP7_75t_SL g985 ( 
.A1(n_984),
.A2(n_978),
.B(n_979),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_978),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_980),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_977),
.Y(n_988)
);

OAI22xp33_ASAP7_75t_L g989 ( 
.A1(n_981),
.A2(n_967),
.B1(n_976),
.B2(n_974),
.Y(n_989)
);

AOI322xp5_ASAP7_75t_L g990 ( 
.A1(n_982),
.A2(n_975),
.A3(n_949),
.B1(n_898),
.B2(n_976),
.C1(n_856),
.C2(n_854),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_983),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_985),
.B(n_981),
.Y(n_992)
);

NOR2x1_ASAP7_75t_L g993 ( 
.A(n_987),
.B(n_947),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_986),
.B(n_882),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_988),
.B(n_890),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_991),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_989),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_995),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_992),
.B(n_828),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_997),
.B(n_990),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_996),
.B(n_935),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_994),
.B(n_937),
.Y(n_1002)
);

AOI211xp5_ASAP7_75t_SL g1003 ( 
.A1(n_993),
.A2(n_796),
.B(n_804),
.C(n_801),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_998),
.Y(n_1004)
);

NOR3xp33_ASAP7_75t_L g1005 ( 
.A(n_999),
.B(n_894),
.C(n_782),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_1002),
.B(n_829),
.Y(n_1006)
);

NAND4xp25_ASAP7_75t_SL g1007 ( 
.A(n_1000),
.B(n_855),
.C(n_823),
.D(n_874),
.Y(n_1007)
);

NAND3xp33_ASAP7_75t_SL g1008 ( 
.A(n_1003),
.B(n_819),
.C(n_771),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_1001),
.B(n_929),
.Y(n_1009)
);

AOI21x1_ASAP7_75t_L g1010 ( 
.A1(n_1004),
.A2(n_937),
.B(n_840),
.Y(n_1010)
);

AOI222xp33_ASAP7_75t_L g1011 ( 
.A1(n_1008),
.A2(n_727),
.B1(n_829),
.B2(n_929),
.C1(n_939),
.C2(n_933),
.Y(n_1011)
);

OAI211xp5_ASAP7_75t_SL g1012 ( 
.A1(n_1006),
.A2(n_823),
.B(n_727),
.C(n_802),
.Y(n_1012)
);

OAI211xp5_ASAP7_75t_SL g1013 ( 
.A1(n_1009),
.A2(n_784),
.B(n_891),
.C(n_829),
.Y(n_1013)
);

AOI221xp5_ASAP7_75t_L g1014 ( 
.A1(n_1007),
.A2(n_829),
.B1(n_847),
.B2(n_896),
.C(n_893),
.Y(n_1014)
);

AOI221xp5_ASAP7_75t_L g1015 ( 
.A1(n_1005),
.A2(n_829),
.B1(n_939),
.B2(n_933),
.C(n_906),
.Y(n_1015)
);

AOI211xp5_ASAP7_75t_SL g1016 ( 
.A1(n_1004),
.A2(n_792),
.B(n_714),
.C(n_834),
.Y(n_1016)
);

OAI221xp5_ASAP7_75t_L g1017 ( 
.A1(n_1015),
.A2(n_864),
.B1(n_803),
.B2(n_897),
.C(n_748),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_1010),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_1014),
.Y(n_1019)
);

OAI322xp33_ASAP7_75t_L g1020 ( 
.A1(n_1011),
.A2(n_854),
.A3(n_919),
.B1(n_907),
.B2(n_865),
.C1(n_864),
.C2(n_909),
.Y(n_1020)
);

AOI211xp5_ASAP7_75t_L g1021 ( 
.A1(n_1012),
.A2(n_818),
.B(n_807),
.C(n_780),
.Y(n_1021)
);

NAND3xp33_ASAP7_75t_L g1022 ( 
.A(n_1016),
.B(n_1013),
.C(n_803),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_SL g1023 ( 
.A1(n_1012),
.A2(n_864),
.B1(n_709),
.B2(n_906),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1010),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_SL g1025 ( 
.A1(n_1012),
.A2(n_714),
.B(n_859),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1019),
.B(n_931),
.Y(n_1026)
);

NAND2x1p5_ASAP7_75t_L g1027 ( 
.A(n_1018),
.B(n_861),
.Y(n_1027)
);

NOR4xp25_ASAP7_75t_L g1028 ( 
.A(n_1024),
.B(n_920),
.C(n_922),
.D(n_903),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_1025),
.A2(n_845),
.B(n_931),
.C(n_923),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1022),
.Y(n_1030)
);

AOI211xp5_ASAP7_75t_L g1031 ( 
.A1(n_1017),
.A2(n_805),
.B(n_797),
.C(n_806),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1023),
.Y(n_1032)
);

AOI221xp5_ASAP7_75t_L g1033 ( 
.A1(n_1020),
.A2(n_913),
.B1(n_922),
.B2(n_920),
.C(n_909),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_SL g1034 ( 
.A1(n_1021),
.A2(n_859),
.B(n_842),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_1019),
.A2(n_897),
.B1(n_760),
.B2(n_923),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1032),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_1030),
.A2(n_931),
.B(n_794),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_1027),
.Y(n_1038)
);

NAND4xp75_ASAP7_75t_L g1039 ( 
.A(n_1026),
.B(n_845),
.C(n_760),
.D(n_877),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_1028),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_1035),
.B(n_897),
.Y(n_1041)
);

AOI222xp33_ASAP7_75t_L g1042 ( 
.A1(n_1034),
.A2(n_852),
.B1(n_858),
.B2(n_841),
.C1(n_867),
.C2(n_712),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1029),
.Y(n_1043)
);

NAND4xp25_ASAP7_75t_SL g1044 ( 
.A(n_1031),
.B(n_919),
.C(n_918),
.D(n_830),
.Y(n_1044)
);

NAND3xp33_ASAP7_75t_SL g1045 ( 
.A(n_1033),
.B(n_848),
.C(n_831),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_1032),
.B(n_861),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1032),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_SL g1048 ( 
.A(n_1027),
.B(n_831),
.C(n_867),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_1036),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_SL g1050 ( 
.A1(n_1047),
.A2(n_861),
.B1(n_708),
.B2(n_897),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_1040),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1038),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_R g1053 ( 
.A(n_1043),
.B(n_169),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_1046),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_1046),
.B(n_918),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_1041),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_1039),
.Y(n_1057)
);

INVxp67_ASAP7_75t_L g1058 ( 
.A(n_1051),
.Y(n_1058)
);

NAND3xp33_ASAP7_75t_L g1059 ( 
.A(n_1052),
.B(n_1042),
.C(n_1037),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1049),
.A2(n_1045),
.B1(n_1044),
.B2(n_1048),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_1054),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1057),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1057),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1056),
.A2(n_851),
.B(n_861),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_1060),
.A2(n_1055),
.B(n_1053),
.Y(n_1065)
);

INVx1_ASAP7_75t_SL g1066 ( 
.A(n_1061),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1058),
.Y(n_1067)
);

OAI31xp67_ASAP7_75t_L g1068 ( 
.A1(n_1062),
.A2(n_1050),
.A3(n_915),
.B(n_912),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1067),
.Y(n_1069)
);

OAI22x1_ASAP7_75t_SL g1070 ( 
.A1(n_1069),
.A2(n_1063),
.B1(n_1066),
.B2(n_1065),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1070),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1071),
.A2(n_1059),
.B1(n_1064),
.B2(n_1068),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_1071),
.A2(n_861),
.B1(n_912),
.B2(n_910),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1072),
.Y(n_1074)
);

OAI222xp33_ASAP7_75t_L g1075 ( 
.A1(n_1073),
.A2(n_915),
.B1(n_910),
.B2(n_852),
.C1(n_857),
.C2(n_871),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_1074),
.A2(n_851),
.B1(n_876),
.B2(n_850),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1075),
.A2(n_851),
.B1(n_857),
.B2(n_173),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1077),
.A2(n_171),
.B(n_172),
.Y(n_1078)
);

AOI211xp5_ASAP7_75t_L g1079 ( 
.A1(n_1078),
.A2(n_1076),
.B(n_177),
.C(n_178),
.Y(n_1079)
);

AOI211xp5_ASAP7_75t_L g1080 ( 
.A1(n_1079),
.A2(n_174),
.B(n_180),
.C(n_182),
.Y(n_1080)
);


endmodule