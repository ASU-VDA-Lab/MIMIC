module real_aes_6540_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_503;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_453;
wire n_374;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_519;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_500;
wire n_307;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g155 ( .A(n_0), .B(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g309 ( .A(n_1), .Y(n_309) );
AOI21xp33_ASAP7_75t_L g216 ( .A1(n_2), .A2(n_217), .B(n_218), .Y(n_216) );
INVx1_ASAP7_75t_L g174 ( .A(n_3), .Y(n_174) );
AND2x6_ASAP7_75t_L g191 ( .A(n_3), .B(n_172), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_3), .B(n_516), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_4), .A2(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g225 ( .A(n_5), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_6), .B(n_277), .Y(n_276) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_7), .A2(n_21), .B1(n_89), .B2(n_90), .Y(n_88) );
INVx1_ASAP7_75t_L g188 ( .A(n_8), .Y(n_188) );
INVx1_ASAP7_75t_L g291 ( .A(n_9), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_10), .A2(n_47), .B1(n_503), .B2(n_504), .Y(n_502) );
INVx1_ASAP7_75t_L g504 ( .A(n_10), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_11), .B(n_236), .Y(n_263) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_12), .A2(n_22), .B1(n_89), .B2(n_94), .Y(n_93) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_13), .B(n_217), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_14), .B(n_213), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_15), .A2(n_289), .B(n_290), .C(n_292), .Y(n_288) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_16), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_17), .B(n_223), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_18), .Y(n_116) );
INVx1_ASAP7_75t_L g201 ( .A(n_19), .Y(n_201) );
INVx2_ASAP7_75t_L g195 ( .A(n_20), .Y(n_195) );
OAI221xp5_ASAP7_75t_L g508 ( .A1(n_22), .A2(n_37), .B1(n_48), .B2(n_509), .C(n_510), .Y(n_508) );
INVxp67_ASAP7_75t_L g511 ( .A(n_22), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_23), .A2(n_191), .B(n_202), .C(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g199 ( .A(n_24), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_25), .B(n_223), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_26), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_27), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_28), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_29), .Y(n_131) );
CKINVDCx16_ASAP7_75t_R g205 ( .A(n_30), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_30), .A2(n_493), .B1(n_505), .B2(n_513), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_31), .B(n_217), .Y(n_279) );
OAI22xp5_ASAP7_75t_SL g499 ( .A1(n_32), .A2(n_55), .B1(n_259), .B2(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_32), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g83 ( .A1(n_33), .A2(n_56), .B1(n_84), .B2(n_99), .Y(n_83) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_34), .A2(n_193), .B1(n_196), .B2(n_202), .Y(n_192) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_34), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_35), .Y(n_256) );
CKINVDCx16_ASAP7_75t_R g306 ( .A(n_36), .Y(n_306) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_37), .A2(n_58), .B1(n_89), .B2(n_94), .Y(n_98) );
INVxp67_ASAP7_75t_L g512 ( .A(n_37), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_38), .A2(n_222), .B(n_224), .C(n_227), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_39), .Y(n_266) );
INVx1_ASAP7_75t_L g219 ( .A(n_40), .Y(n_219) );
INVx1_ASAP7_75t_L g172 ( .A(n_41), .Y(n_172) );
INVx1_ASAP7_75t_L g187 ( .A(n_42), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_43), .A2(n_70), .B1(n_160), .B2(n_164), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_44), .B(n_153), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_45), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_46), .A2(n_69), .B1(n_104), .B2(n_112), .Y(n_103) );
INVx1_ASAP7_75t_L g503 ( .A(n_47), .Y(n_503) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_48), .A2(n_64), .B1(n_89), .B2(n_90), .Y(n_96) );
AOI22xp33_ASAP7_75t_SL g141 ( .A1(n_49), .A2(n_54), .B1(n_142), .B2(n_147), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_SL g235 ( .A1(n_50), .A2(n_227), .B(n_236), .C(n_237), .Y(n_235) );
INVxp67_ASAP7_75t_L g238 ( .A(n_51), .Y(n_238) );
INVx1_ASAP7_75t_L g497 ( .A(n_52), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_53), .Y(n_210) );
INVx1_ASAP7_75t_L g259 ( .A(n_55), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_57), .A2(n_191), .B(n_202), .C(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_59), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g185 ( .A(n_60), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_61), .B(n_236), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g307 ( .A1(n_62), .A2(n_191), .B(n_202), .C(n_308), .Y(n_307) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_63), .B(n_80), .Y(n_79) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_65), .B(n_230), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_66), .Y(n_313) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_67), .A2(n_191), .B(n_202), .C(n_274), .Y(n_273) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_68), .Y(n_281) );
INVx1_ASAP7_75t_L g234 ( .A(n_71), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g287 ( .A(n_72), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_73), .B(n_249), .Y(n_275) );
INVx1_ASAP7_75t_L g89 ( .A(n_74), .Y(n_89) );
INVx1_ASAP7_75t_L g91 ( .A(n_74), .Y(n_91) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_75), .B(n_215), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_76), .A2(n_217), .B(n_233), .Y(n_232) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_167), .B1(n_175), .B2(n_487), .C(n_491), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
OAI322xp33_ASAP7_75t_L g491 ( .A1(n_80), .A2(n_492), .A3(n_517), .B1(n_518), .B2(n_519), .C1(n_522), .C2(n_523), .Y(n_491) );
AND2x2_ASAP7_75t_SL g80 ( .A(n_81), .B(n_135), .Y(n_80) );
INVxp67_ASAP7_75t_L g517 ( .A(n_81), .Y(n_517) );
NOR3xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_115), .C(n_126), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g82 ( .A(n_83), .B(n_103), .Y(n_82) );
BUFx3_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
AND2x4_ASAP7_75t_L g85 ( .A(n_86), .B(n_95), .Y(n_85) );
AND2x4_ASAP7_75t_L g100 ( .A(n_86), .B(n_101), .Y(n_100) );
AND2x2_ASAP7_75t_L g130 ( .A(n_86), .B(n_121), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_86), .B(n_109), .Y(n_134) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_92), .Y(n_86) );
AND2x2_ASAP7_75t_L g111 ( .A(n_87), .B(n_93), .Y(n_111) );
OR2x2_ASAP7_75t_L g120 ( .A(n_87), .B(n_93), .Y(n_120) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g139 ( .A(n_88), .B(n_93), .Y(n_139) );
AND2x2_ASAP7_75t_L g146 ( .A(n_88), .B(n_98), .Y(n_146) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g94 ( .A(n_91), .Y(n_94) );
AND2x2_ASAP7_75t_L g144 ( .A(n_92), .B(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g114 ( .A(n_93), .Y(n_114) );
AND2x6_ASAP7_75t_L g154 ( .A(n_95), .B(n_111), .Y(n_154) );
AND2x4_ASAP7_75t_L g158 ( .A(n_95), .B(n_119), .Y(n_158) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_97), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_96), .B(n_98), .Y(n_102) );
INVx1_ASAP7_75t_L g110 ( .A(n_96), .Y(n_110) );
INVx1_ASAP7_75t_L g122 ( .A(n_96), .Y(n_122) );
INVx1_ASAP7_75t_L g145 ( .A(n_96), .Y(n_145) );
AND2x2_ASAP7_75t_L g121 ( .A(n_97), .B(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_SL g99 ( .A(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OR2x6_ASAP7_75t_L g113 ( .A(n_102), .B(n_114), .Y(n_113) );
INVx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx4_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx8_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
INVx1_ASAP7_75t_L g166 ( .A(n_110), .Y(n_166) );
AND2x4_ASAP7_75t_L g125 ( .A(n_111), .B(n_121), .Y(n_125) );
INVx6_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g163 ( .A(n_114), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_117), .B1(n_123), .B2(n_124), .Y(n_115) );
INVx11_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x6_ASAP7_75t_L g138 ( .A(n_121), .B(n_139), .Y(n_138) );
INVx6_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B1(n_131), .B2(n_132), .Y(n_126) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVxp67_ASAP7_75t_L g518 ( .A(n_135), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_151), .Y(n_135) );
OAI21xp5_ASAP7_75t_SL g136 ( .A1(n_137), .A2(n_140), .B(n_141), .Y(n_136) );
INVx4_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g165 ( .A(n_139), .B(n_166), .Y(n_165) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
INVx1_ASAP7_75t_L g150 ( .A(n_145), .Y(n_150) );
AND2x4_ASAP7_75t_L g149 ( .A(n_146), .B(n_150), .Y(n_149) );
AND2x4_ASAP7_75t_L g162 ( .A(n_146), .B(n_163), .Y(n_162) );
BUFx4f_ASAP7_75t_SL g147 ( .A(n_148), .Y(n_147) );
BUFx12f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NAND3xp33_ASAP7_75t_L g151 ( .A(n_152), .B(n_155), .C(n_159), .Y(n_151) );
BUFx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx2_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_168), .Y(n_167) );
OR2x2_ASAP7_75t_SL g168 ( .A(n_169), .B(n_173), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND3x1_ASAP7_75t_SL g507 ( .A(n_170), .B(n_173), .C(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g513 ( .A(n_170), .B(n_514), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_170), .A2(n_202), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_171), .B(n_174), .Y(n_521) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND3x1_ASAP7_75t_L g176 ( .A(n_177), .B(n_412), .C(n_461), .Y(n_176) );
NOR3xp33_ASAP7_75t_SL g177 ( .A(n_178), .B(n_319), .C(n_357), .Y(n_177) );
OAI222xp33_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_240), .B1(n_294), .B2(n_300), .C1(n_314), .C2(n_317), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_180), .B(n_211), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_180), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_180), .B(n_362), .Y(n_453) );
BUFx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
OR2x2_ASAP7_75t_L g330 ( .A(n_181), .B(n_231), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_181), .B(n_212), .Y(n_338) );
AND2x2_ASAP7_75t_L g373 ( .A(n_181), .B(n_350), .Y(n_373) );
OR2x2_ASAP7_75t_L g397 ( .A(n_181), .B(n_212), .Y(n_397) );
OR2x2_ASAP7_75t_L g405 ( .A(n_181), .B(n_304), .Y(n_405) );
AND2x2_ASAP7_75t_L g408 ( .A(n_181), .B(n_231), .Y(n_408) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
OR2x2_ASAP7_75t_L g302 ( .A(n_182), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g316 ( .A(n_182), .B(n_231), .Y(n_316) );
AND2x2_ASAP7_75t_L g366 ( .A(n_182), .B(n_304), .Y(n_366) );
AND2x2_ASAP7_75t_L g379 ( .A(n_182), .B(n_212), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_182), .B(n_465), .Y(n_486) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_189), .B(n_209), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_183), .B(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g254 ( .A(n_183), .Y(n_254) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_183), .A2(n_305), .B(n_312), .Y(n_304) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_184), .Y(n_215) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
AND2x2_ASAP7_75t_SL g230 ( .A(n_185), .B(n_186), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_192), .B1(n_205), .B2(n_206), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_190), .A2(n_219), .B(n_220), .C(n_221), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_190), .A2(n_220), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g286 ( .A1(n_190), .A2(n_220), .B(n_287), .C(n_288), .Y(n_286) );
INVx4_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
NAND2x1p5_ASAP7_75t_L g206 ( .A(n_191), .B(n_207), .Y(n_206) );
AND2x4_ASAP7_75t_L g217 ( .A(n_191), .B(n_207), .Y(n_217) );
BUFx3_ASAP7_75t_L g490 ( .A(n_191), .Y(n_490) );
INVx2_ASAP7_75t_L g311 ( .A(n_193), .Y(n_311) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g203 ( .A(n_195), .Y(n_203) );
INVx1_ASAP7_75t_L g208 ( .A(n_195), .Y(n_208) );
OAI22xp5_ASAP7_75t_SL g196 ( .A1(n_197), .A2(n_199), .B1(n_200), .B2(n_201), .Y(n_196) );
INVx2_ASAP7_75t_L g200 ( .A(n_197), .Y(n_200) );
INVx4_ASAP7_75t_L g289 ( .A(n_197), .Y(n_289) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g204 ( .A(n_198), .Y(n_204) );
AND2x2_ASAP7_75t_L g207 ( .A(n_198), .B(n_208), .Y(n_207) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_198), .Y(n_223) );
INVx3_ASAP7_75t_L g226 ( .A(n_198), .Y(n_226) );
INVx1_ASAP7_75t_L g236 ( .A(n_198), .Y(n_236) );
INVx5_ASAP7_75t_L g220 ( .A(n_202), .Y(n_220) );
AND2x2_ASAP7_75t_L g489 ( .A(n_202), .B(n_490), .Y(n_489) );
AND2x6_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_203), .Y(n_228) );
BUFx3_ASAP7_75t_L g253 ( .A(n_203), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_205), .A2(n_507), .B1(n_524), .B2(n_525), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_206), .A2(n_259), .B(n_260), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_206), .A2(n_306), .B(n_307), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_L g404 ( .A1(n_211), .A2(n_405), .B(n_406), .C(n_409), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_211), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_211), .B(n_349), .Y(n_471) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_231), .Y(n_211) );
AND2x2_ASAP7_75t_SL g315 ( .A(n_212), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g329 ( .A(n_212), .Y(n_329) );
AND2x2_ASAP7_75t_L g356 ( .A(n_212), .B(n_350), .Y(n_356) );
INVx1_ASAP7_75t_SL g364 ( .A(n_212), .Y(n_364) );
AND2x2_ASAP7_75t_L g387 ( .A(n_212), .B(n_388), .Y(n_387) );
BUFx2_ASAP7_75t_L g465 ( .A(n_212), .Y(n_465) );
OA21x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_216), .B(n_229), .Y(n_212) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NOR2xp33_ASAP7_75t_SL g255 ( .A(n_214), .B(n_256), .Y(n_255) );
INVx4_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_215), .A2(n_232), .B(n_239), .Y(n_231) );
BUFx2_ASAP7_75t_L g285 ( .A(n_217), .Y(n_285) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx4_ASAP7_75t_L g277 ( .A(n_223), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_226), .B(n_238), .Y(n_237) );
INVx5_ASAP7_75t_L g249 ( .A(n_226), .Y(n_249) );
INVx3_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_228), .Y(n_278) );
INVx1_ASAP7_75t_L g267 ( .A(n_230), .Y(n_267) );
INVx2_ASAP7_75t_L g271 ( .A(n_230), .Y(n_271) );
OA21x2_ASAP7_75t_L g283 ( .A1(n_230), .A2(n_284), .B(n_293), .Y(n_283) );
BUFx2_ASAP7_75t_L g301 ( .A(n_231), .Y(n_301) );
INVx1_ASAP7_75t_L g363 ( .A(n_231), .Y(n_363) );
INVx3_ASAP7_75t_L g388 ( .A(n_231), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_240), .B(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_268), .Y(n_240) );
INVx1_ASAP7_75t_L g384 ( .A(n_241), .Y(n_384) );
OAI32xp33_ASAP7_75t_L g390 ( .A1(n_241), .A2(n_329), .A3(n_391), .B1(n_392), .B2(n_393), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_241), .A2(n_395), .B1(n_398), .B2(n_403), .Y(n_394) );
INVx4_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g332 ( .A(n_242), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g410 ( .A(n_242), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g480 ( .A(n_242), .B(n_426), .Y(n_480) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_257), .Y(n_242) );
AND2x2_ASAP7_75t_L g295 ( .A(n_243), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g325 ( .A(n_243), .Y(n_325) );
INVx1_ASAP7_75t_L g344 ( .A(n_243), .Y(n_344) );
OR2x2_ASAP7_75t_L g352 ( .A(n_243), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g359 ( .A(n_243), .B(n_333), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_243), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g380 ( .A(n_243), .B(n_298), .Y(n_380) );
INVx3_ASAP7_75t_L g402 ( .A(n_243), .Y(n_402) );
AND2x2_ASAP7_75t_L g427 ( .A(n_243), .B(n_299), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_243), .B(n_392), .Y(n_475) );
OR2x6_ASAP7_75t_L g243 ( .A(n_244), .B(n_255), .Y(n_243) );
AOI21xp5_ASAP7_75t_SL g244 ( .A1(n_245), .A2(n_246), .B(n_254), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_250), .B(n_251), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g308 ( .A1(n_249), .A2(n_309), .B(n_310), .C(n_311), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_251), .A2(n_262), .B(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g292 ( .A(n_253), .Y(n_292) );
INVx1_ASAP7_75t_L g264 ( .A(n_254), .Y(n_264) );
INVx2_ASAP7_75t_L g299 ( .A(n_257), .Y(n_299) );
AND2x2_ASAP7_75t_L g431 ( .A(n_257), .B(n_269), .Y(n_431) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_264), .B(n_265), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_267), .B(n_281), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_267), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g473 ( .A(n_268), .Y(n_473) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_282), .Y(n_268) );
INVx1_ASAP7_75t_L g318 ( .A(n_269), .Y(n_318) );
AND2x2_ASAP7_75t_L g345 ( .A(n_269), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_269), .B(n_299), .Y(n_353) );
AND2x2_ASAP7_75t_L g411 ( .A(n_269), .B(n_334), .Y(n_411) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g297 ( .A(n_270), .Y(n_297) );
AND2x2_ASAP7_75t_L g324 ( .A(n_270), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g333 ( .A(n_270), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_270), .B(n_299), .Y(n_399) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B(n_280), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_279), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B(n_278), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_282), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g346 ( .A(n_282), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_282), .B(n_299), .Y(n_392) );
AND2x2_ASAP7_75t_L g401 ( .A(n_282), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g426 ( .A(n_282), .Y(n_426) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g298 ( .A(n_283), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g334 ( .A(n_283), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_289), .B(n_291), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_294), .A2(n_304), .B1(n_463), .B2(n_466), .Y(n_462) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
OAI21xp5_ASAP7_75t_SL g485 ( .A1(n_296), .A2(n_407), .B(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_297), .B(n_402), .Y(n_419) );
INVx1_ASAP7_75t_L g444 ( .A(n_297), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_298), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g371 ( .A(n_298), .B(n_324), .Y(n_371) );
INVx2_ASAP7_75t_L g327 ( .A(n_299), .Y(n_327) );
INVx1_ASAP7_75t_L g377 ( .A(n_299), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g468 ( .A1(n_300), .A2(n_452), .B1(n_469), .B2(n_472), .C(n_474), .Y(n_468) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g339 ( .A(n_301), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_301), .B(n_350), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_302), .B(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g393 ( .A(n_302), .B(n_339), .Y(n_393) );
INVx3_ASAP7_75t_SL g434 ( .A(n_302), .Y(n_434) );
AND2x2_ASAP7_75t_L g378 ( .A(n_303), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g407 ( .A(n_303), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_303), .B(n_316), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_303), .B(n_362), .Y(n_448) );
INVx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx3_ASAP7_75t_L g350 ( .A(n_304), .Y(n_350) );
OAI322xp33_ASAP7_75t_L g445 ( .A1(n_304), .A2(n_376), .A3(n_398), .B1(n_446), .B2(n_448), .C1(n_449), .C2(n_450), .Y(n_445) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI21xp33_ASAP7_75t_L g469 ( .A1(n_315), .A2(n_318), .B(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_SL g395 ( .A(n_316), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g417 ( .A(n_316), .B(n_329), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_316), .B(n_356), .Y(n_432) );
INVxp67_ASAP7_75t_L g383 ( .A(n_318), .Y(n_383) );
AOI211xp5_ASAP7_75t_L g389 ( .A1(n_318), .A2(n_390), .B(n_394), .C(n_404), .Y(n_389) );
OAI221xp5_ASAP7_75t_SL g319 ( .A1(n_320), .A2(n_328), .B1(n_331), .B2(n_335), .C(n_340), .Y(n_319) );
INVxp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_326), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g343 ( .A(n_327), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g460 ( .A(n_327), .Y(n_460) );
OAI221xp5_ASAP7_75t_L g476 ( .A1(n_328), .A2(n_477), .B1(n_482), .B2(n_483), .C(n_485), .Y(n_476) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_329), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g376 ( .A(n_329), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_329), .B(n_407), .Y(n_414) );
AND2x2_ASAP7_75t_L g456 ( .A(n_329), .B(n_434), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_330), .B(n_355), .Y(n_354) );
OAI22xp33_ASAP7_75t_L g451 ( .A1(n_330), .A2(n_342), .B1(n_452), .B2(n_453), .Y(n_451) );
OR2x2_ASAP7_75t_L g482 ( .A(n_330), .B(n_350), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g459 ( .A(n_333), .Y(n_459) );
AND2x2_ASAP7_75t_L g484 ( .A(n_333), .B(n_427), .Y(n_484) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_SL g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g348 ( .A(n_338), .B(n_349), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_347), .B1(n_351), .B2(n_354), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
INVx1_ASAP7_75t_L g415 ( .A(n_343), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_343), .B(n_383), .Y(n_450) );
AOI322xp5_ASAP7_75t_L g374 ( .A1(n_345), .A2(n_375), .A3(n_377), .B1(n_378), .B2(n_380), .C1(n_381), .C2(n_385), .Y(n_374) );
INVxp67_ASAP7_75t_L g368 ( .A(n_346), .Y(n_368) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_348), .A2(n_353), .B1(n_370), .B2(n_372), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_349), .B(n_362), .Y(n_449) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_350), .B(n_388), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_350), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g446 ( .A(n_352), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
NAND3xp33_ASAP7_75t_SL g357 ( .A(n_358), .B(n_374), .C(n_389), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B1(n_365), .B2(n_367), .C(n_369), .Y(n_358) );
AND2x2_ASAP7_75t_L g365 ( .A(n_361), .B(n_366), .Y(n_365) );
INVx3_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
AND2x2_ASAP7_75t_L g375 ( .A(n_366), .B(n_376), .Y(n_375) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_368), .Y(n_447) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_373), .B(n_387), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_376), .B(n_434), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_377), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g452 ( .A(n_380), .Y(n_452) );
AND2x2_ASAP7_75t_L g467 ( .A(n_380), .B(n_444), .Y(n_467) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI211xp5_ASAP7_75t_L g461 ( .A1(n_391), .A2(n_462), .B(n_468), .C(n_476), .Y(n_461) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g430 ( .A(n_401), .B(n_431), .Y(n_430) );
NAND2x1_ASAP7_75t_SL g472 ( .A(n_402), .B(n_473), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g442 ( .A(n_405), .Y(n_442) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g437 ( .A(n_411), .Y(n_437) );
AND2x2_ASAP7_75t_L g441 ( .A(n_411), .B(n_427), .Y(n_441) );
NOR5xp2_ASAP7_75t_L g412 ( .A(n_413), .B(n_428), .C(n_445), .D(n_451), .E(n_454), .Y(n_412) );
OAI221xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B1(n_416), .B2(n_418), .C(n_420), .Y(n_413) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_417), .B(n_475), .Y(n_474) );
INVxp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g443 ( .A(n_427), .B(n_444), .Y(n_443) );
OAI221xp5_ASAP7_75t_SL g428 ( .A1(n_429), .A2(n_432), .B1(n_433), .B2(n_435), .C(n_438), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_441), .B1(n_442), .B2(n_443), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g481 ( .A(n_441), .Y(n_481) );
AOI211xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_457), .B(n_459), .C(n_460), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVxp67_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_481), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
CKINVDCx14_ASAP7_75t_R g483 ( .A(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_489), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_493), .Y(n_524) );
OAI22xp5_ASAP7_75t_SL g493 ( .A1(n_494), .A2(n_495), .B1(n_501), .B2(n_502), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B1(n_498), .B2(n_499), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
CKINVDCx14_ASAP7_75t_R g501 ( .A(n_502), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
INVxp67_ASAP7_75t_L g516 ( .A(n_508), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_513), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_515), .Y(n_514) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
CKINVDCx16_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
endmodule