module fake_jpeg_3770_n_96 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_96);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_5),
.B(n_11),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_23),
.B(n_17),
.Y(n_34)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_27),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_25),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_26),
.B(n_29),
.Y(n_40)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_20),
.B(n_0),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_21),
.B1(n_18),
.B2(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_19),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_33),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_53),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_46),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_21),
.B1(n_14),
.B2(n_22),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_50),
.C(n_38),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_22),
.B1(n_12),
.B2(n_14),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_43),
.Y(n_54)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_27),
.A2(n_12),
.B1(n_5),
.B2(n_7),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_49),
.B(n_52),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_30),
.A2(n_6),
.B(n_10),
.Y(n_50)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_29),
.B(n_10),
.Y(n_53)
);

AND2x6_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_35),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_48),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_11),
.Y(n_60)
);

AO22x1_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_50),
.B1(n_36),
.B2(n_40),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_53),
.B1(n_44),
.B2(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_34),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_76),
.B(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_73),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_40),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_70),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_43),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_39),
.B1(n_45),
.B2(n_42),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_54),
.B1(n_58),
.B2(n_65),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_77),
.C(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_47),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_75),
.B1(n_55),
.B2(n_64),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_52),
.C(n_45),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_61),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_84),
.B1(n_73),
.B2(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_81),
.B(n_67),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_54),
.C(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

AOI322xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_88),
.A3(n_78),
.B1(n_82),
.B2(n_84),
.C1(n_60),
.C2(n_59),
.Y(n_91)
);

OAI322xp33_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_56),
.A3(n_59),
.B1(n_60),
.B2(n_62),
.C1(n_82),
.C2(n_85),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_92),
.Y(n_94)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

AOI221xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_88),
.B1(n_90),
.B2(n_89),
.C(n_87),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_93),
.C(n_62),
.Y(n_96)
);


endmodule