module fake_netlist_5_1109_n_1469 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_451, n_408, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_452, n_397, n_111, n_155, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_470, n_325, n_449, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_457, n_297, n_156, n_5, n_225, n_377, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_430, n_313, n_88, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_213, n_129, n_342, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_461, n_333, n_309, n_30, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_85, n_463, n_239, n_466, n_420, n_55, n_49, n_310, n_54, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_441, n_450, n_312, n_429, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_425, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_409, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_391, n_434, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_52, n_278, n_110, n_1469);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_451;
input n_408;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_461;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_85;
input n_463;
input n_239;
input n_466;
input n_420;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_441;
input n_450;
input n_312;
input n_429;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_425;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_409;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_391;
input n_434;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1469;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_1314;
wire n_709;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_976;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_777;
wire n_1070;
wire n_1030;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1459;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_1072;
wire n_832;
wire n_857;
wire n_1319;
wire n_561;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_887;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_868;
wire n_639;
wire n_914;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_759;
wire n_806;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1233;
wire n_526;
wire n_677;
wire n_1333;
wire n_1121;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_514;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_1383;
wire n_1073;
wire n_662;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_860;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_950;
wire n_1346;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_912;
wire n_968;
wire n_619;
wire n_1386;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_753;
wire n_621;
wire n_1048;
wire n_1288;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1149;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1419;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_487;
wire n_665;
wire n_1440;
wire n_1356;
wire n_910;
wire n_768;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_754;
wire n_1125;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_827;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_1086;
wire n_796;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_852;
wire n_1028;
wire n_781;
wire n_542;
wire n_595;
wire n_502;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_480;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_107),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_89),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_377),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_384),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_161),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_417),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_475),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_284),
.Y(n_483)
);

BUFx10_ASAP7_75t_L g484 ( 
.A(n_315),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_162),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_180),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_243),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_233),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_120),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_63),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_331),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_435),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_19),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_338),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_441),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_180),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_264),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_75),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_202),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_425),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_97),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_452),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_198),
.Y(n_503)
);

CKINVDCx14_ASAP7_75t_R g504 ( 
.A(n_56),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_262),
.Y(n_505)
);

BUFx10_ASAP7_75t_L g506 ( 
.A(n_235),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_409),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_465),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_71),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_350),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_422),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_449),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_442),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_138),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_142),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_406),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_49),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_225),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_366),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_32),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_423),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_2),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_267),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_22),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_459),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_404),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_179),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_201),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_340),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_99),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_75),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g532 ( 
.A(n_339),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_356),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_49),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_419),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_372),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_168),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_394),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_140),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_139),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g541 ( 
.A(n_244),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_411),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_463),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_114),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_217),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_396),
.Y(n_546)
);

INVxp33_ASAP7_75t_L g547 ( 
.A(n_309),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_200),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_86),
.Y(n_549)
);

BUFx10_ASAP7_75t_L g550 ( 
.A(n_47),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_205),
.Y(n_551)
);

BUFx5_ASAP7_75t_L g552 ( 
.A(n_351),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_236),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_450),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_307),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_177),
.Y(n_556)
);

BUFx10_ASAP7_75t_L g557 ( 
.A(n_304),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_457),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_324),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_414),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_187),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_405),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_272),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_443),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_462),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_432),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_154),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_344),
.Y(n_568)
);

CKINVDCx14_ASAP7_75t_R g569 ( 
.A(n_448),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_393),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_415),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_21),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_95),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_383),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_116),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_316),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_440),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_385),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_71),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_380),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_226),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_326),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_418),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_388),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_431),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_436),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_323),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_90),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_455),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_337),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_81),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_277),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_122),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_386),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_230),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_251),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_314),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_445),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_281),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_454),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_421),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_399),
.Y(n_602)
);

BUFx10_ASAP7_75t_L g603 ( 
.A(n_6),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_348),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_363),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_120),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_460),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_461),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_473),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_292),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_146),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_329),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_174),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_429),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_458),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_392),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_117),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_430),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_319),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_364),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_426),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_40),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_470),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_73),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_424),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_398),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_44),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_387),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_446),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_456),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_301),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_32),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_401),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_137),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_444),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_165),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_223),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_413),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_60),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_78),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_295),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_193),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_89),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_174),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_325),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_433),
.Y(n_646)
);

BUFx5_ASAP7_75t_L g647 ( 
.A(n_453),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_403),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_306),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_332),
.Y(n_650)
);

CKINVDCx16_ASAP7_75t_R g651 ( 
.A(n_395),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_108),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_273),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_151),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_214),
.Y(n_655)
);

CKINVDCx14_ASAP7_75t_R g656 ( 
.A(n_142),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_439),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_322),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_8),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_250),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_467),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_416),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_428),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_7),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_94),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_447),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_402),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_400),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_119),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_171),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_96),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_135),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_451),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_434),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_438),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_165),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_158),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_162),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_437),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_73),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_420),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_464),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_407),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_410),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_173),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_276),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_69),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_232),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_397),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_128),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_85),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_408),
.Y(n_692)
);

CKINVDCx16_ASAP7_75t_R g693 ( 
.A(n_82),
.Y(n_693)
);

BUFx5_ASAP7_75t_L g694 ( 
.A(n_412),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_427),
.Y(n_695)
);

CKINVDCx16_ASAP7_75t_R g696 ( 
.A(n_693),
.Y(n_696)
);

INVxp33_ASAP7_75t_L g697 ( 
.A(n_622),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_486),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_678),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_486),
.Y(n_700)
);

INVxp33_ASAP7_75t_SL g701 ( 
.A(n_476),
.Y(n_701)
);

INVxp67_ASAP7_75t_SL g702 ( 
.A(n_596),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_482),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_535),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_639),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_489),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_506),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_490),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_599),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_483),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_547),
.B(n_0),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_498),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_610),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_503),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_491),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_509),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_477),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_504),
.B(n_0),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_492),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_698),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_700),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_706),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_708),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_712),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_714),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_717),
.B(n_569),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_716),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_705),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_718),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_699),
.B(n_493),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_711),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_711),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_696),
.A2(n_656),
.B1(n_532),
.B2(n_651),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_707),
.Y(n_734)
);

BUFx2_ASAP7_75t_L g735 ( 
.A(n_703),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_702),
.B(n_710),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_715),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_719),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_701),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_697),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_704),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_709),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_713),
.Y(n_743)
);

INVx4_ASAP7_75t_L g744 ( 
.A(n_729),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_728),
.Y(n_745)
);

OR2x6_ASAP7_75t_L g746 ( 
.A(n_741),
.B(n_516),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_722),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_731),
.B(n_629),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_724),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_735),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_740),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_728),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_729),
.Y(n_753)
);

AND2x6_ASAP7_75t_L g754 ( 
.A(n_733),
.B(n_528),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_723),
.Y(n_755)
);

NOR2x1p5_ASAP7_75t_L g756 ( 
.A(n_739),
.B(n_480),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_726),
.B(n_506),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_725),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_732),
.B(n_680),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_723),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_737),
.B(n_570),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_721),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_727),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_720),
.Y(n_764)
);

AND2x6_ASAP7_75t_L g765 ( 
.A(n_736),
.B(n_478),
.Y(n_765)
);

INVx4_ASAP7_75t_L g766 ( 
.A(n_738),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_734),
.B(n_601),
.Y(n_767)
);

OR2x2_ASAP7_75t_SL g768 ( 
.A(n_743),
.B(n_541),
.Y(n_768)
);

AND2x6_ASAP7_75t_L g769 ( 
.A(n_742),
.B(n_564),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_730),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_723),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_722),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_728),
.Y(n_773)
);

BUFx6f_ASAP7_75t_SL g774 ( 
.A(n_740),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_722),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_730),
.Y(n_776)
);

AND2x2_ASAP7_75t_SL g777 ( 
.A(n_730),
.B(n_539),
.Y(n_777)
);

NAND2x1p5_ASAP7_75t_L g778 ( 
.A(n_744),
.B(n_571),
.Y(n_778)
);

AO22x2_ASAP7_75t_L g779 ( 
.A1(n_776),
.A2(n_642),
.B1(n_537),
.B2(n_545),
.Y(n_779)
);

NAND2x1p5_ASAP7_75t_L g780 ( 
.A(n_753),
.B(n_597),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_747),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_749),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_758),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_777),
.B(n_757),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_772),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_761),
.B(n_626),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_767),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_748),
.A2(n_481),
.B(n_487),
.C(n_479),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_755),
.Y(n_789)
);

AO22x2_ASAP7_75t_L g790 ( 
.A1(n_759),
.A2(n_595),
.B1(n_522),
.B2(n_581),
.Y(n_790)
);

OA22x2_ASAP7_75t_L g791 ( 
.A1(n_751),
.A2(n_488),
.B1(n_499),
.B2(n_496),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_774),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_775),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_764),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_771),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_771),
.Y(n_796)
);

AO22x2_ASAP7_75t_L g797 ( 
.A1(n_754),
.A2(n_573),
.B1(n_644),
.B2(n_593),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_760),
.Y(n_798)
);

AO22x2_ASAP7_75t_L g799 ( 
.A1(n_754),
.A2(n_677),
.B1(n_685),
.B2(n_669),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_756),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_762),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_763),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_745),
.B(n_550),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_763),
.Y(n_804)
);

AO22x2_ASAP7_75t_L g805 ( 
.A1(n_768),
.A2(n_690),
.B1(n_574),
.B2(n_538),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_752),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_765),
.A2(n_695),
.B1(n_650),
.B2(n_645),
.Y(n_807)
);

OR2x2_ASAP7_75t_SL g808 ( 
.A(n_746),
.B(n_485),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_773),
.Y(n_809)
);

OAI221xp5_ASAP7_75t_L g810 ( 
.A1(n_766),
.A2(n_667),
.B1(n_641),
.B2(n_623),
.C(n_683),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_765),
.A2(n_692),
.B1(n_505),
.B2(n_508),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_769),
.B(n_501),
.Y(n_812)
);

AO22x2_ASAP7_75t_L g813 ( 
.A1(n_769),
.A2(n_495),
.B1(n_500),
.B2(n_494),
.Y(n_813)
);

NAND2xp33_ASAP7_75t_L g814 ( 
.A(n_765),
.B(n_497),
.Y(n_814)
);

OAI221xp5_ASAP7_75t_L g815 ( 
.A1(n_761),
.A2(n_604),
.B1(n_619),
.B2(n_594),
.C(n_586),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_747),
.Y(n_816)
);

BUFx8_ASAP7_75t_L g817 ( 
.A(n_774),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_747),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_747),
.Y(n_819)
);

OA22x2_ASAP7_75t_L g820 ( 
.A1(n_770),
.A2(n_515),
.B1(n_517),
.B2(n_514),
.Y(n_820)
);

AO22x2_ASAP7_75t_L g821 ( 
.A1(n_770),
.A2(n_511),
.B1(n_526),
.B2(n_512),
.Y(n_821)
);

OAI221xp5_ASAP7_75t_L g822 ( 
.A1(n_761),
.A2(n_625),
.B1(n_635),
.B2(n_616),
.C(n_608),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_747),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_747),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_750),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_753),
.B(n_580),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_748),
.B(n_587),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_747),
.Y(n_828)
);

OAI221xp5_ASAP7_75t_L g829 ( 
.A1(n_761),
.A2(n_673),
.B1(n_663),
.B2(n_605),
.C(n_609),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_759),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_777),
.A2(n_513),
.B1(n_519),
.B2(n_510),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_777),
.A2(n_523),
.B1(n_525),
.B2(n_521),
.Y(n_832)
);

AO22x2_ASAP7_75t_L g833 ( 
.A1(n_770),
.A2(n_600),
.B1(n_618),
.B2(n_602),
.Y(n_833)
);

OA22x2_ASAP7_75t_L g834 ( 
.A1(n_770),
.A2(n_518),
.B1(n_524),
.B2(n_520),
.Y(n_834)
);

AO22x2_ASAP7_75t_L g835 ( 
.A1(n_770),
.A2(n_620),
.B1(n_631),
.B2(n_628),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_770),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_748),
.B(n_646),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_777),
.A2(n_536),
.B1(n_542),
.B2(n_533),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_748),
.B(n_649),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_770),
.B(n_527),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_750),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_750),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_770),
.B(n_530),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_777),
.A2(n_546),
.B1(n_553),
.B2(n_543),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_755),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_770),
.B(n_550),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_747),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_787),
.B(n_554),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_836),
.B(n_555),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_786),
.B(n_657),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_830),
.B(n_559),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_807),
.B(n_560),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_781),
.B(n_562),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_782),
.B(n_668),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_802),
.B(n_674),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_840),
.B(n_843),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_783),
.B(n_563),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_785),
.B(n_565),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_793),
.B(n_566),
.Y(n_859)
);

NAND2xp33_ASAP7_75t_SL g860 ( 
.A(n_800),
.B(n_611),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_794),
.B(n_568),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_816),
.B(n_675),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_818),
.B(n_502),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_819),
.B(n_576),
.Y(n_864)
);

NAND2xp33_ASAP7_75t_SL g865 ( 
.A(n_812),
.B(n_632),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_823),
.B(n_577),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_824),
.B(n_578),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_828),
.B(n_558),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_847),
.B(n_582),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_811),
.B(n_584),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_831),
.B(n_585),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_832),
.B(n_589),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_838),
.B(n_590),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_844),
.B(n_592),
.Y(n_874)
);

NAND2xp33_ASAP7_75t_SL g875 ( 
.A(n_841),
.B(n_665),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_846),
.B(n_607),
.Y(n_876)
);

NAND2xp33_ASAP7_75t_SL g877 ( 
.A(n_789),
.B(n_691),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_827),
.B(n_612),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_837),
.B(n_614),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_839),
.B(n_615),
.Y(n_880)
);

NAND2xp33_ASAP7_75t_SL g881 ( 
.A(n_801),
.B(n_621),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_803),
.B(n_603),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_804),
.B(n_798),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_795),
.B(n_603),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_826),
.B(n_630),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_796),
.B(n_633),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_825),
.B(n_531),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_845),
.B(n_638),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_791),
.B(n_648),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_806),
.B(n_809),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_797),
.B(n_653),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_778),
.B(n_658),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_842),
.B(n_660),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_SL g894 ( 
.A(n_813),
.B(n_661),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_820),
.B(n_666),
.Y(n_895)
);

NAND2xp33_ASAP7_75t_SL g896 ( 
.A(n_814),
.B(n_681),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_808),
.B(n_687),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_834),
.B(n_682),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_792),
.B(n_780),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_788),
.B(n_684),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_799),
.B(n_686),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_817),
.B(n_689),
.Y(n_902)
);

NAND2xp33_ASAP7_75t_SL g903 ( 
.A(n_805),
.B(n_534),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_810),
.B(n_484),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_815),
.B(n_484),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_822),
.B(n_557),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_835),
.B(n_552),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_829),
.B(n_557),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_821),
.B(n_583),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_833),
.B(n_552),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_790),
.B(n_529),
.Y(n_911)
);

NAND2xp33_ASAP7_75t_SL g912 ( 
.A(n_779),
.B(n_540),
.Y(n_912)
);

NAND2xp33_ASAP7_75t_SL g913 ( 
.A(n_784),
.B(n_544),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_SL g914 ( 
.A(n_784),
.B(n_548),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_SL g915 ( 
.A(n_784),
.B(n_549),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_784),
.B(n_507),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_784),
.B(n_507),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_784),
.B(n_598),
.Y(n_918)
);

NAND2xp33_ASAP7_75t_SL g919 ( 
.A(n_784),
.B(n_551),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_784),
.B(n_598),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_784),
.B(n_662),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_784),
.B(n_662),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_784),
.B(n_679),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_787),
.B(n_556),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_784),
.B(n_679),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_784),
.B(n_552),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_784),
.B(n_552),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_784),
.B(n_647),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_787),
.B(n_561),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_784),
.B(n_647),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_802),
.B(n_237),
.Y(n_931)
);

NAND2xp33_ASAP7_75t_SL g932 ( 
.A(n_784),
.B(n_567),
.Y(n_932)
);

NAND2xp33_ASAP7_75t_SL g933 ( 
.A(n_784),
.B(n_572),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_784),
.B(n_647),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_786),
.B(n_647),
.Y(n_935)
);

NAND2xp33_ASAP7_75t_SL g936 ( 
.A(n_784),
.B(n_575),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_784),
.B(n_694),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_784),
.B(n_694),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_786),
.B(n_694),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_786),
.B(n_694),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_784),
.B(n_579),
.Y(n_941)
);

NAND2xp33_ASAP7_75t_SL g942 ( 
.A(n_784),
.B(n_588),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_786),
.B(n_591),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_784),
.B(n_606),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_784),
.B(n_613),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_802),
.B(n_238),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_786),
.B(n_617),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_786),
.B(n_624),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_784),
.B(n_627),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_784),
.B(n_634),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_784),
.B(n_636),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_787),
.B(n_637),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_786),
.B(n_640),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_784),
.B(n_643),
.Y(n_954)
);

NAND2xp33_ASAP7_75t_SL g955 ( 
.A(n_784),
.B(n_652),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_784),
.B(n_654),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_784),
.B(n_655),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_784),
.B(n_659),
.Y(n_958)
);

NAND2xp33_ASAP7_75t_SL g959 ( 
.A(n_784),
.B(n_664),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_784),
.B(n_670),
.Y(n_960)
);

NAND2x1p5_ASAP7_75t_L g961 ( 
.A(n_931),
.B(n_239),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_943),
.B(n_671),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_850),
.A2(n_676),
.B1(n_688),
.B2(n_672),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_916),
.A2(n_241),
.B(n_240),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_856),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_854),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_947),
.B(n_953),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_SL g968 ( 
.A(n_882),
.B(n_1),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_917),
.A2(n_920),
.B(n_918),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_862),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_883),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_948),
.B(n_1),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_935),
.A2(n_4),
.B(n_2),
.C(n_3),
.Y(n_973)
);

NAND2xp33_ASAP7_75t_L g974 ( 
.A(n_939),
.B(n_242),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_884),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_924),
.B(n_3),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_855),
.B(n_899),
.Y(n_977)
);

AO31x2_ASAP7_75t_L g978 ( 
.A1(n_940),
.A2(n_472),
.A3(n_474),
.B(n_471),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_926),
.A2(n_246),
.B(n_245),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_855),
.B(n_247),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_929),
.B(n_248),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_952),
.B(n_5),
.Y(n_982)
);

OAI21x1_ASAP7_75t_L g983 ( 
.A1(n_927),
.A2(n_252),
.B(n_249),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_928),
.A2(n_254),
.B(n_253),
.Y(n_984)
);

AO22x1_ASAP7_75t_L g985 ( 
.A1(n_887),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_921),
.A2(n_256),
.B1(n_257),
.B2(n_255),
.Y(n_986)
);

OAI21x1_ASAP7_75t_SL g987 ( 
.A1(n_907),
.A2(n_259),
.B(n_258),
.Y(n_987)
);

NAND2x1p5_ASAP7_75t_L g988 ( 
.A(n_931),
.B(n_260),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_913),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_863),
.Y(n_990)
);

AOI21xp33_ASAP7_75t_L g991 ( 
.A1(n_871),
.A2(n_12),
.B(n_13),
.Y(n_991)
);

INVx3_ASAP7_75t_SL g992 ( 
.A(n_902),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_914),
.A2(n_919),
.B(n_932),
.C(n_915),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_946),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_922),
.A2(n_263),
.B(n_261),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_933),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_877),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_923),
.B(n_15),
.Y(n_998)
);

AOI221x1_ASAP7_75t_L g999 ( 
.A1(n_910),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.C(n_20),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_946),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_936),
.A2(n_21),
.B(n_17),
.C(n_18),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_930),
.A2(n_266),
.B(n_265),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_942),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_1003)
);

NOR3xp33_ASAP7_75t_L g1004 ( 
.A(n_875),
.B(n_23),
.C(n_24),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_934),
.A2(n_269),
.B(n_268),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_868),
.Y(n_1006)
);

AO21x1_ASAP7_75t_L g1007 ( 
.A1(n_937),
.A2(n_25),
.B(n_26),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_925),
.A2(n_271),
.B(n_270),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_938),
.A2(n_275),
.B(n_274),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_941),
.B(n_25),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_890),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_SL g1012 ( 
.A1(n_872),
.A2(n_279),
.B(n_280),
.C(n_278),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_873),
.A2(n_283),
.B(n_282),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_L g1014 ( 
.A(n_955),
.B(n_27),
.C(n_28),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_891),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_901),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_889),
.Y(n_1017)
);

AOI221xp5_ASAP7_75t_L g1018 ( 
.A1(n_912),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.C(n_33),
.Y(n_1018)
);

AO31x2_ASAP7_75t_L g1019 ( 
.A1(n_894),
.A2(n_34),
.A3(n_31),
.B(n_33),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_897),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_860),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_851),
.B(n_285),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_959),
.A2(n_287),
.B1(n_288),
.B2(n_286),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_944),
.A2(n_290),
.B1(n_291),
.B2(n_289),
.Y(n_1024)
);

INVxp67_ASAP7_75t_SL g1025 ( 
.A(n_945),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_895),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_853),
.A2(n_294),
.B(n_293),
.Y(n_1027)
);

AO31x2_ASAP7_75t_L g1028 ( 
.A1(n_903),
.A2(n_468),
.A3(n_469),
.B(n_466),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_874),
.A2(n_960),
.B(n_958),
.Y(n_1029)
);

AOI221x1_ASAP7_75t_L g1030 ( 
.A1(n_896),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.C(n_38),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_865),
.B(n_296),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_949),
.A2(n_298),
.B(n_297),
.Y(n_1032)
);

NAND2xp33_ASAP7_75t_R g1033 ( 
.A(n_893),
.B(n_299),
.Y(n_1033)
);

NOR2x1_ASAP7_75t_SL g1034 ( 
.A(n_857),
.B(n_300),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_SL g1035 ( 
.A1(n_892),
.A2(n_303),
.B(n_302),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_858),
.A2(n_861),
.B(n_859),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_848),
.B(n_36),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_950),
.B(n_39),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_951),
.A2(n_308),
.B1(n_310),
.B2(n_305),
.Y(n_1039)
);

XOR2xp5_ASAP7_75t_L g1040 ( 
.A(n_954),
.B(n_311),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_864),
.A2(n_867),
.B(n_866),
.Y(n_1041)
);

OA21x2_ASAP7_75t_L g1042 ( 
.A1(n_969),
.A2(n_869),
.B(n_956),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_SL g1043 ( 
.A1(n_1013),
.A2(n_957),
.B(n_870),
.Y(n_1043)
);

OA21x2_ASAP7_75t_L g1044 ( 
.A1(n_1041),
.A2(n_879),
.B(n_878),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_966),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_965),
.B(n_876),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_962),
.A2(n_852),
.B1(n_906),
.B2(n_905),
.Y(n_1047)
);

OAI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_967),
.A2(n_904),
.B1(n_909),
.B2(n_911),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_970),
.Y(n_1049)
);

OAI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_997),
.A2(n_908),
.B1(n_849),
.B2(n_885),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_1020),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_983),
.A2(n_888),
.B(n_886),
.Y(n_1052)
);

OA21x2_ASAP7_75t_L g1053 ( 
.A1(n_979),
.A2(n_1005),
.B(n_984),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1021),
.B(n_898),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_972),
.A2(n_880),
.B(n_900),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_971),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_976),
.B(n_881),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_975),
.Y(n_1058)
);

NAND3xp33_ASAP7_75t_SL g1059 ( 
.A(n_1004),
.B(n_41),
.C(n_42),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_1002),
.A2(n_313),
.B(n_312),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1006),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_990),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1007),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_1000),
.B(n_977),
.Y(n_1064)
);

AOI221xp5_ASAP7_75t_L g1065 ( 
.A1(n_991),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.C(n_45),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_1009),
.A2(n_318),
.B(n_317),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_1010),
.A2(n_50),
.B1(n_46),
.B2(n_48),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_1017),
.Y(n_1068)
);

AOI21x1_ASAP7_75t_L g1069 ( 
.A1(n_1036),
.A2(n_321),
.B(n_320),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_982),
.B(n_1015),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1038),
.Y(n_1071)
);

AO21x1_ASAP7_75t_L g1072 ( 
.A1(n_1032),
.A2(n_1031),
.B(n_1016),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_980),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1029),
.A2(n_328),
.B(n_327),
.Y(n_1074)
);

NAND2x1_ASAP7_75t_L g1075 ( 
.A(n_1035),
.B(n_330),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_961),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_998),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_1025),
.B(n_333),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_988),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1026),
.B(n_51),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_993),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_1022),
.B(n_334),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_978),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_1037),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_1014),
.A2(n_1018),
.B1(n_968),
.B2(n_1040),
.Y(n_1085)
);

OA21x2_ASAP7_75t_L g1086 ( 
.A1(n_981),
.A2(n_336),
.B(n_335),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_SL g1087 ( 
.A1(n_1034),
.A2(n_342),
.B(n_341),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_963),
.B(n_55),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_964),
.A2(n_345),
.B(n_343),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1019),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_1019),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_1028),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_1019),
.Y(n_1093)
);

AO31x2_ASAP7_75t_L g1094 ( 
.A1(n_973),
.A2(n_996),
.A3(n_1001),
.B(n_989),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_SL g1095 ( 
.A1(n_1027),
.A2(n_347),
.B(n_346),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_974),
.A2(n_352),
.B(n_349),
.Y(n_1096)
);

CKINVDCx16_ASAP7_75t_R g1097 ( 
.A(n_1033),
.Y(n_1097)
);

NAND2xp33_ASAP7_75t_L g1098 ( 
.A(n_1003),
.B(n_353),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_1024),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_995),
.A2(n_355),
.B(n_354),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_985),
.B(n_1039),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1012),
.A2(n_358),
.B(n_357),
.Y(n_1102)
);

NOR2x1_ASAP7_75t_SL g1103 ( 
.A(n_986),
.B(n_359),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_1023),
.B(n_360),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_1008),
.B(n_361),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_978),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_967),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_1107)
);

AOI21xp33_ASAP7_75t_SL g1108 ( 
.A1(n_992),
.A2(n_61),
.B(n_62),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_965),
.Y(n_1109)
);

AO21x1_ASAP7_75t_L g1110 ( 
.A1(n_967),
.A2(n_65),
.B(n_64),
.Y(n_1110)
);

AND2x6_ASAP7_75t_L g1111 ( 
.A(n_1022),
.B(n_362),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_1030),
.A2(n_367),
.A3(n_368),
.B(n_365),
.Y(n_1112)
);

AO32x2_ASAP7_75t_L g1113 ( 
.A1(n_999),
.A2(n_65),
.A3(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_962),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_983),
.A2(n_370),
.B(n_369),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_994),
.B(n_371),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1011),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_965),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_L g1119 ( 
.A(n_962),
.B(n_67),
.C(n_68),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_SL g1120 ( 
.A1(n_987),
.A2(n_374),
.B(n_373),
.Y(n_1120)
);

NOR2xp67_ASAP7_75t_L g1121 ( 
.A(n_975),
.B(n_375),
.Y(n_1121)
);

AOI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1106),
.A2(n_378),
.B(n_376),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_1118),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_1064),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1062),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1045),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_1051),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_1079),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_1116),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_1109),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_1073),
.B(n_379),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1049),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1061),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1058),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1117),
.Y(n_1135)
);

AOI221xp5_ASAP7_75t_SL g1136 ( 
.A1(n_1088),
.A2(n_74),
.B1(n_70),
.B2(n_72),
.C(n_76),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1076),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1046),
.B(n_76),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1071),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1077),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_1068),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1090),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1093),
.Y(n_1143)
);

AOI221xp5_ASAP7_75t_L g1144 ( 
.A1(n_1085),
.A2(n_1048),
.B1(n_1059),
.B2(n_1099),
.C(n_1101),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1063),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1091),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_1078),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_1105),
.Y(n_1148)
);

OA21x2_ASAP7_75t_L g1149 ( 
.A1(n_1083),
.A2(n_382),
.B(n_381),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1070),
.B(n_77),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1097),
.B(n_77),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1056),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1042),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_1054),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1075),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1094),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_1086),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1069),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_1084),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1047),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1082),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_1080),
.B(n_80),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1050),
.B(n_81),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_1111),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1113),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1067),
.B(n_1114),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1060),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1066),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_1057),
.B(n_82),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1110),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1104),
.B(n_83),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_1129),
.B(n_1121),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1144),
.B(n_1072),
.Y(n_1173)
);

INVxp67_ASAP7_75t_L g1174 ( 
.A(n_1130),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1141),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_1161),
.B(n_1108),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1147),
.B(n_1119),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_1154),
.Y(n_1178)
);

BUFx10_ASAP7_75t_L g1179 ( 
.A(n_1127),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_R g1180 ( 
.A(n_1161),
.B(n_1098),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_R g1181 ( 
.A(n_1147),
.B(n_1092),
.Y(n_1181)
);

INVxp67_ASAP7_75t_L g1182 ( 
.A(n_1123),
.Y(n_1182)
);

CKINVDCx16_ASAP7_75t_R g1183 ( 
.A(n_1151),
.Y(n_1183)
);

NAND2xp33_ASAP7_75t_R g1184 ( 
.A(n_1134),
.B(n_1169),
.Y(n_1184)
);

NAND2xp33_ASAP7_75t_R g1185 ( 
.A(n_1150),
.B(n_1044),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1138),
.B(n_1081),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1142),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1126),
.Y(n_1188)
);

OR2x6_ASAP7_75t_L g1189 ( 
.A(n_1164),
.B(n_1043),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1124),
.B(n_1055),
.Y(n_1190)
);

NAND2xp33_ASAP7_75t_R g1191 ( 
.A(n_1163),
.B(n_1053),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1171),
.B(n_1107),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1148),
.B(n_1052),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1139),
.B(n_1065),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1128),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1140),
.B(n_1074),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_1131),
.B(n_1089),
.Y(n_1197)
);

OR2x6_ASAP7_75t_L g1198 ( 
.A(n_1159),
.B(n_1120),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1132),
.Y(n_1199)
);

OAI221xp5_ASAP7_75t_L g1200 ( 
.A1(n_1192),
.A2(n_1136),
.B1(n_1160),
.B2(n_1162),
.C(n_1166),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1187),
.Y(n_1201)
);

AND2x4_ASAP7_75t_SL g1202 ( 
.A(n_1179),
.B(n_1137),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1188),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1178),
.B(n_1146),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1199),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1182),
.Y(n_1206)
);

NAND2x1p5_ASAP7_75t_SL g1207 ( 
.A(n_1173),
.B(n_1153),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_1175),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1193),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1183),
.B(n_1135),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1174),
.B(n_1177),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1196),
.B(n_1125),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1195),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1186),
.B(n_1190),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1194),
.B(n_1143),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1181),
.Y(n_1216)
);

OR2x2_ASAP7_75t_L g1217 ( 
.A(n_1189),
.B(n_1145),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1189),
.B(n_1156),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1176),
.B(n_1170),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1197),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1198),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1185),
.Y(n_1222)
);

NOR2xp67_ASAP7_75t_L g1223 ( 
.A(n_1172),
.B(n_1152),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1180),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1191),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1184),
.B(n_1133),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1203),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1205),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1211),
.B(n_1165),
.Y(n_1229)
);

AO21x2_ASAP7_75t_L g1230 ( 
.A1(n_1225),
.A2(n_1122),
.B(n_1158),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1201),
.Y(n_1231)
);

INVxp67_ASAP7_75t_SL g1232 ( 
.A(n_1222),
.Y(n_1232)
);

OAI221xp5_ASAP7_75t_SL g1233 ( 
.A1(n_1200),
.A2(n_1102),
.B1(n_1155),
.B2(n_1168),
.C(n_1167),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1201),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1224),
.A2(n_1096),
.B1(n_1149),
.B2(n_1157),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1209),
.Y(n_1236)
);

AND2x2_ASAP7_75t_SL g1237 ( 
.A(n_1216),
.B(n_1149),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1206),
.B(n_1112),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1204),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1209),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1208),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1214),
.B(n_1112),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1215),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1217),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1220),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1212),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1219),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1226),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1218),
.Y(n_1249)
);

INVx2_ASAP7_75t_SL g1250 ( 
.A(n_1202),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1224),
.B(n_1115),
.Y(n_1251)
);

NOR2x1_ASAP7_75t_SL g1252 ( 
.A(n_1207),
.B(n_1103),
.Y(n_1252)
);

OR2x2_ASAP7_75t_SL g1253 ( 
.A(n_1213),
.B(n_84),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_1221),
.B(n_1100),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1203),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1210),
.B(n_84),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1203),
.Y(n_1257)
);

INVx5_ASAP7_75t_L g1258 ( 
.A(n_1216),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1201),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1201),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1210),
.B(n_87),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1223),
.B(n_1087),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1259),
.Y(n_1263)
);

OR2x6_ASAP7_75t_L g1264 ( 
.A(n_1250),
.B(n_1095),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1236),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1240),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1244),
.B(n_88),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1247),
.B(n_91),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1231),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1246),
.B(n_1243),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1258),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1232),
.B(n_91),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1234),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1260),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1239),
.B(n_92),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1227),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1249),
.B(n_93),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1228),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1229),
.B(n_96),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1255),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1257),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1245),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1241),
.B(n_98),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1233),
.A2(n_1237),
.B(n_1262),
.C(n_1235),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1242),
.B(n_99),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1238),
.B(n_100),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1230),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1251),
.B(n_101),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1256),
.B(n_102),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1261),
.B(n_102),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1254),
.B(n_103),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1252),
.B(n_104),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1253),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1259),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1249),
.B(n_105),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1249),
.B(n_106),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1259),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_1248),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1263),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1298),
.B(n_106),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1271),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1270),
.B(n_109),
.Y(n_1302)
);

NAND2xp33_ASAP7_75t_SL g1303 ( 
.A(n_1295),
.B(n_110),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1295),
.Y(n_1304)
);

AO221x2_ASAP7_75t_L g1305 ( 
.A1(n_1291),
.A2(n_1288),
.B1(n_1286),
.B2(n_1265),
.C(n_1266),
.Y(n_1305)
);

NAND2xp33_ASAP7_75t_SL g1306 ( 
.A(n_1296),
.B(n_1272),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1289),
.B(n_111),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1281),
.B(n_112),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1282),
.B(n_113),
.Y(n_1309)
);

XNOR2xp5_ASAP7_75t_L g1310 ( 
.A(n_1290),
.B(n_114),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1276),
.B(n_115),
.Y(n_1311)
);

INVxp67_ASAP7_75t_L g1312 ( 
.A(n_1292),
.Y(n_1312)
);

INVx5_ASAP7_75t_L g1313 ( 
.A(n_1277),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1278),
.B(n_118),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1294),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1280),
.B(n_121),
.Y(n_1316)
);

BUFx12f_ASAP7_75t_L g1317 ( 
.A(n_1283),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1264),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_1318)
);

NOR2x1_ASAP7_75t_L g1319 ( 
.A(n_1287),
.B(n_126),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1267),
.B(n_126),
.Y(n_1320)
);

AO221x2_ASAP7_75t_L g1321 ( 
.A1(n_1297),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.C(n_130),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1285),
.B(n_131),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1274),
.B(n_131),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1269),
.B(n_132),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1273),
.B(n_133),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1279),
.B(n_134),
.Y(n_1326)
);

NAND2xp33_ASAP7_75t_SL g1327 ( 
.A(n_1268),
.B(n_136),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1275),
.B(n_137),
.Y(n_1328)
);

NOR2x1_ASAP7_75t_L g1329 ( 
.A(n_1284),
.B(n_141),
.Y(n_1329)
);

NAND2xp33_ASAP7_75t_SL g1330 ( 
.A(n_1293),
.B(n_143),
.Y(n_1330)
);

OAI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1293),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_1331)
);

NOR2x1_ASAP7_75t_L g1332 ( 
.A(n_1284),
.B(n_145),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1293),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1298),
.B(n_150),
.Y(n_1334)
);

AO21x2_ASAP7_75t_L g1335 ( 
.A1(n_1300),
.A2(n_152),
.B(n_153),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1317),
.Y(n_1336)
);

AO22x1_ASAP7_75t_L g1337 ( 
.A1(n_1332),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1315),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1313),
.B(n_159),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1301),
.B(n_160),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1324),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1325),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1330),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1311),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1304),
.B(n_163),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1314),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1316),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1323),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1308),
.B(n_164),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1309),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1334),
.B(n_166),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1327),
.Y(n_1352)
);

INVxp67_ASAP7_75t_L g1353 ( 
.A(n_1307),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1302),
.B(n_167),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1322),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1328),
.B(n_169),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1326),
.Y(n_1357)
);

AO21x2_ASAP7_75t_L g1358 ( 
.A1(n_1331),
.A2(n_1333),
.B(n_1310),
.Y(n_1358)
);

INVx1_ASAP7_75t_SL g1359 ( 
.A(n_1303),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1321),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1320),
.B(n_170),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1318),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1305),
.B(n_172),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1305),
.B(n_173),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1299),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1299),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1299),
.Y(n_1367)
);

INVxp67_ASAP7_75t_SL g1368 ( 
.A(n_1319),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_1306),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1313),
.B(n_175),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1306),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1299),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1305),
.B(n_176),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1299),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1299),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1312),
.B(n_178),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1312),
.B(n_179),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1329),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_1378)
);

BUFx2_ASAP7_75t_SL g1379 ( 
.A(n_1313),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1329),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1368),
.B(n_188),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1362),
.B(n_189),
.Y(n_1382)
);

AOI211xp5_ASAP7_75t_L g1383 ( 
.A1(n_1337),
.A2(n_192),
.B(n_190),
.C(n_191),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1355),
.B(n_194),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1357),
.B(n_194),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1336),
.Y(n_1386)
);

AOI22x1_ASAP7_75t_L g1387 ( 
.A1(n_1379),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1363),
.B(n_199),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1365),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1366),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1367),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1364),
.B(n_203),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1369),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_1393)
);

AOI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1371),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_1394)
);

AOI21xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1358),
.A2(n_210),
.B(n_211),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1372),
.Y(n_1396)
);

O2A1O1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1373),
.A2(n_214),
.B(n_212),
.C(n_213),
.Y(n_1397)
);

AOI322xp5_ASAP7_75t_L g1398 ( 
.A1(n_1360),
.A2(n_215),
.A3(n_216),
.B1(n_217),
.B2(n_218),
.C1(n_219),
.C2(n_220),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1374),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1370),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1375),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1352),
.B(n_221),
.Y(n_1402)
);

NOR2x1_ASAP7_75t_L g1403 ( 
.A(n_1339),
.B(n_222),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1343),
.A2(n_223),
.B(n_224),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1359),
.A2(n_1380),
.B(n_1378),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1338),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1341),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1342),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1344),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1346),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1347),
.Y(n_1411)
);

OAI211xp5_ASAP7_75t_SL g1412 ( 
.A1(n_1350),
.A2(n_229),
.B(n_227),
.C(n_228),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1348),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1376),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1335),
.B(n_231),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1353),
.B(n_234),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1395),
.B(n_1351),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1386),
.Y(n_1418)
);

NOR2x1_ASAP7_75t_L g1419 ( 
.A(n_1403),
.B(n_1340),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1400),
.B(n_1377),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1382),
.B(n_1354),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1389),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1414),
.B(n_1345),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1405),
.B(n_1349),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1390),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1391),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1397),
.B(n_1356),
.Y(n_1427)
);

NOR2x1_ASAP7_75t_L g1428 ( 
.A(n_1381),
.B(n_1361),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1396),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1399),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1388),
.B(n_1392),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1401),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1404),
.B(n_389),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1407),
.B(n_390),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1406),
.B(n_391),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_1419),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1418),
.Y(n_1437)
);

INVx8_ASAP7_75t_L g1438 ( 
.A(n_1423),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1422),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1423),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1417),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1425),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1426),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1429),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1430),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1432),
.Y(n_1446)
);

NAND3xp33_ASAP7_75t_L g1447 ( 
.A(n_1436),
.B(n_1383),
.C(n_1398),
.Y(n_1447)
);

OAI21xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1441),
.A2(n_1424),
.B(n_1427),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1438),
.Y(n_1449)
);

OAI211xp5_ASAP7_75t_L g1450 ( 
.A1(n_1437),
.A2(n_1387),
.B(n_1394),
.C(n_1393),
.Y(n_1450)
);

NOR2x1_ASAP7_75t_L g1451 ( 
.A(n_1440),
.B(n_1415),
.Y(n_1451)
);

XOR2x2_ASAP7_75t_L g1452 ( 
.A(n_1447),
.B(n_1428),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1451),
.Y(n_1453)
);

NOR2x1_ASAP7_75t_L g1454 ( 
.A(n_1449),
.B(n_1402),
.Y(n_1454)
);

NOR3xp33_ASAP7_75t_L g1455 ( 
.A(n_1448),
.B(n_1431),
.C(n_1439),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1454),
.B(n_1420),
.Y(n_1456)
);

NAND2x1p5_ASAP7_75t_L g1457 ( 
.A(n_1453),
.B(n_1435),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1452),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1456),
.B(n_1455),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_R g1460 ( 
.A(n_1458),
.B(n_1433),
.Y(n_1460)
);

NAND3xp33_ASAP7_75t_SL g1461 ( 
.A(n_1459),
.B(n_1457),
.C(n_1450),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1461),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1462),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1463),
.A2(n_1460),
.B1(n_1442),
.B2(n_1444),
.Y(n_1464)
);

NAND5xp2_ASAP7_75t_L g1465 ( 
.A(n_1464),
.B(n_1445),
.C(n_1446),
.D(n_1443),
.E(n_1421),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1465),
.A2(n_1412),
.B1(n_1409),
.B2(n_1410),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1466),
.Y(n_1467)
);

AOI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1467),
.A2(n_1434),
.B1(n_1385),
.B2(n_1384),
.C(n_1411),
.Y(n_1468)
);

AOI211xp5_ASAP7_75t_L g1469 ( 
.A1(n_1468),
.A2(n_1416),
.B(n_1413),
.C(n_1408),
.Y(n_1469)
);


endmodule