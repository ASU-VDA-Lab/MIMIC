module fake_jpeg_30482_n_391 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_391);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_391;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_18),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_9),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_55),
.Y(n_88)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_23),
.B(n_8),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_53),
.B(n_56),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_8),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_23),
.B(n_10),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_34),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_73),
.Y(n_80)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_24),
.B(n_10),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_60),
.B(n_69),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_39),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g115 ( 
.A(n_62),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_63),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_24),
.B(n_7),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_70),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_46),
.B(n_0),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_37),
.B(n_7),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_30),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_30),
.B(n_12),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_44),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_25),
.B1(n_43),
.B2(n_27),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_81),
.A2(n_89),
.B1(n_93),
.B2(n_108),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_87),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_85),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_88),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_25),
.B1(n_27),
.B2(n_35),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_59),
.A2(n_25),
.B1(n_26),
.B2(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_R g96 ( 
.A(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_96),
.B(n_14),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_22),
.B1(n_47),
.B2(n_33),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_99),
.A2(n_38),
.B1(n_32),
.B2(n_14),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_26),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_107),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_31),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_31),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_72),
.A2(n_39),
.B1(n_32),
.B2(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_40),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_111),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_79),
.B1(n_78),
.B2(n_44),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_121),
.A2(n_132),
.B1(n_141),
.B2(n_149),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_40),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_128),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_129),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_36),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_126),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_96),
.A2(n_39),
.B1(n_48),
.B2(n_47),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_22),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_99),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_139),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_65),
.B1(n_48),
.B2(n_29),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_142),
.Y(n_175)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_137),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_88),
.B(n_36),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_117),
.C(n_95),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_88),
.B(n_33),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_145),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_91),
.A2(n_29),
.B1(n_39),
.B2(n_36),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_143),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_104),
.B(n_16),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_150),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_91),
.A2(n_36),
.B(n_32),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_19),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_95),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_109),
.A2(n_38),
.B1(n_32),
.B2(n_16),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_94),
.A2(n_38),
.B1(n_6),
.B2(n_17),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_32),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_156),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_38),
.B1(n_6),
.B2(n_17),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_114),
.B1(n_90),
.B2(n_113),
.Y(n_157)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_105),
.Y(n_180)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_157),
.A2(n_150),
.B1(n_122),
.B2(n_141),
.Y(n_188)
);

OA22x2_ASAP7_75t_SL g158 ( 
.A1(n_147),
.A2(n_90),
.B1(n_105),
.B2(n_38),
.Y(n_158)
);

OR2x4_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_154),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_120),
.B(n_112),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_159),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_185),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_153),
.B(n_123),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_171),
.B(n_178),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_120),
.B(n_112),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_115),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_128),
.B(n_19),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g179 ( 
.A(n_155),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_179),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_125),
.B(n_115),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_181),
.B(n_138),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_145),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_139),
.B(n_124),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_137),
.B1(n_134),
.B2(n_156),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_188),
.A2(n_196),
.B1(n_210),
.B2(n_159),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_189),
.B(n_199),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_125),
.C(n_126),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_198),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_205),
.Y(n_227)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_121),
.B1(n_132),
.B2(n_152),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_197),
.B1(n_209),
.B2(n_159),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_186),
.A2(n_161),
.B1(n_176),
.B2(n_168),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_138),
.B1(n_149),
.B2(n_126),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_201),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_161),
.A2(n_138),
.B(n_148),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_162),
.B(n_181),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_155),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_146),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_212),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_180),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_207),
.B(n_208),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_158),
.A2(n_116),
.B1(n_92),
.B2(n_133),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_151),
.C(n_140),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_184),
.C(n_198),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_193),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_213),
.B(n_218),
.Y(n_245)
);

NOR2x1_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_161),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_224),
.Y(n_241)
);

CKINVDCx12_ASAP7_75t_R g216 ( 
.A(n_204),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_216),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_236),
.C(n_197),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_178),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_184),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_219),
.A2(n_228),
.B(n_231),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_212),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_222),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_230),
.B1(n_158),
.B2(n_180),
.Y(n_259)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_187),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_187),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_210),
.A2(n_159),
.B1(n_182),
.B2(n_158),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_198),
.A2(n_161),
.B(n_164),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_202),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_234),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_159),
.C(n_172),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_168),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_237),
.A2(n_238),
.B(n_194),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_158),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_190),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_242),
.C(n_248),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_190),
.Y(n_242)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_227),
.B(n_192),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_247),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_191),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_216),
.A2(n_209),
.B(n_200),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_249),
.A2(n_266),
.B(n_231),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_251),
.C(n_253),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_169),
.C(n_200),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_207),
.Y(n_252)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_219),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_169),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_256),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_165),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_224),
.A2(n_188),
.B1(n_209),
.B2(n_195),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_230),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_259),
.A2(n_174),
.B1(n_166),
.B2(n_157),
.Y(n_286)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_214),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_263),
.Y(n_282)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_214),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_220),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_228),
.A2(n_165),
.B(n_202),
.Y(n_266)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_269),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_272),
.A2(n_276),
.B1(n_281),
.B2(n_280),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_252),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_274),
.B(n_286),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_258),
.A2(n_225),
.B1(n_238),
.B2(n_222),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_276),
.A2(n_280),
.B1(n_281),
.B2(n_287),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_277),
.A2(n_284),
.B(n_285),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_265),
.A2(n_232),
.B1(n_233),
.B2(n_163),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_235),
.Y(n_279)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_262),
.A2(n_238),
.B1(n_237),
.B2(n_215),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_262),
.A2(n_237),
.B1(n_215),
.B2(n_213),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_206),
.Y(n_283)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_232),
.Y(n_284)
);

NAND2x1_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_174),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_241),
.A2(n_160),
.B1(n_166),
.B2(n_183),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_241),
.A2(n_160),
.B(n_117),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_288),
.A2(n_289),
.B(n_244),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_249),
.A2(n_163),
.B(n_117),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_277),
.B(n_253),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_294),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_293),
.A2(n_286),
.B1(n_290),
.B2(n_285),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_250),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_268),
.B(n_266),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_296),
.B(n_301),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_240),
.C(n_251),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_300),
.C(n_303),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_248),
.C(n_242),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_268),
.B(n_264),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_270),
.B(n_244),
.C(n_246),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_305),
.A2(n_289),
.B(n_272),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_256),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_312),
.C(n_271),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_267),
.Y(n_307)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_307),
.Y(n_314)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_282),
.Y(n_308)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_309),
.Y(n_327)
);

MAJx2_ASAP7_75t_L g312 ( 
.A(n_273),
.B(n_243),
.C(n_254),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_271),
.CI(n_274),
.CON(n_313),
.SN(n_313)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_313),
.B(n_316),
.Y(n_346)
);

NAND4xp25_ASAP7_75t_SL g316 ( 
.A(n_298),
.B(n_267),
.C(n_245),
.D(n_284),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_272),
.B1(n_287),
.B2(n_290),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_317),
.A2(n_331),
.B1(n_170),
.B2(n_183),
.Y(n_344)
);

INVxp33_ASAP7_75t_SL g319 ( 
.A(n_295),
.Y(n_319)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_319),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_294),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_326),
.Y(n_333)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_297),
.Y(n_324)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_324),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_299),
.B(n_203),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_325),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_310),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_328),
.A2(n_239),
.B1(n_267),
.B2(n_255),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_273),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_329),
.A2(n_284),
.B(n_261),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_304),
.B(n_203),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_330),
.B(n_304),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_311),
.A2(n_275),
.B1(n_285),
.B2(n_263),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_335),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_334),
.B(n_344),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_293),
.Y(n_335)
);

AOI322xp5_ASAP7_75t_SL g336 ( 
.A1(n_322),
.A2(n_292),
.A3(n_312),
.B1(n_303),
.B2(n_302),
.C1(n_300),
.C2(n_275),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_336),
.B(n_313),
.Y(n_357)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_338),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_260),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_340),
.B(n_342),
.C(n_345),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_315),
.B(n_260),
.C(n_239),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_343),
.B(n_324),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_320),
.B(n_170),
.C(n_173),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_329),
.B(n_317),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_347),
.A2(n_354),
.B(n_357),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_344),
.A2(n_323),
.B1(n_327),
.B2(n_318),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_349),
.A2(n_333),
.B1(n_345),
.B2(n_314),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_339),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_356),
.Y(n_365)
);

INVx11_ASAP7_75t_L g352 ( 
.A(n_337),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_352),
.B(n_341),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_342),
.B(n_320),
.C(n_331),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_338),
.A2(n_326),
.B1(n_313),
.B2(n_316),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_358),
.Y(n_363)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_360),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_352),
.B(n_340),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_362),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_347),
.A2(n_335),
.B(n_334),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_364),
.A2(n_349),
.B1(n_82),
.B2(n_19),
.Y(n_376)
);

AOI221xp5_ASAP7_75t_L g366 ( 
.A1(n_356),
.A2(n_333),
.B1(n_167),
.B2(n_170),
.C(n_144),
.Y(n_366)
);

OAI221xp5_ASAP7_75t_L g378 ( 
.A1(n_366),
.A2(n_368),
.B1(n_18),
.B2(n_20),
.C(n_5),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_183),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_367),
.B(n_350),
.Y(n_370)
);

OAI221xp5_ASAP7_75t_L g368 ( 
.A1(n_348),
.A2(n_173),
.B1(n_133),
.B2(n_136),
.C(n_18),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_136),
.C(n_142),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_369),
.B(n_354),
.C(n_353),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_370),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_371),
.A2(n_372),
.B(n_373),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_355),
.C(n_353),
.Y(n_372)
);

AO21x1_ASAP7_75t_L g373 ( 
.A1(n_365),
.A2(n_348),
.B(n_358),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_376),
.A2(n_377),
.B(n_378),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_363),
.A2(n_119),
.B1(n_92),
.B2(n_116),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_374),
.A2(n_363),
.B(n_366),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_381),
.C(n_370),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_375),
.A2(n_142),
.B(n_131),
.Y(n_381)
);

NOR3xp33_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_110),
.C(n_5),
.Y(n_384)
);

AOI21x1_ASAP7_75t_SL g386 ( 
.A1(n_384),
.A2(n_20),
.B(n_1),
.Y(n_386)
);

AOI322xp5_ASAP7_75t_L g388 ( 
.A1(n_385),
.A2(n_386),
.A3(n_387),
.B1(n_383),
.B2(n_382),
.C1(n_110),
.C2(n_3),
.Y(n_388)
);

AOI321xp33_ASAP7_75t_L g387 ( 
.A1(n_380),
.A2(n_131),
.A3(n_82),
.B1(n_110),
.B2(n_95),
.C(n_0),
.Y(n_387)
);

OAI22xp33_ASAP7_75t_L g390 ( 
.A1(n_388),
.A2(n_389),
.B1(n_3),
.B2(n_1),
.Y(n_390)
);

AOI322xp5_ASAP7_75t_L g389 ( 
.A1(n_385),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_383),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_390),
.B(n_3),
.Y(n_391)
);


endmodule