module real_jpeg_3943_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_11;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_9;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_4),
.B(n_14),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_4),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_4),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_4),
.B(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_40),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_38),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_25),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_11),
.B(n_25),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_17),
.C(n_21),
.Y(n_11)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_12),
.A2(n_13),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_12),
.A2(n_13),
.B1(n_17),
.B2(n_54),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_21),
.A2(n_44),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_21),
.A2(n_44),
.B1(n_45),
.B2(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_57),
.C(n_58),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_22),
.A2(n_46),
.B1(n_57),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_22),
.Y(n_80)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_89),
.Y(n_40)
);

NAND3xp33_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_55),
.C(n_70),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_42),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_51),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_43),
.B(n_51),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.C(n_46),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_57),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_47),
.A2(n_73),
.B(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_66),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_66),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_58),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_59),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_83),
.B(n_88),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);


endmodule