module real_jpeg_17517_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_470;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_215;
wire n_286;
wire n_176;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_500),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_0),
.B(n_501),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_1),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_1),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g149 ( 
.A(n_1),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_1),
.B(n_41),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_1),
.B(n_62),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_1),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_1),
.B(n_174),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_2),
.B(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_2),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_2),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_2),
.B(n_362),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_2),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_2),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_2),
.B(n_423),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_3),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_3),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g360 ( 
.A(n_3),
.Y(n_360)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_4),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_4),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_4),
.Y(n_224)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_4),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_5),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_5),
.B(n_96),
.Y(n_95)
);

AND2x4_ASAP7_75t_L g155 ( 
.A(n_5),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_5),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_5),
.B(n_262),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_5),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_5),
.B(n_75),
.Y(n_455)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g369 ( 
.A(n_6),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_7),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_7),
.A2(n_8),
.B1(n_64),
.B2(n_69),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_7),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_7),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_7),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_7),
.B(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_7),
.B(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_8),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_8),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_8),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_8),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_8),
.B(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_8),
.B(n_496),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_9),
.Y(n_85)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_9),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_9),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_9),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_9),
.Y(n_217)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_10),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_10),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_10),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_10),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_10),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_10),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_10),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_10),
.B(n_369),
.Y(n_368)
);

INVxp33_ASAP7_75t_L g501 ( 
.A(n_11),
.Y(n_501)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_12),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_12),
.Y(n_148)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_12),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_13),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_13),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_13),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_13),
.B(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_13),
.B(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_13),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_15),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_15),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_15),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_15),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_15),
.B(n_336),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_15),
.B(n_420),
.Y(n_419)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_16),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g374 ( 
.A(n_16),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_16),
.Y(n_408)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g174 ( 
.A(n_17),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_17),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_17),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_471),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_440),
.B(n_470),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2x1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_323),
.Y(n_22)
);

A2O1A1O1Ixp25_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_237),
.B(n_286),
.C(n_287),
.D(n_322),
.Y(n_23)
);

OAI21x1_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_186),
.B(n_236),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_139),
.Y(n_25)
);

NOR2xp67_ASAP7_75t_SL g439 ( 
.A(n_26),
.B(n_139),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_87),
.C(n_123),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_27),
.B(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_49),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_28),
.B(n_50),
.C(n_73),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_37),
.C(n_43),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_29),
.B(n_331),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_30),
.A2(n_176),
.B1(n_177),
.B2(n_180),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_30),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_30),
.B(n_173),
.C(n_177),
.Y(n_198)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_32),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_33),
.A2(n_232),
.B1(n_233),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_33),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_33),
.B(n_233),
.C(n_268),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_33),
.A2(n_108),
.B1(n_127),
.B2(n_273),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_33),
.B(n_180),
.Y(n_333)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_37),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_331)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_48),
.Y(n_220)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_48),
.Y(n_315)
);

INVx3_ASAP7_75t_SL g498 ( 
.A(n_48),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_73),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_59),
.B(n_63),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_52),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_52),
.B(n_229),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_57),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_62),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_63),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_63),
.Y(n_183)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_70),
.B(n_310),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_71),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_72),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_74),
.B(n_79),
.C(n_82),
.Y(n_168)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_77),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B1(n_82),
.B2(n_86),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_79),
.B(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_81),
.A2(n_82),
.B1(n_108),
.B2(n_127),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_81),
.A2(n_82),
.B1(n_149),
.B2(n_153),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_82),
.B(n_127),
.C(n_463),
.Y(n_483)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_86),
.B(n_278),
.C(n_283),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_87),
.A2(n_88),
.B1(n_123),
.B2(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_112),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_99),
.B2(n_100),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_90),
.B(n_100),
.C(n_112),
.Y(n_169)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_95),
.A2(n_129),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_96),
.Y(n_119)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJx2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.C(n_108),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_108),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_125),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_106),
.Y(n_282)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_106),
.Y(n_392)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_108),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_108),
.B(n_273),
.C(n_309),
.Y(n_467)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_110),
.Y(n_166)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_111),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_113),
.B(n_117),
.C(n_120),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_123),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.C(n_130),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_124),
.B(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_128),
.B(n_130),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_129),
.B(n_228),
.C(n_233),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.C(n_137),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_131),
.B(n_137),
.Y(n_381)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_134),
.B(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_170),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_171),
.C(n_185),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_169),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_159),
.Y(n_141)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_154),
.B2(n_155),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_144)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_145),
.B(n_153),
.C(n_154),
.Y(n_226)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_154),
.A2(n_155),
.B1(n_317),
.B2(n_321),
.Y(n_316)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_155),
.B(n_314),
.C(n_321),
.Y(n_466)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx6_ASAP7_75t_L g365 ( 
.A(n_158),
.Y(n_365)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_168),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_164),
.B1(n_165),
.B2(n_167),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_161),
.A2(n_165),
.B(n_168),
.C(n_208),
.Y(n_207)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_190),
.C(n_191),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_185),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_181),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_183),
.C(n_184),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_178),
.Y(n_342)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

NOR2x1_ASAP7_75t_L g438 ( 
.A(n_186),
.B(n_439),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_187),
.B(n_188),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_189),
.B(n_239),
.C(n_240),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_211),
.B2(n_212),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_195),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_196)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_206),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_198),
.Y(n_206)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_201),
.B(n_206),
.C(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_203),
.Y(n_338)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_204),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_207),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_243),
.C(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_225),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_226),
.C(n_234),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g263 ( 
.A(n_214),
.B(n_219),
.C(n_221),
.Y(n_263)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_220),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_221),
.A2(n_451),
.B1(n_452),
.B2(n_453),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_221),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_221),
.B(n_452),
.C(n_455),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_223),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_224),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_234),
.B2(n_235),
.Y(n_225)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_226),
.Y(n_235)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_227),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_232),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_232),
.B(n_340),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_233),
.B(n_340),
.Y(n_339)
);

NAND4xp25_ASAP7_75t_L g323 ( 
.A(n_237),
.B(n_287),
.C(n_324),
.D(n_438),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_238),
.B(n_241),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_242),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_266),
.B1(n_284),
.B2(n_285),
.Y(n_245)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_265),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_247),
.B(n_250),
.C(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_254),
.B2(n_264),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_263),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_260),
.B2(n_261),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_260),
.C(n_263),
.Y(n_298)
);

BUFx12f_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_260),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_260),
.A2(n_459),
.B1(n_494),
.B2(n_495),
.Y(n_493)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_261),
.B(n_301),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_264),
.Y(n_292)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_284),
.C(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_274),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_275),
.C(n_276),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_272),
.Y(n_267)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_283),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_281),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_290),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_291),
.B(n_306),
.C(n_469),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_306),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_294),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_305),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_295),
.B(n_298),
.C(n_299),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

AO22x1_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_299)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_301),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_302),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_304),
.B(n_458),
.C(n_459),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_311),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_307),
.B(n_312),
.C(n_313),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_310),
.B(n_464),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_310),
.B(n_486),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

XNOR2x1_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_316),
.Y(n_313)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_346),
.B(n_437),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_343),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_326),
.B(n_343),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_330),
.C(n_332),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_327),
.A2(n_328),
.B1(n_434),
.B2(n_435),
.Y(n_433)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_330),
.B(n_332),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.C(n_339),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_333),
.A2(n_334),
.B1(n_335),
.B2(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_333),
.Y(n_384)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_339),
.B(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_431),
.B(n_436),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_385),
.B(n_430),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_377),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_349),
.B(n_377),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_366),
.C(n_375),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_350),
.A2(n_351),
.B1(n_396),
.B2(n_398),
.Y(n_395)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_361),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_359),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_359),
.C(n_361),
.Y(n_379)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_366),
.A2(n_375),
.B1(n_376),
.B2(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_366),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_370),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_367),
.A2(n_368),
.B1(n_370),
.B2(n_371),
.Y(n_388)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_374),
.Y(n_421)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_382),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_379),
.B(n_380),
.C(n_382),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_399),
.B(n_429),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_395),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_387),
.B(n_395),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.C(n_393),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_412),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_389),
.A2(n_390),
.B1(n_393),
.B2(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_393),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_396),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_400),
.A2(n_414),
.B(n_428),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_411),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_401),
.B(n_411),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_409),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_402),
.B(n_409),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_418),
.B(n_427),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_416),
.B(n_417),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_422),
.Y(n_418)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_433),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_432),
.B(n_433),
.Y(n_436)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

CKINVDCx14_ASAP7_75t_R g440 ( 
.A(n_441),
.Y(n_440)
);

OR2x6_ASAP7_75t_SL g441 ( 
.A(n_442),
.B(n_468),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_442),
.B(n_468),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_444),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_443),
.B(n_445),
.C(n_460),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_460),
.Y(n_444)
);

XNOR2x1_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_446),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_457),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_457),
.C(n_477),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_450),
.B1(n_455),
.B2(n_456),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_455),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_465),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_461),
.B(n_466),
.C(n_467),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_499),
.Y(n_471)
);

INVxp33_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_474),
.B(n_475),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_478),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_480),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_481),
.A2(n_482),
.B1(n_490),
.B2(n_491),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.Y(n_482)
);

XNOR2x1_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_489),
.Y(n_484)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx6_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_497),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);


endmodule