module real_aes_7951_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_552;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_500;
wire n_307;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g286 ( .A(n_0), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g163 ( .A1(n_1), .A2(n_3), .B1(n_164), .B2(n_166), .C(n_170), .Y(n_163) );
AOI21xp33_ASAP7_75t_L g254 ( .A1(n_2), .A2(n_229), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g549 ( .A(n_2), .Y(n_549) );
INVx1_ASAP7_75t_L g212 ( .A(n_4), .Y(n_212) );
AND2x6_ASAP7_75t_L g234 ( .A(n_4), .B(n_210), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_4), .B(n_543), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_5), .A2(n_336), .B(n_337), .Y(n_335) );
INVx1_ASAP7_75t_L g261 ( .A(n_6), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_7), .B(n_328), .Y(n_327) );
AO22x2_ASAP7_75t_L g90 ( .A1(n_8), .A2(n_26), .B1(n_91), .B2(n_92), .Y(n_90) );
INVx1_ASAP7_75t_L g227 ( .A(n_9), .Y(n_227) );
INVx1_ASAP7_75t_L g342 ( .A(n_10), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_11), .B(n_242), .Y(n_315) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_12), .A2(n_27), .B1(n_91), .B2(n_95), .Y(n_94) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_13), .B(n_229), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_14), .B(n_250), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_15), .A2(n_192), .B1(n_193), .B2(n_194), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_15), .Y(n_192) );
AOI221xp5_ASAP7_75t_L g142 ( .A1(n_16), .A2(n_77), .B1(n_143), .B2(n_148), .C(n_152), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g339 ( .A1(n_17), .A2(n_340), .B(n_341), .C(n_343), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_18), .A2(n_81), .B1(n_182), .B2(n_183), .Y(n_80) );
INVx1_ASAP7_75t_L g182 ( .A(n_18), .Y(n_182) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_19), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_20), .B(n_259), .Y(n_288) );
INVx1_ASAP7_75t_L g171 ( .A(n_21), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_22), .Y(n_84) );
INVx1_ASAP7_75t_L g275 ( .A(n_23), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_24), .Y(n_122) );
INVx2_ASAP7_75t_L g232 ( .A(n_25), .Y(n_232) );
OAI221xp5_ASAP7_75t_L g203 ( .A1(n_27), .A2(n_42), .B1(n_50), .B2(n_204), .C(n_205), .Y(n_203) );
INVxp67_ASAP7_75t_L g206 ( .A(n_27), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_28), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_29), .A2(n_81), .B1(n_183), .B2(n_551), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_29), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_L g299 ( .A1(n_30), .A2(n_234), .B(n_237), .C(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g273 ( .A(n_31), .Y(n_273) );
OAI22xp5_ASAP7_75t_SL g185 ( .A1(n_32), .A2(n_54), .B1(n_186), .B2(n_187), .Y(n_185) );
INVx1_ASAP7_75t_L g187 ( .A(n_32), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_33), .B(n_259), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_34), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_35), .Y(n_134) );
CKINVDCx16_ASAP7_75t_R g276 ( .A(n_36), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_37), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_38), .B(n_229), .Y(n_330) );
OAI22xp5_ASAP7_75t_SL g195 ( .A1(n_39), .A2(n_58), .B1(n_196), .B2(n_197), .Y(n_195) );
CKINVDCx16_ASAP7_75t_R g196 ( .A(n_39), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_39), .A2(n_237), .B1(n_269), .B2(n_271), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_40), .Y(n_308) );
CKINVDCx16_ASAP7_75t_R g283 ( .A(n_41), .Y(n_283) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_42), .A2(n_60), .B1(n_91), .B2(n_95), .Y(n_100) );
INVxp67_ASAP7_75t_L g207 ( .A(n_42), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_43), .A2(n_246), .B(n_258), .C(n_260), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_44), .Y(n_318) );
INVx1_ASAP7_75t_L g256 ( .A(n_45), .Y(n_256) );
AOI22xp5_ASAP7_75t_SL g539 ( .A1(n_45), .A2(n_81), .B1(n_183), .B2(n_256), .Y(n_539) );
INVx1_ASAP7_75t_L g210 ( .A(n_46), .Y(n_210) );
INVx1_ASAP7_75t_L g226 ( .A(n_47), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_48), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_49), .B(n_124), .Y(n_123) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_50), .A2(n_66), .B1(n_91), .B2(n_92), .Y(n_98) );
A2O1A1Ixp33_ASAP7_75t_SL g241 ( .A1(n_51), .A2(n_242), .B(n_243), .C(n_246), .Y(n_241) );
INVxp67_ASAP7_75t_L g244 ( .A(n_52), .Y(n_244) );
INVx1_ASAP7_75t_L g177 ( .A(n_53), .Y(n_177) );
INVx1_ASAP7_75t_L g186 ( .A(n_54), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_55), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g279 ( .A(n_56), .Y(n_279) );
INVx1_ASAP7_75t_L g311 ( .A(n_57), .Y(n_311) );
INVx1_ASAP7_75t_L g197 ( .A(n_58), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g312 ( .A1(n_58), .A2(n_234), .B(n_237), .C(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g193 ( .A(n_59), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_61), .B(n_287), .Y(n_301) );
INVx2_ASAP7_75t_L g224 ( .A(n_62), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_63), .B(n_242), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_64), .A2(n_234), .B(n_237), .C(n_285), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_65), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_67), .B(n_263), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_68), .Y(n_291) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_69), .A2(n_234), .B(n_237), .C(n_325), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_70), .Y(n_332) );
INVx1_ASAP7_75t_L g240 ( .A(n_71), .Y(n_240) );
CKINVDCx16_ASAP7_75t_R g338 ( .A(n_72), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_73), .B(n_287), .Y(n_326) );
INVx1_ASAP7_75t_L g91 ( .A(n_74), .Y(n_91) );
INVx1_ASAP7_75t_L g93 ( .A(n_74), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_75), .B(n_222), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_76), .A2(n_229), .B(n_235), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_200), .B1(n_213), .B2(n_537), .C(n_538), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_184), .Y(n_79) );
INVx1_ASAP7_75t_L g183 ( .A(n_81), .Y(n_183) );
AND3x1_ASAP7_75t_L g81 ( .A(n_82), .B(n_142), .C(n_163), .Y(n_81) );
NOR3xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_106), .C(n_128), .Y(n_82) );
OAI22xp5_ASAP7_75t_L g83 ( .A1(n_84), .A2(n_85), .B1(n_101), .B2(n_102), .Y(n_83) );
INVx1_ASAP7_75t_SL g85 ( .A(n_86), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
OR2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_96), .Y(n_87) );
INVx2_ASAP7_75t_L g176 ( .A(n_88), .Y(n_176) );
OR2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_94), .Y(n_88) );
AND2x2_ASAP7_75t_L g105 ( .A(n_89), .B(n_94), .Y(n_105) );
AND2x2_ASAP7_75t_L g147 ( .A(n_89), .B(n_120), .Y(n_147) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
AND2x2_ASAP7_75t_L g110 ( .A(n_90), .B(n_94), .Y(n_110) );
AND2x2_ASAP7_75t_L g121 ( .A(n_90), .B(n_100), .Y(n_121) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g95 ( .A(n_93), .Y(n_95) );
INVx2_ASAP7_75t_L g120 ( .A(n_94), .Y(n_120) );
INVx1_ASAP7_75t_L g162 ( .A(n_94), .Y(n_162) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
NAND2x1p5_ASAP7_75t_L g104 ( .A(n_97), .B(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g146 ( .A(n_97), .B(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_99), .Y(n_97) );
INVx1_ASAP7_75t_L g112 ( .A(n_98), .Y(n_112) );
INVx1_ASAP7_75t_L g119 ( .A(n_98), .Y(n_119) );
INVx1_ASAP7_75t_L g141 ( .A(n_98), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_98), .B(n_100), .Y(n_151) );
AND2x2_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g156 ( .A(n_100), .B(n_141), .Y(n_156) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_105), .B(n_156), .Y(n_155) );
AND2x4_ASAP7_75t_L g181 ( .A(n_105), .B(n_111), .Y(n_181) );
OAI221xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_113), .B1(n_114), .B2(n_122), .C(n_123), .Y(n_106) );
INVx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x6_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g138 ( .A(n_110), .Y(n_138) );
AND2x2_ASAP7_75t_L g165 ( .A(n_111), .B(n_147), .Y(n_165) );
AND2x6_ASAP7_75t_L g175 ( .A(n_111), .B(n_176), .Y(n_175) );
INVx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_121), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
INVx1_ASAP7_75t_L g127 ( .A(n_119), .Y(n_127) );
INVx1_ASAP7_75t_L g133 ( .A(n_120), .Y(n_133) );
AND2x4_ASAP7_75t_L g126 ( .A(n_121), .B(n_127), .Y(n_126) );
NAND2x1p5_ASAP7_75t_L g132 ( .A(n_121), .B(n_133), .Y(n_132) );
BUFx4f_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
BUFx12f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_130), .B1(n_134), .B2(n_135), .Y(n_128) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx4_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g136 ( .A(n_137), .Y(n_136) );
OR2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx4_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g149 ( .A(n_147), .B(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g169 ( .A(n_147), .B(n_156), .Y(n_169) );
BUFx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OR2x6_ASAP7_75t_L g161 ( .A(n_151), .B(n_162), .Y(n_161) );
OAI22xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B1(n_157), .B2(n_158), .Y(n_152) );
BUFx2_ASAP7_75t_R g154 ( .A(n_155), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_159), .Y(n_158) );
BUFx4f_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
INVx6_ASAP7_75t_SL g160 ( .A(n_161), .Y(n_160) );
BUFx2_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B1(n_177), .B2(n_178), .Y(n_170) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx4_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx11_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx6_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_188), .B1(n_189), .B2(n_199), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_185), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_189), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B1(n_195), .B2(n_198), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g194 ( .A(n_193), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_195), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_201), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_202), .Y(n_201) );
AND3x1_ASAP7_75t_SL g202 ( .A(n_203), .B(n_208), .C(n_211), .Y(n_202) );
INVxp67_ASAP7_75t_L g543 ( .A(n_203), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g544 ( .A(n_208), .Y(n_544) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_208), .A2(n_230), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g555 ( .A(n_208), .Y(n_555) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_209), .B(n_212), .Y(n_548) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_SL g554 ( .A(n_211), .B(n_555), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_212), .Y(n_211) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND4x1_ASAP7_75t_L g214 ( .A(n_215), .B(n_455), .C(n_502), .D(n_522), .Y(n_214) );
NOR3xp33_ASAP7_75t_SL g215 ( .A(n_216), .B(n_385), .C(n_410), .Y(n_215) );
OAI211xp5_ASAP7_75t_SL g216 ( .A1(n_217), .A2(n_293), .B(n_345), .C(n_375), .Y(n_216) );
INVxp67_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_219), .B(n_264), .Y(n_218) );
INVx3_ASAP7_75t_SL g427 ( .A(n_219), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_219), .B(n_358), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_219), .B(n_280), .Y(n_508) );
AND2x2_ASAP7_75t_L g531 ( .A(n_219), .B(n_397), .Y(n_531) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_252), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g349 ( .A(n_221), .B(n_253), .Y(n_349) );
INVx3_ASAP7_75t_L g362 ( .A(n_221), .Y(n_362) );
AND2x2_ASAP7_75t_L g367 ( .A(n_221), .B(n_252), .Y(n_367) );
OR2x2_ASAP7_75t_L g418 ( .A(n_221), .B(n_359), .Y(n_418) );
BUFx2_ASAP7_75t_L g438 ( .A(n_221), .Y(n_438) );
AND2x2_ASAP7_75t_L g448 ( .A(n_221), .B(n_359), .Y(n_448) );
AND2x2_ASAP7_75t_L g454 ( .A(n_221), .B(n_265), .Y(n_454) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_228), .B(n_249), .Y(n_221) );
INVx4_ASAP7_75t_L g251 ( .A(n_222), .Y(n_251) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g266 ( .A(n_223), .Y(n_266) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
AND2x2_ASAP7_75t_SL g263 ( .A(n_224), .B(n_225), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
BUFx2_ASAP7_75t_L g336 ( .A(n_229), .Y(n_336) );
AND2x4_ASAP7_75t_L g229 ( .A(n_230), .B(n_234), .Y(n_229) );
NAND2x1p5_ASAP7_75t_L g277 ( .A(n_230), .B(n_234), .Y(n_277) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g238 ( .A(n_232), .Y(n_238) );
INVx1_ASAP7_75t_L g270 ( .A(n_232), .Y(n_270) );
INVx1_ASAP7_75t_L g239 ( .A(n_233), .Y(n_239) );
INVx1_ASAP7_75t_L g242 ( .A(n_233), .Y(n_242) );
INVx3_ASAP7_75t_L g245 ( .A(n_233), .Y(n_245) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_233), .Y(n_259) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_233), .Y(n_272) );
INVx4_ASAP7_75t_SL g248 ( .A(n_234), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_240), .B(n_241), .C(n_248), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_236), .A2(n_248), .B(n_256), .C(n_257), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g337 ( .A1(n_236), .A2(n_248), .B(n_338), .C(n_339), .Y(n_337) );
INVx5_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x6_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_238), .Y(n_247) );
BUFx3_ASAP7_75t_L g305 ( .A(n_238), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_245), .B(n_261), .Y(n_260) );
INVx5_ASAP7_75t_L g287 ( .A(n_245), .Y(n_287) );
INVx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_247), .Y(n_329) );
OAI22xp33_ASAP7_75t_L g267 ( .A1(n_248), .A2(n_268), .B1(n_276), .B2(n_277), .Y(n_267) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_250), .A2(n_254), .B(n_262), .Y(n_253) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_SL g307 ( .A(n_251), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_253), .B(n_359), .Y(n_373) );
INVx2_ASAP7_75t_L g383 ( .A(n_253), .Y(n_383) );
AND2x2_ASAP7_75t_L g396 ( .A(n_253), .B(n_362), .Y(n_396) );
OR2x2_ASAP7_75t_L g407 ( .A(n_253), .B(n_359), .Y(n_407) );
AND2x2_ASAP7_75t_SL g453 ( .A(n_253), .B(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g465 ( .A(n_253), .Y(n_465) );
AND2x2_ASAP7_75t_L g511 ( .A(n_253), .B(n_265), .Y(n_511) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx4_ASAP7_75t_L g328 ( .A(n_259), .Y(n_328) );
INVx1_ASAP7_75t_L g292 ( .A(n_263), .Y(n_292) );
INVx2_ASAP7_75t_L g322 ( .A(n_263), .Y(n_322) );
OA21x2_ASAP7_75t_L g334 ( .A1(n_263), .A2(n_335), .B(n_344), .Y(n_334) );
INVx3_ASAP7_75t_SL g384 ( .A(n_264), .Y(n_384) );
OR2x2_ASAP7_75t_L g437 ( .A(n_264), .B(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_280), .Y(n_264) );
INVx3_ASAP7_75t_L g359 ( .A(n_265), .Y(n_359) );
AND2x2_ASAP7_75t_L g426 ( .A(n_265), .B(n_281), .Y(n_426) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_265), .Y(n_494) );
AOI33xp33_ASAP7_75t_L g498 ( .A1(n_265), .A2(n_427), .A3(n_434), .B1(n_443), .B2(n_499), .B3(n_500), .Y(n_498) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .B(n_278), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_266), .B(n_279), .Y(n_278) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_266), .A2(n_282), .B(n_290), .Y(n_281) );
INVx2_ASAP7_75t_L g306 ( .A(n_266), .Y(n_306) );
INVx2_ASAP7_75t_L g289 ( .A(n_269), .Y(n_289) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OAI22xp5_ASAP7_75t_SL g271 ( .A1(n_272), .A2(n_273), .B1(n_274), .B2(n_275), .Y(n_271) );
INVx2_ASAP7_75t_L g274 ( .A(n_272), .Y(n_274) );
INVx4_ASAP7_75t_L g340 ( .A(n_272), .Y(n_340) );
OAI21xp5_ASAP7_75t_L g282 ( .A1(n_277), .A2(n_283), .B(n_284), .Y(n_282) );
OAI21xp5_ASAP7_75t_L g310 ( .A1(n_277), .A2(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_L g347 ( .A(n_280), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_280), .B(n_362), .Y(n_361) );
NOR3xp33_ASAP7_75t_L g421 ( .A(n_280), .B(n_422), .C(n_424), .Y(n_421) );
AND2x2_ASAP7_75t_L g447 ( .A(n_280), .B(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_280), .B(n_454), .Y(n_457) );
AND2x2_ASAP7_75t_L g510 ( .A(n_280), .B(n_511), .Y(n_510) );
INVx3_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx3_ASAP7_75t_L g366 ( .A(n_281), .Y(n_366) );
OR2x2_ASAP7_75t_L g460 ( .A(n_281), .B(n_359), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_288), .C(n_289), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_292), .B(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_292), .B(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_319), .Y(n_293) );
AOI32xp33_ASAP7_75t_L g411 ( .A1(n_294), .A2(n_412), .A3(n_414), .B1(n_416), .B2(n_419), .Y(n_411) );
NOR2xp67_ASAP7_75t_L g484 ( .A(n_294), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g514 ( .A(n_294), .Y(n_514) );
INVx4_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g446 ( .A(n_295), .B(n_430), .Y(n_446) );
AND2x2_ASAP7_75t_L g466 ( .A(n_295), .B(n_392), .Y(n_466) );
AND2x2_ASAP7_75t_L g534 ( .A(n_295), .B(n_452), .Y(n_534) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_309), .Y(n_295) );
INVx3_ASAP7_75t_L g355 ( .A(n_296), .Y(n_355) );
AND2x2_ASAP7_75t_L g369 ( .A(n_296), .B(n_353), .Y(n_369) );
OR2x2_ASAP7_75t_L g374 ( .A(n_296), .B(n_352), .Y(n_374) );
INVx1_ASAP7_75t_L g381 ( .A(n_296), .Y(n_381) );
AND2x2_ASAP7_75t_L g389 ( .A(n_296), .B(n_363), .Y(n_389) );
AND2x2_ASAP7_75t_L g391 ( .A(n_296), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_296), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g444 ( .A(n_296), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_296), .B(n_529), .Y(n_528) );
OR2x6_ASAP7_75t_L g296 ( .A(n_297), .B(n_307), .Y(n_296) );
AOI21xp5_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_299), .B(n_306), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B(n_303), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_303), .A2(n_314), .B(n_315), .Y(n_313) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g343 ( .A(n_305), .Y(n_343) );
INVx1_ASAP7_75t_L g316 ( .A(n_306), .Y(n_316) );
INVx2_ASAP7_75t_L g353 ( .A(n_309), .Y(n_353) );
AND2x2_ASAP7_75t_L g399 ( .A(n_309), .B(n_320), .Y(n_399) );
AND2x2_ASAP7_75t_L g409 ( .A(n_309), .B(n_334), .Y(n_409) );
AO21x2_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_316), .B(n_317), .Y(n_309) );
INVx2_ASAP7_75t_L g529 ( .A(n_319), .Y(n_529) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_333), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_320), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g370 ( .A(n_320), .Y(n_370) );
AND2x2_ASAP7_75t_L g414 ( .A(n_320), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g430 ( .A(n_320), .B(n_393), .Y(n_430) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g378 ( .A(n_321), .Y(n_378) );
AND2x2_ASAP7_75t_L g392 ( .A(n_321), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g443 ( .A(n_321), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_321), .B(n_353), .Y(n_475) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_323), .B(n_331), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_330), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B(n_329), .Y(n_325) );
AND2x2_ASAP7_75t_L g354 ( .A(n_333), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g415 ( .A(n_333), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_333), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g452 ( .A(n_333), .Y(n_452) );
INVx1_ASAP7_75t_L g485 ( .A(n_333), .Y(n_485) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g363 ( .A(n_334), .B(n_353), .Y(n_363) );
INVx1_ASAP7_75t_L g393 ( .A(n_334), .Y(n_393) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_336), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_340), .B(n_342), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_350), .B1(n_356), .B2(n_363), .C(n_364), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_347), .B(n_367), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_347), .B(n_430), .Y(n_507) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_349), .B(n_397), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_349), .B(n_358), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_349), .B(n_372), .Y(n_501) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_354), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g423 ( .A(n_353), .Y(n_423) );
AND2x2_ASAP7_75t_L g398 ( .A(n_354), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g476 ( .A(n_354), .Y(n_476) );
AND2x2_ASAP7_75t_L g408 ( .A(n_355), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_355), .B(n_378), .Y(n_424) );
AND2x2_ASAP7_75t_L g488 ( .A(n_355), .B(n_414), .Y(n_488) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g397 ( .A(n_359), .B(n_366), .Y(n_397) );
AND2x2_ASAP7_75t_L g493 ( .A(n_360), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_362), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_363), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_363), .B(n_370), .Y(n_458) );
AND2x2_ASAP7_75t_L g478 ( .A(n_363), .B(n_378), .Y(n_478) );
AND2x2_ASAP7_75t_L g499 ( .A(n_363), .B(n_443), .Y(n_499) );
OAI32xp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_368), .A3(n_370), .B1(n_371), .B2(n_374), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_SL g372 ( .A(n_366), .Y(n_372) );
NAND2x1_ASAP7_75t_L g413 ( .A(n_366), .B(n_396), .Y(n_413) );
OR2x2_ASAP7_75t_L g417 ( .A(n_366), .B(n_418), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_366), .B(n_465), .Y(n_518) );
INVx1_ASAP7_75t_L g386 ( .A(n_367), .Y(n_386) );
OAI221xp5_ASAP7_75t_SL g504 ( .A1(n_368), .A2(n_459), .B1(n_505), .B2(n_508), .C(n_509), .Y(n_504) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g376 ( .A(n_369), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g419 ( .A(n_369), .B(n_392), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_369), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g497 ( .A(n_369), .B(n_430), .Y(n_497) );
INVxp67_ASAP7_75t_L g433 ( .A(n_370), .Y(n_433) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
AND2x2_ASAP7_75t_L g503 ( .A(n_372), .B(n_490), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_372), .B(n_453), .Y(n_526) );
INVx1_ASAP7_75t_L g401 ( .A(n_374), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_374), .B(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g519 ( .A(n_374), .B(n_520), .Y(n_519) );
OAI21xp5_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_379), .B(n_382), .Y(n_375) );
AND2x2_ASAP7_75t_L g388 ( .A(n_377), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g472 ( .A(n_381), .B(n_392), .Y(n_472) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
AND2x2_ASAP7_75t_L g490 ( .A(n_383), .B(n_448), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_383), .B(n_447), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_384), .B(n_396), .Y(n_470) );
OAI211xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B(n_390), .C(n_400), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_386), .A2(n_421), .B1(n_425), .B2(n_428), .C(n_431), .Y(n_420) );
AOI31xp33_ASAP7_75t_L g515 ( .A1(n_386), .A2(n_516), .A3(n_517), .B(n_519), .Y(n_515) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_394), .B1(n_396), .B2(n_398), .Y(n_390) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g516 ( .A(n_396), .Y(n_516) );
INVx1_ASAP7_75t_L g479 ( .A(n_397), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_399), .A2(n_523), .B(n_525), .C(n_527), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_404), .B2(n_408), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_405), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI221xp5_ASAP7_75t_SL g495 ( .A1(n_407), .A2(n_441), .B1(n_460), .B2(n_496), .C(n_498), .Y(n_495) );
INVx1_ASAP7_75t_L g491 ( .A(n_408), .Y(n_491) );
INVx1_ASAP7_75t_L g445 ( .A(n_409), .Y(n_445) );
NAND3xp33_ASAP7_75t_SL g410 ( .A(n_411), .B(n_420), .C(n_435), .Y(n_410) );
OAI21xp33_ASAP7_75t_L g461 ( .A1(n_412), .A2(n_462), .B(n_466), .Y(n_461) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_414), .B(n_514), .Y(n_513) );
INVxp67_ASAP7_75t_L g521 ( .A(n_415), .Y(n_521) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g459 ( .A(n_422), .B(n_442), .Y(n_459) );
INVx1_ASAP7_75t_L g434 ( .A(n_423), .Y(n_434) );
AND2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_L g432 ( .A(n_426), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_426), .B(n_464), .Y(n_463) );
NOR4xp25_ASAP7_75t_L g431 ( .A(n_427), .B(n_432), .C(n_433), .D(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI222xp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_440), .B1(n_446), .B2(n_447), .C1(n_449), .C2(n_453), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_437), .B(n_439), .Y(n_436) );
INVx1_ASAP7_75t_L g533 ( .A(n_437), .Y(n_533) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_445), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_449), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI21xp5_ASAP7_75t_SL g509 ( .A1(n_454), .A2(n_510), .B(n_512), .Y(n_509) );
NOR4xp25_ASAP7_75t_L g455 ( .A(n_456), .B(n_467), .C(n_480), .D(n_495), .Y(n_455) );
OAI221xp5_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_458), .B1(n_459), .B2(n_460), .C(n_461), .Y(n_456) );
INVx1_ASAP7_75t_L g536 ( .A(n_457), .Y(n_536) );
INVx1_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_464), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
OAI222xp33_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_471), .B1(n_473), .B2(n_474), .C1(n_477), .C2(n_479), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AOI211xp5_ASAP7_75t_L g502 ( .A1(n_472), .A2(n_503), .B(n_504), .C(n_515), .Y(n_502) );
OR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
OAI222xp33_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_486), .B1(n_487), .B2(n_489), .C1(n_491), .C2(n_492), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVxp67_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_497), .A2(n_500), .B1(n_533), .B2(n_534), .Y(n_532) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OAI211xp5_ASAP7_75t_SL g527 ( .A1(n_528), .A2(n_530), .B(n_532), .C(n_535), .Y(n_527) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OAI322xp33_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .A3(n_544), .B1(n_545), .B2(n_549), .C1(n_550), .C2(n_552), .Y(n_538) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_546), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_547), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_553), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_554), .Y(n_553) );
endmodule