module fake_jpeg_29130_n_333 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_333);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_6),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_44),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_47),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_54),
.Y(n_91)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_57),
.Y(n_70)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_63),
.Y(n_88)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_66),
.A2(n_75),
.B1(n_95),
.B2(n_63),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_69),
.B(n_101),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_45),
.A2(n_65),
.B1(n_51),
.B2(n_60),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_102),
.B1(n_104),
.B2(n_108),
.Y(n_121)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_28),
.B(n_22),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_84),
.B(n_109),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_35),
.B1(n_23),
.B2(n_28),
.Y(n_86)
);

AO22x1_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_63),
.B1(n_54),
.B2(n_27),
.Y(n_120)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_61),
.A2(n_30),
.B1(n_21),
.B2(n_37),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_46),
.B(n_26),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_45),
.A2(n_30),
.B1(n_19),
.B2(n_37),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_57),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_107),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_51),
.A2(n_35),
.B1(n_23),
.B2(n_41),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_57),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_59),
.A2(n_60),
.B1(n_65),
.B2(n_58),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_47),
.B(n_19),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_73),
.A2(n_23),
.B(n_35),
.C(n_36),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_111),
.B(n_99),
.Y(n_168)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_127),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_81),
.Y(n_122)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_81),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_138),
.Y(n_164)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_130),
.B1(n_131),
.B2(n_135),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_63),
.B(n_54),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_32),
.B1(n_25),
.B2(n_24),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_73),
.A2(n_32),
.B1(n_36),
.B2(n_41),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_80),
.A2(n_40),
.B1(n_29),
.B2(n_41),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_143),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_40),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_133),
.B(n_134),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_0),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_86),
.A2(n_57),
.B1(n_1),
.B2(n_2),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_77),
.A2(n_57),
.B1(n_2),
.B2(n_3),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_79),
.B(n_0),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_70),
.A2(n_96),
.B1(n_78),
.B2(n_68),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_86),
.B(n_0),
.C(n_3),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_131),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_98),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_72),
.A2(n_4),
.B(n_5),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_70),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_99),
.Y(n_158)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_124),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_152),
.B(n_179),
.Y(n_209)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_158),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_166),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_116),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_177),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_168),
.B(n_171),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_82),
.B1(n_87),
.B2(n_76),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_128),
.B1(n_117),
.B2(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_170),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_130),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g172 ( 
.A(n_120),
.B(n_85),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_129),
.C(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_147),
.B1(n_141),
.B2(n_12),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_114),
.B(n_100),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_114),
.B(n_87),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_180),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_121),
.A2(n_71),
.B1(n_9),
.B2(n_10),
.Y(n_179)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_113),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_182),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_183),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_172),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_132),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_187),
.B(n_198),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_76),
.B1(n_67),
.B2(n_111),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_188),
.A2(n_194),
.B1(n_199),
.B2(n_201),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_146),
.C(n_115),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_193),
.B(n_200),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_153),
.A2(n_146),
.B1(n_67),
.B2(n_123),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_161),
.A2(n_118),
.B(n_110),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_164),
.B(n_162),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_112),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_153),
.A2(n_123),
.B1(n_118),
.B2(n_71),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_110),
.C(n_147),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_179),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_205),
.A2(n_207),
.B1(n_210),
.B2(n_214),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_156),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_165),
.A2(n_13),
.B1(n_15),
.B2(n_113),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_161),
.B(n_113),
.C(n_13),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_211),
.B(n_176),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_161),
.A2(n_15),
.B1(n_154),
.B2(n_163),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_175),
.B(n_163),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_165),
.A2(n_156),
.B1(n_172),
.B2(n_154),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_198),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_215),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_216),
.A2(n_229),
.B1(n_230),
.B2(n_233),
.Y(n_255)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_219),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_226),
.B(n_230),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_213),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_227),
.Y(n_250)
);

OAI32xp33_ASAP7_75t_L g228 ( 
.A1(n_192),
.A2(n_150),
.A3(n_148),
.B1(n_160),
.B2(n_149),
.Y(n_228)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_149),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_191),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_236),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_185),
.B(n_151),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_235),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_151),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_190),
.B(n_200),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_238),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_199),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_240),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_241),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_209),
.B1(n_214),
.B2(n_210),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_244),
.A2(n_216),
.B1(n_229),
.B2(n_225),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_233),
.A2(n_187),
.B1(n_188),
.B2(n_186),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_246),
.A2(n_255),
.B1(n_209),
.B2(n_263),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_190),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_259),
.C(n_239),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_222),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_258),
.B(n_217),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_183),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_272),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_231),
.Y(n_265)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_266),
.A2(n_268),
.B1(n_272),
.B2(n_280),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_256),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_270),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_209),
.B1(n_218),
.B2(n_220),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_231),
.Y(n_269)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_269),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_219),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_275),
.B1(n_279),
.B2(n_247),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_246),
.A2(n_220),
.B1(n_215),
.B2(n_205),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_274),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_245),
.A2(n_207),
.B1(n_212),
.B2(n_211),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_242),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_224),
.C(n_223),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_260),
.C(n_243),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_248),
.Y(n_278)
);

NOR3xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_250),
.C(n_227),
.Y(n_285)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_242),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_249),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_195),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_266),
.Y(n_298)
);

BUFx12_ASAP7_75t_L g283 ( 
.A(n_277),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_271),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_289),
.C(n_262),
.Y(n_303)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_244),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_268),
.A2(n_260),
.B(n_247),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_290),
.A2(n_280),
.B(n_228),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_264),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_293),
.A2(n_262),
.B1(n_250),
.B2(n_254),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_297),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_300),
.B(n_305),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_288),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_301),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_261),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_303),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_257),
.Y(n_304)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_304),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_196),
.Y(n_305)
);

AOI321xp33_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_286),
.A3(n_294),
.B1(n_284),
.B2(n_289),
.C(n_291),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_301),
.B(n_302),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_295),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_310),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_287),
.C(n_282),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_282),
.B(n_261),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_313),
.A2(n_213),
.B(n_184),
.Y(n_318)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_315),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_SL g316 ( 
.A1(n_311),
.A2(n_254),
.B(n_249),
.C(n_221),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_318),
.B(n_321),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_236),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_320),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_306),
.A2(n_314),
.B1(n_309),
.B2(n_232),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_189),
.B(n_197),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_317),
.B(n_148),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_323),
.A2(n_324),
.B(n_157),
.Y(n_329)
);

NAND4xp25_ASAP7_75t_SL g325 ( 
.A(n_316),
.B(n_182),
.C(n_166),
.D(n_174),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_324),
.C(n_181),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_159),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_327),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_328),
.C(n_329),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_331),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_326),
.Y(n_333)
);


endmodule