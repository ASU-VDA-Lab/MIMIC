module fake_jpeg_5131_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_40),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_8),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_42),
.Y(n_53)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_29),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_45),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_33),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_17),
.B1(n_26),
.B2(n_27),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_48),
.B1(n_37),
.B2(n_23),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_17),
.B1(n_26),
.B2(n_30),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_50),
.B(n_14),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_17),
.B1(n_42),
.B2(n_35),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_19),
.B1(n_20),
.B2(n_30),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_19),
.B1(n_20),
.B2(n_18),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_18),
.B1(n_34),
.B2(n_21),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_44),
.C(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_23),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_67),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_68),
.Y(n_91)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_75),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_51),
.B1(n_54),
.B2(n_49),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_83),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_69),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_76),
.B(n_81),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_77),
.A2(n_79),
.B(n_84),
.Y(n_120)
);

OR2x4_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_23),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_23),
.B1(n_28),
.B2(n_16),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_90),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_36),
.C(n_38),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_89),
.C(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_16),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_96),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_67),
.A2(n_36),
.B(n_43),
.Y(n_89)
);

OR2x2_ASAP7_75t_SL g90 ( 
.A(n_52),
.B(n_62),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_61),
.A2(n_28),
.B1(n_16),
.B2(n_14),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_68),
.B1(n_56),
.B2(n_15),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_62),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_52),
.A2(n_38),
.B(n_16),
.C(n_45),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_61),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_95),
.B1(n_76),
.B2(n_81),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_115),
.B(n_128),
.C(n_98),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_123),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_108),
.B(n_121),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_65),
.B1(n_59),
.B2(n_64),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_72),
.B1(n_78),
.B2(n_83),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_53),
.C(n_49),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_71),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_111),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_71),
.Y(n_111)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_119),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_89),
.A2(n_48),
.B1(n_47),
.B2(n_64),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_78),
.B(n_43),
.Y(n_150)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_53),
.C(n_68),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_69),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_68),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_127),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_56),
.B1(n_33),
.B2(n_32),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_100),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_130),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_99),
.B(n_90),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_131),
.B(n_45),
.Y(n_192)
);

AOI22x1_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_132),
.A2(n_122),
.B1(n_119),
.B2(n_113),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx6p67_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_144),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_92),
.B(n_91),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_143),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_142),
.B1(n_147),
.B2(n_126),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_117),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_141),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_63),
.B1(n_56),
.B2(n_75),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_73),
.Y(n_144)
);

NAND2x1_ASAP7_75t_SL g145 ( 
.A(n_106),
.B(n_91),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_145),
.A2(n_150),
.B(n_45),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_146),
.A2(n_105),
.B1(n_127),
.B2(n_122),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_91),
.B(n_75),
.C(n_72),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_149),
.Y(n_174)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_110),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_151),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_111),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_154),
.Y(n_187)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_97),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_157),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_74),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_24),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_158),
.B(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_2),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_3),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_161),
.A2(n_147),
.B1(n_142),
.B2(n_133),
.Y(n_201)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_180),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_102),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_163),
.B(n_175),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_101),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_165),
.A2(n_171),
.B(n_178),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_120),
.C(n_114),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_170),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_114),
.C(n_105),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_172),
.A2(n_189),
.B1(n_146),
.B2(n_137),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_139),
.B1(n_154),
.B2(n_150),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_173),
.A2(n_134),
.B1(n_32),
.B2(n_22),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_38),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_176),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_177),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_43),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_181),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_149),
.B(n_109),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_184),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_3),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_155),
.B(n_13),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_186),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_188),
.A2(n_192),
.B(n_129),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_140),
.A2(n_142),
.B1(n_135),
.B2(n_147),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_116),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_190),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_3),
.Y(n_191)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_191),
.Y(n_197)
);

NAND2x1p5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_145),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_194),
.A2(n_199),
.B(n_204),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_174),
.B(n_148),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_196),
.B(n_200),
.Y(n_228)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_172),
.A2(n_142),
.B1(n_145),
.B2(n_152),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_203),
.A2(n_218),
.B(n_205),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_164),
.A2(n_135),
.B(n_129),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_160),
.B(n_151),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_209),
.Y(n_226)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_219),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_193),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_212),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_178),
.A2(n_140),
.B1(n_159),
.B2(n_137),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_215),
.A2(n_220),
.B1(n_203),
.B2(n_201),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_216),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_217),
.A2(n_165),
.B1(n_189),
.B2(n_170),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_168),
.A2(n_141),
.B(n_130),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_178),
.A2(n_122),
.B1(n_158),
.B2(n_134),
.Y(n_220)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_223),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_163),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_225),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_168),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_175),
.C(n_169),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_229),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_192),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_184),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_231),
.B(n_233),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_232),
.A2(n_200),
.B1(n_198),
.B2(n_220),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_219),
.C(n_181),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_211),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_236),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_212),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_194),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_238),
.B(n_247),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_215),
.A2(n_165),
.B1(n_160),
.B2(n_185),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_240),
.A2(n_217),
.B1(n_209),
.B2(n_205),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_194),
.B(n_179),
.C(n_185),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_244),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_193),
.C(n_183),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_182),
.C(n_166),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_246),
.B(n_214),
.Y(n_259)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_208),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_248),
.B(n_214),
.Y(n_254)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_243),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_250),
.Y(n_282)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

XOR2x2_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_195),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_259),
.B(n_265),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_229),
.B(n_204),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_239),
.Y(n_274)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_258),
.A2(n_261),
.B1(n_266),
.B2(n_267),
.Y(n_271)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_263),
.B(n_264),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_230),
.Y(n_264)
);

A2O1A1O1Ixp25_ASAP7_75t_L g265 ( 
.A1(n_246),
.A2(n_222),
.B(n_196),
.C(n_207),
.D(n_197),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_232),
.A2(n_207),
.B1(n_176),
.B2(n_197),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_234),
.A2(n_202),
.B1(n_191),
.B2(n_166),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_227),
.B1(n_240),
.B2(n_233),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_223),
.B(n_202),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_239),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_262),
.A2(n_244),
.B1(n_226),
.B2(n_241),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_268),
.B1(n_253),
.B2(n_270),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_275),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_224),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_255),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_279),
.C(n_283),
.Y(n_289)
);

A2O1A1O1Ixp25_ASAP7_75t_L g278 ( 
.A1(n_252),
.A2(n_225),
.B(n_231),
.C(n_228),
.D(n_242),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_278),
.B(n_287),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_134),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_237),
.Y(n_280)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

O2A1O1Ixp33_ASAP7_75t_SL g281 ( 
.A1(n_257),
.A2(n_116),
.B(n_22),
.C(n_6),
.Y(n_281)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_38),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_116),
.C(n_38),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_269),
.C(n_266),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_265),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_288),
.A2(n_292),
.B(n_293),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_290),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_269),
.C(n_255),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_251),
.C(n_22),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_294),
.A2(n_295),
.B(n_298),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_45),
.C(n_28),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_284),
.A2(n_276),
.B1(n_282),
.B2(n_285),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_297),
.B(n_278),
.Y(n_308)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_273),
.A2(n_45),
.B(n_10),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_271),
.A2(n_10),
.B(n_13),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_300),
.B(n_295),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_274),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_305),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_275),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_289),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_281),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_294),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_296),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_313),
.C(n_289),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_302),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_11),
.B1(n_15),
.B2(n_9),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_312),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_290),
.A2(n_4),
.B(n_5),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_11),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_317),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_304),
.B(n_296),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_318),
.A2(n_321),
.B(n_322),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_323),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_309),
.A2(n_9),
.B(n_10),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_12),
.C(n_13),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_320),
.A2(n_311),
.B1(n_312),
.B2(n_310),
.Y(n_325)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_325),
.Y(n_331)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

NAND3xp33_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_330),
.C(n_7),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_314),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_329),
.A2(n_12),
.B(n_6),
.C(n_7),
.Y(n_332)
);

NOR3xp33_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_12),
.C(n_6),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_332),
.B(n_333),
.Y(n_334)
);

OAI221xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_327),
.B1(n_329),
.B2(n_328),
.C(n_324),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_335),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_331),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_7),
.Y(n_338)
);


endmodule