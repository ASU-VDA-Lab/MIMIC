module real_jpeg_1950_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_215;
wire n_176;
wire n_221;
wire n_249;
wire n_286;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_297;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_97;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_213;
wire n_179;
wire n_295;
wire n_133;
wire n_202;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_1),
.B(n_35),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_1),
.B(n_48),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_1),
.B(n_29),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_1),
.B(n_71),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_1),
.B(n_54),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_2),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_2),
.B(n_58),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_2),
.B(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_2),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_2),
.B(n_54),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_2),
.B(n_35),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_3),
.B(n_58),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_3),
.B(n_26),
.Y(n_275)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_5),
.B(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_5),
.B(n_35),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_5),
.B(n_71),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_5),
.B(n_26),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_6),
.B(n_29),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_6),
.B(n_71),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_6),
.B(n_48),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_6),
.B(n_54),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_6),
.B(n_26),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_6),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_6),
.B(n_58),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_9),
.B(n_26),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_9),
.B(n_58),
.Y(n_65)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_9),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_9),
.B(n_43),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_9),
.B(n_54),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_9),
.B(n_48),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_9),
.B(n_35),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_13),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_13),
.B(n_48),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_13),
.B(n_29),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_14),
.B(n_71),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_14),
.B(n_35),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_14),
.B(n_48),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_14),
.B(n_29),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_165),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_164),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_127),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_20),
.B(n_127),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_83),
.C(n_107),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_21),
.B(n_107),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_62),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_22),
.B(n_63),
.C(n_72),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.C(n_50),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_23),
.A2(n_50),
.B1(n_51),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_23),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_33),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_24)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_26),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_28),
.B(n_32),
.C(n_33),
.Y(n_117)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_29),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_34),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_34),
.B(n_41),
.Y(n_253)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_38),
.B(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.C(n_45),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_39),
.A2(n_45),
.B1(n_46),
.B2(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_39),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_40),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_41),
.B(n_208),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_41),
.B(n_97),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_41),
.B(n_47),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_42),
.B(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_45),
.A2(n_46),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_47),
.B(n_149),
.Y(n_206)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.C(n_60),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_53),
.B1(n_60),
.B2(n_61),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_56),
.B(n_82),
.Y(n_252)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_72),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.C(n_68),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_68),
.A2(n_69),
.B(n_70),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_71),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_78),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_74),
.B(n_77),
.C(n_78),
.Y(n_155)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_76),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.C(n_81),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_81),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_100),
.B1(n_101),
.B2(n_104),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_81),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_81),
.A2(n_102),
.B1(n_133),
.B2(n_134),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_83),
.B(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_98),
.C(n_105),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_84),
.B(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.C(n_91),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_85),
.B(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_87),
.B(n_91),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_113),
.Y(n_202)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_90),
.B(n_112),
.C(n_114),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.C(n_95),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_92),
.B(n_95),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_94),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_94),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_96),
.B(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_98),
.A2(n_99),
.B1(n_105),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_102),
.B(n_133),
.Y(n_176)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_116),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_117),
.C(n_118),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_114),
.B2(n_115),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_112),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_111),
.A2(n_112),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_112),
.B(n_243),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_114),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_124),
.C(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_123),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_124),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_163),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_150),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_144),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_142),
.B2(n_143),
.Y(n_130)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_141),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_162),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_160),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_215),
.Y(n_165)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_191),
.B(n_214),
.Y(n_167)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_168),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_189),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_169),
.B(n_189),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.C(n_186),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_186),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_181),
.C(n_183),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_181),
.B1(n_182),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.C(n_179),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_175),
.A2(n_176),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_192),
.B(n_194),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_209),
.C(n_211),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_195),
.A2(n_196),
.B1(n_209),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_202),
.C(n_203),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_197),
.A2(n_198),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_202),
.B(n_203),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.C(n_207),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_206),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_207),
.B(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_209),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_211),
.B(n_294),
.Y(n_293)
);

NOR3xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_297),
.C(n_298),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_291),
.B(n_296),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_279),
.B(n_290),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_265),
.B(n_278),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_246),
.B(n_264),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_221),
.B(n_229),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.C(n_228),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_222),
.A2(n_223),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_223),
.A2(n_224),
.B(n_225),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_228),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_237),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_238),
.C(n_242),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_235),
.C(n_236),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_234),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_241),
.B1(n_242),
.B2(n_245),
.Y(n_237)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_245),
.A2(n_257),
.B(n_258),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_255),
.B(n_263),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_251),
.B(n_254),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_249),
.B(n_250),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_256),
.B(n_259),
.Y(n_263)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_266),
.B(n_267),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_273),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_272),
.C(n_273),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_276),
.C(n_277),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_280),
.B(n_281),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_286),
.C(n_287),
.Y(n_292)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_292),
.B(n_293),
.Y(n_296)
);


endmodule