module real_aes_16087_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g115 ( .A(n_0), .B(n_116), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_1), .A2(n_4), .B1(n_255), .B2(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_2), .A2(n_40), .B1(n_150), .B2(n_152), .Y(n_149) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_3), .A2(n_22), .B1(n_152), .B2(n_195), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_5), .A2(n_15), .B1(n_177), .B2(n_246), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_6), .A2(n_57), .B1(n_197), .B2(n_222), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_7), .A2(n_16), .B1(n_150), .B2(n_181), .Y(n_611) );
INVx1_ASAP7_75t_L g116 ( .A(n_8), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_9), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_10), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_11), .A2(n_17), .B1(n_179), .B2(n_221), .Y(n_220) );
BUFx2_ASAP7_75t_L g107 ( .A(n_12), .Y(n_107) );
OR2x2_ASAP7_75t_L g123 ( .A(n_12), .B(n_36), .Y(n_123) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_13), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_14), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_18), .A2(n_97), .B1(n_177), .B2(n_255), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_19), .A2(n_37), .B1(n_213), .B2(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_20), .B(n_178), .Y(n_210) );
OAI21x1_ASAP7_75t_L g166 ( .A1(n_21), .A2(n_54), .B(n_167), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_23), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_24), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_25), .B(n_156), .Y(n_519) );
INVx4_ASAP7_75t_R g574 ( .A(n_26), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g157 ( .A1(n_27), .A2(n_44), .B1(n_158), .B2(n_160), .Y(n_157) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_28), .A2(n_50), .B1(n_160), .B2(n_177), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_29), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_30), .B(n_213), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_31), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_32), .B(n_152), .Y(n_526) );
INVx1_ASAP7_75t_L g535 ( .A(n_33), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_SL g592 ( .A1(n_34), .A2(n_150), .B(n_162), .C(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_35), .A2(n_51), .B1(n_150), .B2(n_160), .Y(n_508) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_36), .Y(n_105) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_38), .A2(n_82), .B1(n_150), .B2(n_194), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_39), .A2(n_43), .B1(n_150), .B2(n_181), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_41), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_42), .A2(n_56), .B1(n_177), .B2(n_232), .Y(n_257) );
INVx1_ASAP7_75t_L g523 ( .A(n_45), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_46), .B(n_150), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_47), .Y(n_544) );
INVx2_ASAP7_75t_L g129 ( .A(n_48), .Y(n_129) );
INVx1_ASAP7_75t_L g110 ( .A(n_49), .Y(n_110) );
BUFx3_ASAP7_75t_L g132 ( .A(n_49), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_52), .A2(n_134), .B1(n_840), .B2(n_841), .Y(n_133) );
INVx1_ASAP7_75t_L g840 ( .A(n_52), .Y(n_840) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_53), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_55), .A2(n_84), .B1(n_150), .B2(n_160), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_58), .A2(n_71), .B1(n_158), .B2(n_232), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_59), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_60), .A2(n_73), .B1(n_150), .B2(n_181), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_61), .A2(n_95), .B1(n_177), .B2(n_179), .Y(n_176) );
AND2x4_ASAP7_75t_L g146 ( .A(n_62), .B(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g167 ( .A(n_63), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_64), .Y(n_119) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_65), .A2(n_88), .B1(n_158), .B2(n_160), .Y(n_531) );
AO22x1_ASAP7_75t_L g561 ( .A1(n_66), .A2(n_72), .B1(n_243), .B2(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g147 ( .A(n_67), .Y(n_147) );
AND2x2_ASAP7_75t_L g595 ( .A(n_68), .B(n_164), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_69), .B(n_197), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_70), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_74), .B(n_152), .Y(n_545) );
INVx2_ASAP7_75t_L g156 ( .A(n_75), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_76), .B(n_164), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_77), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_78), .A2(n_96), .B1(n_160), .B2(n_197), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_79), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_80), .B(n_174), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_81), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g854 ( .A(n_83), .Y(n_854) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_85), .A2(n_135), .B1(n_848), .B2(n_849), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_85), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_86), .A2(n_100), .B1(n_102), .B2(n_117), .Y(n_99) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_87), .B(n_164), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_89), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_90), .B(n_164), .Y(n_541) );
INVx1_ASAP7_75t_L g114 ( .A(n_91), .Y(n_114) );
NAND2xp33_ASAP7_75t_L g214 ( .A(n_92), .B(n_178), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g569 ( .A1(n_93), .A2(n_183), .B(n_197), .C(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g576 ( .A(n_94), .B(n_577), .Y(n_576) );
NAND2xp33_ASAP7_75t_L g549 ( .A(n_98), .B(n_159), .Y(n_549) );
HB1xp67_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx8_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OR2x6_ASAP7_75t_L g102 ( .A(n_103), .B(n_108), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
NOR2x1p5_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
AND3x2_ASAP7_75t_L g121 ( .A(n_109), .B(n_113), .C(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_115), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g494 ( .A(n_114), .Y(n_494) );
OR2x6_ASAP7_75t_L g117 ( .A(n_118), .B(n_124), .Y(n_117) );
INVxp67_ASAP7_75t_SL g850 ( .A(n_118), .Y(n_850) );
NOR2x1_ASAP7_75t_R g118 ( .A(n_119), .B(n_120), .Y(n_118) );
INVx3_ASAP7_75t_L g846 ( .A(n_120), .Y(n_846) );
INVx4_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_122), .B(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NOR2x1_ASAP7_75t_L g860 ( .A(n_123), .B(n_132), .Y(n_860) );
OAI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_133), .B(n_842), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
BUFx12f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x6_ASAP7_75t_SL g127 ( .A(n_128), .B(n_130), .Y(n_127) );
BUFx3_ASAP7_75t_L g852 ( .A(n_128), .Y(n_852) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_129), .B(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g841 ( .A(n_134), .Y(n_841) );
OA22x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_491), .B1(n_495), .B2(n_497), .Y(n_134) );
INVx2_ASAP7_75t_L g849 ( .A(n_135), .Y(n_849) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_387), .Y(n_135) );
NOR2x1_ASAP7_75t_L g136 ( .A(n_137), .B(n_339), .Y(n_136) );
NAND3xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_286), .C(n_324), .Y(n_137) );
AOI221xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_217), .B1(n_237), .B2(n_265), .C(n_271), .Y(n_138) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_139), .A2(n_464), .B1(n_467), .B2(n_468), .Y(n_463) );
INVx2_ASAP7_75t_SL g139 ( .A(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_188), .Y(n_140) );
INVx1_ASAP7_75t_L g378 ( .A(n_141), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_170), .Y(n_141) );
INVx1_ASAP7_75t_L g330 ( .A(n_142), .Y(n_330) );
AND2x4_ASAP7_75t_L g373 ( .A(n_142), .B(n_294), .Y(n_373) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g301 ( .A(n_143), .B(n_204), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_143), .B(n_270), .Y(n_361) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g269 ( .A(n_144), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g285 ( .A(n_144), .B(n_190), .Y(n_285) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_144), .Y(n_292) );
INVx1_ASAP7_75t_L g348 ( .A(n_144), .Y(n_348) );
AO31x2_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_148), .A3(n_163), .B(n_168), .Y(n_144) );
INVx2_ASAP7_75t_L g185 ( .A(n_145), .Y(n_185) );
AO31x2_ASAP7_75t_L g218 ( .A1(n_145), .A2(n_172), .A3(n_219), .B(n_225), .Y(n_218) );
AO31x2_ASAP7_75t_L g240 ( .A1(n_145), .A2(n_191), .A3(n_241), .B(n_248), .Y(n_240) );
AO31x2_ASAP7_75t_L g609 ( .A1(n_145), .A2(n_236), .A3(n_610), .B(n_613), .Y(n_609) );
BUFx10_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g200 ( .A(n_146), .Y(n_200) );
BUFx10_ASAP7_75t_L g510 ( .A(n_146), .Y(n_510) );
INVx1_ASAP7_75t_L g565 ( .A(n_146), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_153), .B1(n_157), .B2(n_161), .Y(n_148) );
INVx1_ASAP7_75t_L g179 ( .A(n_150), .Y(n_179) );
INVx4_ASAP7_75t_L g181 ( .A(n_150), .Y(n_181) );
INVx1_ASAP7_75t_L g232 ( .A(n_150), .Y(n_232) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_151), .Y(n_152) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_151), .Y(n_160) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_151), .Y(n_178) );
INVx2_ASAP7_75t_L g195 ( .A(n_151), .Y(n_195) );
INVx1_ASAP7_75t_L g197 ( .A(n_151), .Y(n_197) );
INVx1_ASAP7_75t_L g223 ( .A(n_151), .Y(n_223) );
INVx1_ASAP7_75t_L g244 ( .A(n_151), .Y(n_244) );
INVx1_ASAP7_75t_L g247 ( .A(n_151), .Y(n_247) );
INVx1_ASAP7_75t_L g256 ( .A(n_151), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_152), .B(n_588), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_153), .A2(n_161), .B1(n_231), .B2(n_233), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_153), .A2(n_161), .B1(n_242), .B2(n_245), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_153), .A2(n_161), .B1(n_254), .B2(n_257), .Y(n_253) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g509 ( .A(n_154), .Y(n_509) );
BUFx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g547 ( .A(n_155), .Y(n_547) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx8_ASAP7_75t_L g162 ( .A(n_156), .Y(n_162) );
INVx1_ASAP7_75t_L g183 ( .A(n_156), .Y(n_183) );
INVx1_ASAP7_75t_L g522 ( .A(n_156), .Y(n_522) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g213 ( .A(n_159), .Y(n_213) );
OAI22xp33_ASAP7_75t_L g573 ( .A1(n_159), .A2(n_247), .B1(n_574), .B2(n_575), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_160), .B(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g533 ( .A(n_160), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g175 ( .A1(n_161), .A2(n_176), .B1(n_180), .B2(n_182), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_161), .A2(n_193), .B1(n_196), .B2(n_198), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_161), .A2(n_212), .B(n_214), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_161), .A2(n_182), .B1(n_220), .B2(n_224), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_161), .A2(n_507), .B1(n_508), .B2(n_509), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_161), .A2(n_198), .B1(n_531), .B2(n_532), .Y(n_530) );
OAI22x1_ASAP7_75t_L g610 ( .A1(n_161), .A2(n_198), .B1(n_611), .B2(n_612), .Y(n_610) );
INVx6_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
O2A1O1Ixp5_ASAP7_75t_L g208 ( .A1(n_162), .A2(n_181), .B(n_209), .C(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_162), .A2(n_549), .B(n_550), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_162), .B(n_561), .Y(n_560) );
A2O1A1Ixp33_ASAP7_75t_L g623 ( .A1(n_162), .A2(n_557), .B(n_561), .C(n_564), .Y(n_623) );
AO31x2_ASAP7_75t_L g505 ( .A1(n_163), .A2(n_506), .A3(n_510), .B(n_511), .Y(n_505) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2x1_ASAP7_75t_L g551 ( .A(n_164), .B(n_552), .Y(n_551) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_165), .B(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_165), .B(n_187), .Y(n_186) );
BUFx3_ASAP7_75t_L g191 ( .A(n_165), .Y(n_191) );
INVx2_ASAP7_75t_SL g206 ( .A(n_165), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_165), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g527 ( .A(n_165), .B(n_510), .Y(n_527) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g174 ( .A(n_166), .Y(n_174) );
INVx3_ASAP7_75t_L g268 ( .A(n_170), .Y(n_268) );
AND2x2_ASAP7_75t_L g283 ( .A(n_170), .B(n_204), .Y(n_283) );
INVx2_ASAP7_75t_L g289 ( .A(n_170), .Y(n_289) );
AND2x4_ASAP7_75t_L g351 ( .A(n_170), .B(n_190), .Y(n_351) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_170), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_170), .B(n_484), .Y(n_483) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g300 ( .A(n_171), .B(n_190), .Y(n_300) );
AND2x2_ASAP7_75t_L g328 ( .A(n_171), .B(n_329), .Y(n_328) );
BUFx2_ASAP7_75t_L g407 ( .A(n_171), .Y(n_407) );
AO31x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .A3(n_184), .B(n_186), .Y(n_171) );
AO31x2_ASAP7_75t_L g529 ( .A1(n_172), .A2(n_199), .A3(n_530), .B(n_534), .Y(n_529) );
AOI21x1_ASAP7_75t_L g584 ( .A1(n_172), .A2(n_585), .B(n_595), .Y(n_584) );
BUFx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_173), .B(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_173), .B(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g577 ( .A(n_173), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_173), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g202 ( .A(n_174), .Y(n_202) );
INVx2_ASAP7_75t_L g236 ( .A(n_174), .Y(n_236) );
OAI21xp33_ASAP7_75t_L g564 ( .A1(n_174), .A2(n_559), .B(n_565), .Y(n_564) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVxp67_ASAP7_75t_SL g562 ( .A(n_178), .Y(n_562) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_181), .A2(n_544), .B(n_545), .C(n_546), .Y(n_543) );
INVx1_ASAP7_75t_SL g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g198 ( .A(n_183), .Y(n_198) );
AO31x2_ASAP7_75t_L g252 ( .A1(n_184), .A2(n_228), .A3(n_253), .B(n_258), .Y(n_252) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_185), .A2(n_569), .B(n_572), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_204), .Y(n_188) );
INVx1_ASAP7_75t_L g363 ( .A(n_189), .Y(n_363) );
NAND2x1_ASAP7_75t_L g391 ( .A(n_189), .B(n_283), .Y(n_391) );
BUFx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OR2x2_ASAP7_75t_L g293 ( .A(n_190), .B(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g329 ( .A(n_190), .Y(n_329) );
INVx1_ASAP7_75t_L g405 ( .A(n_190), .Y(n_405) );
AO31x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .A3(n_199), .B(n_201), .Y(n_190) );
INVx2_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_195), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_198), .B(n_573), .Y(n_572) );
AO31x2_ASAP7_75t_L g227 ( .A1(n_199), .A2(n_228), .A3(n_230), .B(n_234), .Y(n_227) );
INVx2_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_SL g215 ( .A(n_200), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
NOR2xp33_ASAP7_75t_SL g225 ( .A(n_202), .B(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g229 ( .A(n_202), .Y(n_229) );
AND2x4_ASAP7_75t_L g344 ( .A(n_204), .B(n_329), .Y(n_344) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
BUFx2_ASAP7_75t_L g366 ( .A(n_205), .Y(n_366) );
OAI21x1_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_216), .Y(n_205) );
OAI21x1_ASAP7_75t_L g270 ( .A1(n_206), .A2(n_207), .B(n_216), .Y(n_270) );
OAI21x1_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_211), .B(n_215), .Y(n_207) );
AND2x4_ASAP7_75t_L g238 ( .A(n_217), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_227), .Y(n_217) );
INVx4_ASAP7_75t_SL g262 ( .A(n_218), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_218), .B(n_264), .Y(n_274) );
BUFx2_ASAP7_75t_L g338 ( .A(n_218), .Y(n_338) );
AND2x2_ASAP7_75t_L g382 ( .A(n_218), .B(n_240), .Y(n_382) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_223), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g260 ( .A(n_227), .Y(n_260) );
OR2x2_ASAP7_75t_L g298 ( .A(n_227), .B(n_240), .Y(n_298) );
INVx2_ASAP7_75t_L g309 ( .A(n_227), .Y(n_309) );
AND2x4_ASAP7_75t_L g312 ( .A(n_227), .B(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_227), .Y(n_353) );
INVx1_ASAP7_75t_L g394 ( .A(n_227), .Y(n_394) );
AO21x2_ASAP7_75t_L g567 ( .A1(n_228), .A2(n_568), .B(n_576), .Y(n_567) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_236), .B(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_250), .Y(n_237) );
INVx2_ASAP7_75t_L g487 ( .A(n_238), .Y(n_487) );
AND2x4_ASAP7_75t_L g448 ( .A(n_239), .B(n_251), .Y(n_448) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g264 ( .A(n_240), .Y(n_264) );
INVx2_ASAP7_75t_L g313 ( .A(n_240), .Y(n_313) );
INVx1_ASAP7_75t_L g369 ( .A(n_240), .Y(n_369) );
AND2x2_ASAP7_75t_L g395 ( .A(n_240), .B(n_320), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_240), .B(n_308), .Y(n_399) );
OAI21xp33_ASAP7_75t_SL g518 ( .A1(n_243), .A2(n_519), .B(n_520), .Y(n_518) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_261), .Y(n_250) );
INVx3_ASAP7_75t_L g376 ( .A(n_251), .Y(n_376) );
AND2x4_ASAP7_75t_L g251 ( .A(n_252), .B(n_260), .Y(n_251) );
INVx2_ASAP7_75t_L g280 ( .A(n_252), .Y(n_280) );
INVx2_ASAP7_75t_L g320 ( .A(n_252), .Y(n_320) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_256), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_260), .B(n_262), .Y(n_321) );
AND2x2_ASAP7_75t_L g349 ( .A(n_260), .B(n_320), .Y(n_349) );
INVx1_ASAP7_75t_L g275 ( .A(n_261), .Y(n_275) );
NAND2x1_ASAP7_75t_L g411 ( .A(n_261), .B(n_385), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_261), .B(n_349), .Y(n_460) );
AND2x4_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g278 ( .A(n_262), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_262), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g368 ( .A(n_262), .B(n_369), .Y(n_368) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_262), .Y(n_445) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_265), .A2(n_458), .B1(n_459), .B2(n_461), .Y(n_457) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_267), .B(n_301), .Y(n_336) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x4_ASAP7_75t_L g359 ( .A(n_268), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g458 ( .A(n_268), .B(n_269), .Y(n_458) );
AND2x2_ASAP7_75t_L g331 ( .A(n_269), .B(n_300), .Y(n_331) );
AND2x4_ASAP7_75t_L g350 ( .A(n_269), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g401 ( .A(n_269), .B(n_328), .Y(n_401) );
INVx1_ASAP7_75t_L g294 ( .A(n_270), .Y(n_294) );
AOI31xp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_275), .A3(n_276), .B(n_281), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_273), .B(n_316), .Y(n_315) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_273), .Y(n_467) );
OAI21xp33_ASAP7_75t_L g485 ( .A1(n_273), .A2(n_275), .B(n_305), .Y(n_485) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g327 ( .A(n_274), .Y(n_327) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g462 ( .A(n_277), .B(n_298), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx2_ASAP7_75t_L g296 ( .A(n_278), .Y(n_296) );
INVx1_ASAP7_75t_L g317 ( .A(n_279), .Y(n_317) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_279), .Y(n_424) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g306 ( .A(n_280), .Y(n_306) );
OR2x2_ASAP7_75t_L g334 ( .A(n_280), .B(n_309), .Y(n_334) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NOR2x1p5_ASAP7_75t_L g323 ( .A(n_285), .B(n_289), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_295), .B1(n_299), .B2(n_302), .C(n_314), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2x1_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g403 ( .A(n_292), .B(n_306), .Y(n_403) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
OR2x2_ASAP7_75t_L g333 ( .A(n_296), .B(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g420 ( .A(n_296), .B(n_312), .Y(n_420) );
AND2x4_ASAP7_75t_L g337 ( .A(n_297), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g356 ( .A(n_298), .B(n_319), .Y(n_356) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AND2x4_ASAP7_75t_SL g372 ( .A(n_300), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g413 ( .A(n_300), .Y(n_413) );
INVx2_ASAP7_75t_L g422 ( .A(n_300), .Y(n_422) );
AND2x2_ASAP7_75t_L g436 ( .A(n_300), .B(n_366), .Y(n_436) );
INVx1_ASAP7_75t_L g414 ( .A(n_301), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_310), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_307), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_304), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2x1p5_ASAP7_75t_L g346 ( .A(n_305), .B(n_312), .Y(n_346) );
AND2x2_ASAP7_75t_L g367 ( .A(n_305), .B(n_368), .Y(n_367) );
NAND2x1_ASAP7_75t_L g475 ( .A(n_305), .B(n_337), .Y(n_475) );
INVx3_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_318), .B(n_322), .Y(n_314) );
NAND2x1_ASAP7_75t_L g476 ( .A(n_316), .B(n_420), .Y(n_476) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_317), .B(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx4_ASAP7_75t_L g385 ( .A(n_319), .Y(n_385) );
AND2x2_ASAP7_75t_L g455 ( .A(n_319), .B(n_360), .Y(n_455) );
INVx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g352 ( .A(n_320), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g365 ( .A(n_323), .B(n_366), .Y(n_365) );
NOR2x1_ASAP7_75t_L g435 ( .A(n_323), .B(n_436), .Y(n_435) );
AOI322xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_328), .A3(n_330), .B1(n_331), .B2(n_332), .C1(n_335), .C2(n_337), .Y(n_324) );
INVxp67_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g418 ( .A(n_328), .B(n_366), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_328), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g442 ( .A(n_328), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g447 ( .A(n_328), .B(n_432), .Y(n_447) );
INVx1_ASAP7_75t_L g456 ( .A(n_328), .Y(n_456) );
OR2x2_ASAP7_75t_L g342 ( .A(n_330), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g469 ( .A(n_330), .Y(n_469) );
AND2x2_ASAP7_75t_L g472 ( .A(n_331), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NOR3xp33_ASAP7_75t_L g408 ( .A(n_334), .B(n_348), .C(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g450 ( .A(n_334), .Y(n_450) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND3xp33_ASAP7_75t_SL g339 ( .A(n_340), .B(n_354), .C(n_364), .Y(n_339) );
AOI222xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_345), .B1(n_347), .B2(n_349), .C1(n_350), .C2(n_352), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OAI22x1_ASAP7_75t_L g486 ( .A1(n_343), .A2(n_487), .B1(n_488), .B2(n_489), .Y(n_486) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g347 ( .A(n_344), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_344), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g440 ( .A(n_344), .B(n_406), .Y(n_440) );
AND2x4_ASAP7_75t_L g470 ( .A(n_344), .B(n_407), .Y(n_470) );
AND2x2_ASAP7_75t_L g451 ( .A(n_345), .B(n_418), .Y(n_451) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g443 ( .A(n_348), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_349), .B(n_382), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_349), .B(n_368), .Y(n_466) );
INVx1_ASAP7_75t_L g386 ( .A(n_350), .Y(n_386) );
INVx2_ASAP7_75t_L g430 ( .A(n_352), .Y(n_430) );
INVx1_ASAP7_75t_L g380 ( .A(n_353), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2x1p5_ASAP7_75t_L g358 ( .A(n_359), .B(n_362), .Y(n_358) );
AOI221xp5_ASAP7_75t_SL g446 ( .A1(n_359), .A2(n_447), .B1(n_448), .B2(n_449), .C(n_451), .Y(n_446) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g432 ( .A(n_361), .Y(n_432) );
INVxp67_ASAP7_75t_SL g484 ( .A(n_361), .Y(n_484) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_363), .B(n_469), .Y(n_478) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_367), .B1(n_370), .B2(n_381), .C(n_383), .Y(n_364) );
OR2x2_ASAP7_75t_L g421 ( .A(n_366), .B(n_422), .Y(n_421) );
AOI32xp33_ASAP7_75t_L g402 ( .A1(n_368), .A2(n_382), .A3(n_403), .B1(n_404), .B2(n_408), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_368), .B(n_424), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_374), .B1(n_377), .B2(n_379), .Y(n_370) );
INVx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_373), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g444 ( .A(n_376), .B(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g437 ( .A(n_380), .B(n_382), .Y(n_437) );
AND2x2_ASAP7_75t_L g490 ( .A(n_380), .B(n_395), .Y(n_490) );
AND2x2_ASAP7_75t_L g449 ( .A(n_381), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_382), .B(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
NOR2x1_ASAP7_75t_L g387 ( .A(n_388), .B(n_452), .Y(n_387) );
NAND4xp75_ASAP7_75t_L g388 ( .A(n_389), .B(n_415), .C(n_433), .D(n_446), .Y(n_388) );
AOI211x1_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B(n_396), .C(n_410), .Y(n_389) );
INVxp67_ASAP7_75t_L g488 ( .A(n_390), .Y(n_488) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OAI21xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_400), .B(n_402), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
BUFx2_ASAP7_75t_L g409 ( .A(n_405), .Y(n_409) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g481 ( .A(n_409), .Y(n_481) );
NOR3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .C(n_414), .Y(n_410) );
INVx2_ASAP7_75t_L g473 ( .A(n_411), .Y(n_473) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NOR2x1_ASAP7_75t_L g415 ( .A(n_416), .B(n_425), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_419), .B1(n_421), .B2(n_423), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B1(n_430), .B2(n_431), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_437), .B(n_438), .Y(n_433) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI21xp33_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_441), .B(n_444), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_445), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g465 ( .A(n_448), .Y(n_465) );
NAND4xp75_ASAP7_75t_SL g452 ( .A(n_453), .B(n_463), .C(n_471), .D(n_479), .Y(n_452) );
OA21x2_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_456), .B(n_457), .Y(n_453) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
NOR2xp67_ASAP7_75t_SL g471 ( .A(n_472), .B(n_474), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_477), .Y(n_474) );
INVxp67_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
AOI21x1_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_485), .B(n_486), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx8_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx12f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_494), .Y(n_493) );
BUFx8_ASAP7_75t_SL g496 ( .A(n_494), .Y(n_496) );
AND2x2_ASAP7_75t_L g859 ( .A(n_494), .B(n_860), .Y(n_859) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_L g497 ( .A(n_498), .B(n_730), .Y(n_497) );
NOR4xp25_ASAP7_75t_L g498 ( .A(n_499), .B(n_630), .C(n_672), .D(n_704), .Y(n_498) );
OAI211xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_536), .B(n_578), .C(n_615), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_513), .Y(n_502) );
INVx2_ASAP7_75t_L g643 ( .A(n_503), .Y(n_643) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g722 ( .A(n_504), .B(n_515), .Y(n_722) );
BUFx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_505), .B(n_529), .Y(n_581) );
AND2x2_ASAP7_75t_L g604 ( .A(n_505), .B(n_605), .Y(n_604) );
INVx2_ASAP7_75t_SL g629 ( .A(n_505), .Y(n_629) );
OR2x2_ASAP7_75t_L g692 ( .A(n_505), .B(n_529), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_509), .A2(n_525), .B(n_526), .Y(n_524) );
OAI21x1_ASAP7_75t_L g557 ( .A1(n_509), .A2(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g552 ( .A(n_510), .Y(n_552) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g626 ( .A(n_514), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g638 ( .A(n_514), .Y(n_638) );
INVxp67_ASAP7_75t_SL g816 ( .A(n_514), .Y(n_816) );
OR2x2_ASAP7_75t_L g829 ( .A(n_514), .B(n_830), .Y(n_829) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_528), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_515), .B(n_583), .Y(n_582) );
INVx3_ASAP7_75t_L g602 ( .A(n_515), .Y(n_602) );
AND2x2_ASAP7_75t_L g649 ( .A(n_515), .B(n_650), .Y(n_649) );
NAND2x1p5_ASAP7_75t_SL g668 ( .A(n_515), .B(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_515), .B(n_603), .Y(n_718) );
INVx1_ASAP7_75t_L g807 ( .A(n_515), .Y(n_807) );
AND2x2_ASAP7_75t_L g836 ( .A(n_515), .B(n_529), .Y(n_836) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_524), .B(n_527), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
BUFx4f_ASAP7_75t_L g591 ( .A(n_522), .Y(n_591) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g603 ( .A(n_529), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_529), .B(n_629), .Y(n_651) );
INVx1_ASAP7_75t_L g671 ( .A(n_529), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_529), .B(n_605), .Y(n_723) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_553), .Y(n_537) );
OR2x2_ASAP7_75t_L g620 ( .A(n_538), .B(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g727 ( .A(n_538), .B(n_676), .Y(n_727) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g636 ( .A(n_539), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_539), .B(n_656), .Y(n_655) );
NOR2x1_ASAP7_75t_L g741 ( .A(n_539), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g599 ( .A(n_540), .Y(n_599) );
BUFx3_ASAP7_75t_L g647 ( .A(n_540), .Y(n_647) );
AND2x2_ASAP7_75t_L g683 ( .A(n_540), .B(n_664), .Y(n_683) );
AND2x2_ASAP7_75t_L g763 ( .A(n_540), .B(n_609), .Y(n_763) );
AND2x2_ASAP7_75t_L g776 ( .A(n_540), .B(n_567), .Y(n_776) );
NAND2x1p5_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
OAI21x1_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_548), .B(n_551), .Y(n_542) );
INVx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g716 ( .A(n_553), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_553), .B(n_646), .Y(n_724) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_566), .Y(n_553) );
AND2x2_ASAP7_75t_L g635 ( .A(n_554), .B(n_567), .Y(n_635) );
INVx1_ASAP7_75t_L g743 ( .A(n_554), .Y(n_743) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x4_ASAP7_75t_L g597 ( .A(n_555), .B(n_567), .Y(n_597) );
AND2x2_ASAP7_75t_L g660 ( .A(n_555), .B(n_566), .Y(n_660) );
AOI21x1_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_560), .B(n_563), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_565), .A2(n_586), .B(n_592), .Y(n_585) );
AND2x2_ASAP7_75t_L g618 ( .A(n_566), .B(n_609), .Y(n_618) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g608 ( .A(n_567), .B(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g676 ( .A(n_567), .B(n_609), .Y(n_676) );
INVx1_ASAP7_75t_L g687 ( .A(n_567), .Y(n_687) );
AND2x2_ASAP7_75t_L g750 ( .A(n_567), .B(n_599), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_596), .B1(n_600), .B2(n_606), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_579), .A2(n_649), .B1(n_652), .B2(n_654), .Y(n_648) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
OR2x2_ASAP7_75t_L g728 ( .A(n_581), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g834 ( .A(n_581), .Y(n_834) );
INVx1_ASAP7_75t_L g693 ( .A(n_582), .Y(n_693) );
OR2x2_ASAP7_75t_L g756 ( .A(n_582), .B(n_651), .Y(n_756) );
OR2x2_ASAP7_75t_L g627 ( .A(n_583), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_583), .B(n_602), .Y(n_703) );
AND2x2_ASAP7_75t_L g720 ( .A(n_583), .B(n_647), .Y(n_720) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_583), .Y(n_737) );
INVxp67_ASAP7_75t_L g785 ( .A(n_583), .Y(n_785) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g605 ( .A(n_584), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_589), .B(n_591), .Y(n_586) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_597), .Y(n_695) );
INVx3_ASAP7_75t_L g700 ( .A(n_597), .Y(n_700) );
AND2x2_ASAP7_75t_L g713 ( .A(n_597), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g813 ( .A(n_597), .B(n_775), .Y(n_813) );
INVx1_ASAP7_75t_L g607 ( .A(n_598), .Y(n_607) );
OR2x2_ASAP7_75t_L g790 ( .A(n_598), .B(n_765), .Y(n_790) );
BUFx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g714 ( .A(n_599), .B(n_624), .Y(n_714) );
AND2x2_ASAP7_75t_L g735 ( .A(n_599), .B(n_660), .Y(n_735) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_604), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_601), .B(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g736 ( .A(n_601), .Y(n_736) );
AND2x2_ASAP7_75t_L g778 ( .A(n_601), .B(n_779), .Y(n_778) );
AND2x4_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx2_ASAP7_75t_L g679 ( .A(n_602), .Y(n_679) );
AND2x2_ASAP7_75t_L g710 ( .A(n_602), .B(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_602), .B(n_669), .Y(n_729) );
AND2x2_ASAP7_75t_L g678 ( .A(n_604), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g794 ( .A(n_604), .Y(n_794) );
AND2x2_ASAP7_75t_L g817 ( .A(n_604), .B(n_807), .Y(n_817) );
INVx1_ASAP7_75t_L g830 ( .A(n_604), .Y(n_830) );
INVx2_ASAP7_75t_L g669 ( .A(n_605), .Y(n_669) );
OR2x2_ASAP7_75t_L g765 ( .A(n_605), .B(n_629), .Y(n_765) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_608), .B(n_646), .Y(n_653) );
INVx2_ASAP7_75t_L g624 ( .A(n_609), .Y(n_624) );
INVx2_ASAP7_75t_L g664 ( .A(n_609), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_609), .B(n_622), .Y(n_686) );
OAI21xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_619), .B(n_625), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_618), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g759 ( .A(n_621), .B(n_760), .Y(n_759) );
OR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
INVx2_ASAP7_75t_L g665 ( .A(n_622), .Y(n_665) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g656 ( .A(n_624), .Y(n_656) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g639 ( .A(n_627), .Y(n_639) );
INVxp67_ASAP7_75t_L g810 ( .A(n_627), .Y(n_810) );
OR2x2_ASAP7_75t_L g712 ( .A(n_628), .B(n_669), .Y(n_712) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND4xp25_ASAP7_75t_L g630 ( .A(n_631), .B(n_640), .C(n_648), .D(n_657), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_637), .C(n_639), .Y(n_631) );
INVx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_L g826 ( .A1(n_633), .A2(n_827), .B(n_829), .C(n_831), .Y(n_826) );
OR2x6_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_635), .B(n_683), .Y(n_682) );
NOR3xp33_ASAP7_75t_L g738 ( .A(n_635), .B(n_739), .C(n_741), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_635), .B(n_714), .Y(n_819) );
AOI221xp5_ASAP7_75t_L g831 ( .A1(n_635), .A2(n_740), .B1(n_832), .B2(n_835), .C(n_837), .Y(n_831) );
INVx1_ASAP7_75t_L g822 ( .A(n_636), .Y(n_822) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_644), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g757 ( .A1(n_641), .A2(n_649), .B1(n_684), .B2(n_758), .C(n_761), .Y(n_757) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_643), .B(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g708 ( .A(n_644), .Y(n_708) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2x1p5_ASAP7_75t_L g662 ( .A(n_646), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g823 ( .A(n_646), .B(n_674), .Y(n_823) );
INVx3_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
BUFx2_ASAP7_75t_L g659 ( .A(n_647), .Y(n_659) );
AND3x1_ASAP7_75t_L g832 ( .A(n_647), .B(n_833), .C(n_834), .Y(n_832) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g702 ( .A(n_651), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g772 ( .A(n_654), .Y(n_772) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g748 ( .A(n_656), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g775 ( .A(n_656), .Y(n_775) );
OAI21xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_661), .B(n_666), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NAND2x1_ASAP7_75t_L g673 ( .A(n_659), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g740 ( .A(n_660), .Y(n_740) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g696 ( .A(n_664), .Y(n_696) );
OR2x2_ASAP7_75t_L g675 ( .A(n_665), .B(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g788 ( .A(n_665), .Y(n_788) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_667), .B(n_815), .Y(n_814) );
OR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
OR2x2_ASAP7_75t_L g744 ( .A(n_668), .B(n_692), .Y(n_744) );
INVx2_ASAP7_75t_L g833 ( .A(n_668), .Y(n_833) );
INVx1_ASAP7_75t_L g707 ( .A(n_669), .Y(n_707) );
NOR4xp25_ASAP7_75t_L g837 ( .A(n_669), .B(n_700), .C(n_838), .D(n_839), .Y(n_837) );
INVx1_ASAP7_75t_L g839 ( .A(n_670), .Y(n_839) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
BUFx3_ASAP7_75t_L g825 ( .A(n_671), .Y(n_825) );
OAI211xp5_ASAP7_75t_SL g672 ( .A1(n_673), .A2(n_677), .B(n_680), .C(n_688), .Y(n_672) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g812 ( .A(n_675), .Y(n_812) );
INVx2_ASAP7_75t_L g797 ( .A(n_676), .Y(n_797) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g680 ( .A1(n_678), .A2(n_681), .B(n_684), .Y(n_680) );
OR2x2_ASAP7_75t_L g764 ( .A(n_679), .B(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g782 ( .A(n_679), .B(n_783), .Y(n_782) );
INVxp67_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g698 ( .A(n_683), .Y(n_698) );
AND2x4_ASAP7_75t_SL g787 ( .A(n_683), .B(n_788), .Y(n_787) );
INVx3_ASAP7_75t_R g684 ( .A(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_686), .Y(n_753) );
INVx1_ASAP7_75t_L g760 ( .A(n_687), .Y(n_760) );
AOI32xp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_694), .A3(n_696), .B1(n_697), .B2(n_701), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_691), .B(n_707), .Y(n_706) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_691), .Y(n_752) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g769 ( .A(n_692), .B(n_707), .Y(n_769) );
INVx2_ASAP7_75t_L g783 ( .A(n_692), .Y(n_783) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g762 ( .A(n_700), .B(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI211xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_708), .B(n_709), .C(n_725), .Y(n_704) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_713), .B(n_715), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g766 ( .A(n_714), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_714), .B(n_801), .Y(n_800) );
OAI32xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .A3(n_719), .B1(n_721), .B2(n_724), .Y(n_715) );
INVx1_ASAP7_75t_L g801 ( .A(n_716), .Y(n_801) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OR2x2_ASAP7_75t_L g793 ( .A(n_718), .B(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVxp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
NOR2x1_ASAP7_75t_L g730 ( .A(n_731), .B(n_802), .Y(n_730) );
NAND4xp25_ASAP7_75t_L g731 ( .A(n_732), .B(n_757), .C(n_770), .D(n_798), .Y(n_731) );
NOR2xp67_ASAP7_75t_L g732 ( .A(n_733), .B(n_745), .Y(n_732) );
OAI32xp33_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_736), .A3(n_737), .B1(n_738), .B2(n_744), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
OR2x2_ASAP7_75t_L g784 ( .A(n_736), .B(n_785), .Y(n_784) );
OAI32xp33_ASAP7_75t_L g789 ( .A1(n_736), .A2(n_790), .A3(n_791), .B1(n_793), .B2(n_795), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_737), .B(n_825), .Y(n_824) );
NAND2xp5_ASAP7_75t_SL g803 ( .A(n_739), .B(n_804), .Y(n_803) );
INVx3_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g796 ( .A(n_742), .B(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g828 ( .A(n_742), .Y(n_828) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g792 ( .A(n_743), .Y(n_792) );
OAI22x1_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_751), .B1(n_753), .B2(n_754), .Y(n_745) );
INVx2_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_755), .B(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx3_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NOR2x1_ASAP7_75t_L g821 ( .A(n_759), .B(n_822), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_764), .B1(n_766), .B2(n_767), .Y(n_761) );
NAND2x1_ASAP7_75t_L g827 ( .A(n_763), .B(n_828), .Y(n_827) );
INVx2_ASAP7_75t_L g838 ( .A(n_763), .Y(n_838) );
INVx2_ASAP7_75t_L g779 ( .A(n_765), .Y(n_779) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NOR3xp33_ASAP7_75t_SL g770 ( .A(n_771), .B(n_780), .C(n_789), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .B(n_777), .Y(n_771) );
NAND2xp33_ASAP7_75t_L g799 ( .A(n_773), .B(n_800), .Y(n_799) );
INVx2_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AND2x4_ASAP7_75t_L g835 ( .A(n_779), .B(n_836), .Y(n_835) );
AOI21xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_784), .B(n_786), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
AND2x4_ASAP7_75t_L g806 ( .A(n_783), .B(n_807), .Y(n_806) );
INVxp67_ASAP7_75t_SL g805 ( .A(n_785), .Y(n_805) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVxp67_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NAND3xp33_ASAP7_75t_SL g802 ( .A(n_803), .B(n_808), .C(n_820), .Y(n_802) );
AND2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
INVx1_ASAP7_75t_L g811 ( .A(n_807), .Y(n_811) );
AOI222xp33_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_812), .B1(n_813), .B2(n_814), .C1(n_817), .C2(n_818), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
O2A1O1Ixp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_823), .B(n_824), .C(n_826), .Y(n_820) );
AOI21xp5_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_851), .B(n_853), .Y(n_842) );
OAI21xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_847), .B(n_850), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_854), .B(n_855), .Y(n_853) );
INVx6_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
BUFx10_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
endmodule