module fake_jpeg_27844_n_57 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_57);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_57;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_2),
.Y(n_11)
);

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_17),
.Y(n_22)
);

OR2x2_ASAP7_75t_SL g17 ( 
.A(n_8),
.B(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_19),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_17),
.B(n_8),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_11),
.B1(n_16),
.B2(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_30),
.Y(n_36)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_15),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_13),
.C(n_15),
.Y(n_37)
);

AO22x1_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_25),
.C(n_10),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_31),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_41),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_13),
.B1(n_32),
.B2(n_14),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_40),
.B1(n_44),
.B2(n_41),
.Y(n_48)
);

XNOR2x1_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_12),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_12),
.C(n_14),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_0),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_40),
.B1(n_43),
.B2(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_45),
.B(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_12),
.B1(n_14),
.B2(n_4),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_48),
.B(n_0),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_45),
.B(n_5),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

AOI322xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_51),
.A3(n_50),
.B1(n_7),
.B2(n_5),
.C1(n_3),
.C2(n_14),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_7),
.Y(n_57)
);


endmodule