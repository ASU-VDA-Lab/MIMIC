module fake_jpeg_31333_n_540 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_540);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_540;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_11),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_16),
.B(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_52),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_53),
.Y(n_151)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_54),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_55),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_57),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_58),
.B(n_89),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_18),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_65),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx2_ASAP7_75t_R g130 ( 
.A(n_70),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_71),
.B(n_76),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_74),
.Y(n_138)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_35),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_79),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_86),
.Y(n_135)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_81),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_25),
.B(n_17),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_38),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_19),
.Y(n_139)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_107),
.B(n_108),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_52),
.B(n_25),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_111),
.B(n_139),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_86),
.A2(n_22),
.B(n_20),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_41),
.C(n_31),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_56),
.A2(n_33),
.B1(n_20),
.B2(n_29),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_136),
.A2(n_33),
.B1(n_41),
.B2(n_82),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_74),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_144),
.B(n_149),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_59),
.B(n_19),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_147),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_59),
.B(n_49),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_91),
.B(n_49),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_91),
.B(n_48),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_157),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_75),
.B(n_48),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_93),
.B(n_50),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_160),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_63),
.B(n_50),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_64),
.B(n_46),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_165),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_67),
.A2(n_36),
.B1(n_34),
.B2(n_29),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_162),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_167),
.B(n_207),
.Y(n_249)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_168),
.Y(n_268)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_170),
.Y(n_245)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_171),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_172),
.Y(n_236)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_173),
.Y(n_238)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_174),
.Y(n_272)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_175),
.Y(n_241)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_176),
.Y(n_253)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_177),
.Y(n_271)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_178),
.Y(n_279)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_179),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_181),
.B(n_182),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_114),
.B(n_33),
.Y(n_182)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

AO21x1_ASAP7_75t_L g228 ( 
.A1(n_185),
.A2(n_219),
.B(n_222),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

BUFx2_ASAP7_75t_SL g260 ( 
.A(n_186),
.Y(n_260)
);

CKINVDCx12_ASAP7_75t_R g189 ( 
.A(n_130),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_189),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_138),
.A2(n_32),
.B1(n_84),
.B2(n_78),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_190),
.A2(n_200),
.B1(n_215),
.B2(n_217),
.Y(n_256)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_192),
.Y(n_251)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_129),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_195),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_114),
.B(n_34),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_216),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_198),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_138),
.A2(n_88),
.B1(n_72),
.B2(n_69),
.Y(n_200)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_134),
.Y(n_201)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_201),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_135),
.B(n_46),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_202),
.B(n_204),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_145),
.B(n_40),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_221),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_118),
.B(n_40),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_151),
.Y(n_205)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_205),
.Y(n_265)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_142),
.Y(n_206)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_206),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_106),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_128),
.B(n_26),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_208),
.B(n_209),
.Y(n_263)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_137),
.Y(n_209)
);

CKINVDCx12_ASAP7_75t_R g210 ( 
.A(n_126),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_210),
.B(n_211),
.Y(n_273)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_124),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_113),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_212),
.B(n_213),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_122),
.B(n_26),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_166),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_104),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_141),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_113),
.Y(n_217)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_218),
.A2(n_224),
.B1(n_227),
.B2(n_131),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_163),
.B(n_26),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_151),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_220),
.A2(n_223),
.B1(n_205),
.B2(n_161),
.Y(n_250)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_124),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_127),
.B(n_34),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_109),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_163),
.B(n_17),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_226),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_141),
.B(n_36),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_125),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_121),
.B1(n_110),
.B2(n_148),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_232),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_197),
.A2(n_136),
.B1(n_121),
.B2(n_156),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_237),
.A2(n_239),
.B1(n_258),
.B2(n_270),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_196),
.A2(n_125),
.B1(n_143),
.B2(n_110),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_193),
.B(n_131),
.C(n_115),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_243),
.B(n_264),
.C(n_140),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_182),
.A2(n_148),
.B1(n_143),
.B2(n_68),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_185),
.A2(n_152),
.B1(n_54),
.B2(n_57),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_199),
.A2(n_152),
.B1(n_53),
.B2(n_55),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_250),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_200),
.A2(n_161),
.B1(n_158),
.B2(n_166),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_187),
.B(n_36),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_177),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_180),
.B(n_155),
.C(n_30),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_184),
.A2(n_30),
.B1(n_29),
.B2(n_155),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_269),
.A2(n_223),
.B1(n_170),
.B2(n_162),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_190),
.A2(n_150),
.B1(n_41),
.B2(n_133),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_183),
.A2(n_150),
.B1(n_41),
.B2(n_133),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_274),
.A2(n_278),
.B1(n_198),
.B2(n_195),
.Y(n_299)
);

A2O1A1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_188),
.A2(n_41),
.B(n_162),
.C(n_133),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_276),
.A2(n_178),
.B(n_214),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_220),
.A2(n_140),
.B1(n_16),
.B2(n_15),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_186),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_280),
.B(n_282),
.Y(n_357)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_281),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_261),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_243),
.B(n_186),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_283),
.B(n_286),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_284),
.B(n_291),
.Y(n_334)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_251),
.Y(n_285)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_285),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_231),
.B(n_206),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_251),
.Y(n_287)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_287),
.Y(n_345)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_249),
.Y(n_288)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_288),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_240),
.B(n_191),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_300),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_230),
.B(n_201),
.Y(n_291)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_292),
.Y(n_342)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_233),
.Y(n_293)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_293),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_228),
.A2(n_212),
.B(n_217),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_294),
.A2(n_2),
.B(n_3),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_252),
.B(n_168),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_295),
.B(n_309),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_228),
.A2(n_227),
.B1(n_224),
.B2(n_218),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_296),
.A2(n_299),
.B1(n_313),
.B2(n_326),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_298),
.Y(n_331)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_238),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_234),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_302),
.B(n_307),
.Y(n_367)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_260),
.Y(n_303)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_303),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_267),
.B(n_176),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_304),
.B(n_306),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_305),
.A2(n_258),
.B1(n_299),
.B2(n_270),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_16),
.Y(n_306)
);

INVx13_ASAP7_75t_L g307 ( 
.A(n_279),
.Y(n_307)
);

INVx13_ASAP7_75t_L g308 ( 
.A(n_279),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_310),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_230),
.B(n_242),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_268),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_242),
.B(n_0),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_311),
.B(n_312),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_253),
.Y(n_312)
);

INVx11_ASAP7_75t_L g313 ( 
.A(n_268),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_252),
.B(n_15),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_315),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_264),
.B(n_2),
.Y(n_315)
);

CKINVDCx12_ASAP7_75t_R g316 ( 
.A(n_266),
.Y(n_316)
);

OAI22x1_ASAP7_75t_L g368 ( 
.A1(n_316),
.A2(n_327),
.B1(n_8),
.B2(n_4),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_317),
.B(n_274),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_275),
.B(n_2),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_318),
.B(n_319),
.Y(n_341)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_238),
.Y(n_319)
);

INVx6_ASAP7_75t_SL g320 ( 
.A(n_248),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_320),
.B(n_321),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_253),
.Y(n_321)
);

AND2x6_ASAP7_75t_L g322 ( 
.A(n_254),
.B(n_140),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_322),
.A2(n_276),
.B(n_254),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_259),
.B(n_10),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_325),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_237),
.B(n_2),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_272),
.Y(n_326)
);

INVx13_ASAP7_75t_L g327 ( 
.A(n_235),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_332),
.A2(n_358),
.B1(n_360),
.B2(n_320),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_301),
.A2(n_256),
.B1(n_246),
.B2(n_269),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_333),
.A2(n_346),
.B1(n_347),
.B2(n_349),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_254),
.C(n_232),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_348),
.C(n_352),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_343),
.Y(n_380)
);

OAI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_288),
.A2(n_235),
.B1(n_255),
.B2(n_247),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_301),
.A2(n_244),
.B1(n_229),
.B2(n_255),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_325),
.A2(n_278),
.B1(n_265),
.B2(n_262),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_309),
.B(n_266),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_315),
.B(n_277),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_354),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_284),
.B(n_311),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_291),
.A2(n_265),
.B1(n_241),
.B2(n_277),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_347),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_289),
.A2(n_241),
.B1(n_236),
.B2(n_233),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_297),
.A2(n_294),
.B1(n_289),
.B2(n_323),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_359),
.A2(n_323),
.B1(n_297),
.B2(n_305),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_295),
.A2(n_236),
.B1(n_245),
.B2(n_272),
.Y(n_360)
);

OAI32xp33_ASAP7_75t_L g362 ( 
.A1(n_322),
.A2(n_248),
.A3(n_245),
.B1(n_234),
.B2(n_10),
.Y(n_362)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_362),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_365),
.A2(n_366),
.B(n_3),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_298),
.A2(n_3),
.B(n_4),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_368),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_339),
.B(n_314),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_369),
.B(n_370),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_339),
.B(n_318),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_371),
.A2(n_378),
.B1(n_3),
.B2(n_4),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_374),
.B(n_375),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_336),
.B(n_287),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_344),
.Y(n_376)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_302),
.Y(n_377)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_377),
.Y(n_411)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_344),
.Y(n_379)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_379),
.Y(n_412)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_330),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_381),
.B(n_384),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_382),
.A2(n_400),
.B(n_351),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_312),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_332),
.A2(n_285),
.B1(n_293),
.B2(n_281),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_385),
.B(n_387),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_340),
.Y(n_386)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_345),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_336),
.B(n_326),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_388),
.B(n_392),
.Y(n_432)
);

CKINVDCx10_ASAP7_75t_R g390 ( 
.A(n_368),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_390),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_353),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_391),
.B(n_307),
.Y(n_425)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_340),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_350),
.B(n_321),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_393),
.B(n_394),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_334),
.B(n_319),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_334),
.B(n_300),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_395),
.B(n_396),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_356),
.B(n_316),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_329),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_397),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_359),
.B(n_356),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_307),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_367),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_341),
.B(n_310),
.Y(n_401)
);

OAI21x1_ASAP7_75t_L g423 ( 
.A1(n_401),
.A2(n_335),
.B(n_328),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_331),
.A2(n_303),
.B(n_313),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_402),
.A2(n_331),
.B(n_367),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_338),
.B(n_327),
.C(n_308),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_348),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_404),
.B(n_406),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_391),
.B(n_354),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_407),
.Y(n_457)
);

A2O1A1Ixp33_ASAP7_75t_SL g408 ( 
.A1(n_402),
.A2(n_365),
.B(n_362),
.C(n_366),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_408),
.A2(n_419),
.B(n_431),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_372),
.A2(n_361),
.B1(n_343),
.B2(n_337),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_409),
.A2(n_417),
.B1(n_420),
.B2(n_374),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_413),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_380),
.A2(n_351),
.B(n_337),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_401),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_372),
.A2(n_363),
.B1(n_341),
.B2(n_342),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_415),
.A2(n_424),
.B1(n_414),
.B2(n_389),
.Y(n_448)
);

OAI22xp33_ASAP7_75t_SL g417 ( 
.A1(n_390),
.A2(n_292),
.B1(n_355),
.B2(n_335),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_400),
.A2(n_335),
.B(n_328),
.Y(n_419)
);

OAI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_399),
.A2(n_400),
.B1(n_378),
.B2(n_385),
.Y(n_420)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_423),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_425),
.B(n_433),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_428),
.A2(n_399),
.B1(n_398),
.B2(n_389),
.Y(n_440)
);

XOR2x2_ASAP7_75t_L g431 ( 
.A(n_380),
.B(n_5),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_383),
.B(n_5),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_383),
.B(n_373),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_434),
.B(n_403),
.C(n_373),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_436),
.B(n_449),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_438),
.A2(n_419),
.B(n_407),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_411),
.B(n_375),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_439),
.B(n_444),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_440),
.A2(n_448),
.B1(n_456),
.B2(n_459),
.Y(n_470)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_405),
.Y(n_441)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_441),
.Y(n_468)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_412),
.Y(n_442)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_388),
.Y(n_443)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_443),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_432),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_432),
.Y(n_445)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_445),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_410),
.B(n_395),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_447),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_410),
.B(n_394),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_424),
.B(n_387),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_450),
.A2(n_451),
.B1(n_453),
.B2(n_455),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_418),
.B(n_392),
.Y(n_451)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_422),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_416),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_430),
.B(n_376),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_458),
.A2(n_460),
.B(n_447),
.Y(n_467)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_426),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_430),
.B(n_379),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_461),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_452),
.B(n_406),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_465),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_437),
.A2(n_413),
.B(n_382),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_464),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_436),
.B(n_434),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_404),
.C(n_425),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_472),
.C(n_475),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_467),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_433),
.C(n_409),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_431),
.C(n_426),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_438),
.B(n_421),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_477),
.B(n_480),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_459),
.A2(n_427),
.B1(n_408),
.B2(n_428),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_478),
.A2(n_470),
.B1(n_461),
.B2(n_457),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_438),
.B(n_453),
.Y(n_480)
);

FAx1_ASAP7_75t_SL g481 ( 
.A(n_443),
.B(n_408),
.CI(n_427),
.CON(n_481),
.SN(n_481)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_481),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_477),
.B(n_474),
.Y(n_486)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_486),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_455),
.Y(n_487)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_487),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_489),
.A2(n_386),
.B1(n_7),
.B2(n_8),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_463),
.B(n_457),
.C(n_435),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_490),
.B(n_463),
.C(n_475),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_435),
.C(n_446),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_491),
.B(n_494),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_468),
.B(n_441),
.Y(n_492)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_492),
.Y(n_509)
);

XOR2x2_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_446),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_408),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_437),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_480),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_495),
.B(n_440),
.Y(n_506)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_469),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_442),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_502),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_484),
.A2(n_473),
.B1(n_471),
.B2(n_476),
.Y(n_502)
);

FAx1_ASAP7_75t_SL g503 ( 
.A(n_490),
.B(n_449),
.CI(n_464),
.CON(n_503),
.SN(n_503)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_506),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_483),
.B(n_466),
.C(n_472),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_504),
.A2(n_505),
.B(n_510),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_483),
.B(n_462),
.C(n_445),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_508),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_495),
.B(n_456),
.C(n_416),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_511),
.B(n_512),
.Y(n_522)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_510),
.Y(n_513)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_513),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_503),
.B(n_498),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_514),
.B(n_518),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_503),
.B(n_485),
.Y(n_518)
);

AOI21x1_ASAP7_75t_SL g519 ( 
.A1(n_511),
.A2(n_488),
.B(n_493),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_519),
.A2(n_482),
.B(n_496),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_501),
.A2(n_482),
.B1(n_488),
.B2(n_494),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_520),
.A2(n_509),
.B(n_512),
.Y(n_528)
);

AOI21xp33_ASAP7_75t_L g523 ( 
.A1(n_517),
.A2(n_499),
.B(n_507),
.Y(n_523)
);

AOI21xp33_ASAP7_75t_L g530 ( 
.A1(n_523),
.A2(n_527),
.B(n_519),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_521),
.A2(n_504),
.B(n_505),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_524),
.B(n_516),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_528),
.B(n_520),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_529),
.B(n_530),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_531),
.B(n_532),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_526),
.B(n_515),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_533),
.A2(n_531),
.B(n_525),
.Y(n_535)
);

BUFx24_ASAP7_75t_SL g536 ( 
.A(n_535),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_500),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_537),
.A2(n_534),
.B1(n_522),
.B2(n_8),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_538),
.B(n_522),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_539),
.A2(n_7),
.B(n_8),
.Y(n_540)
);


endmodule