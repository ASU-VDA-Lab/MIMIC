module real_jpeg_14637_n_12 (n_5, n_4, n_8, n_0, n_306, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_306;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_300;
wire n_221;
wire n_292;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_285;
wire n_45;
wire n_160;
wire n_304;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_205;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_185;
wire n_240;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_295;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_210;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g108 ( 
.A(n_0),
.Y(n_108)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_3),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_3),
.A2(n_42),
.B1(n_46),
.B2(n_113),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_113),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_113),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_35),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_4),
.A2(n_35),
.B1(n_42),
.B2(n_46),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_4),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_7),
.A2(n_42),
.B1(n_46),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_53),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_53),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_7),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_7),
.B(n_58),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_7),
.B(n_45),
.C(n_49),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_7),
.B(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_7),
.B(n_47),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_7),
.A2(n_24),
.B(n_60),
.C(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_7),
.B(n_20),
.Y(n_183)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_30),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_10),
.A2(n_30),
.B1(n_48),
.B2(n_49),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_10),
.A2(n_30),
.B1(n_42),
.B2(n_46),
.Y(n_233)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_93),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_91),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_83),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_15),
.B(n_83),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_69),
.C(n_75),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_16),
.A2(n_17),
.B1(n_69),
.B2(n_77),
.Y(n_301)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_36),
.B1(n_37),
.B2(n_68),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_18),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_25),
.B(n_31),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_19),
.A2(n_73),
.B(n_74),
.Y(n_278)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_20),
.B(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_20),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_20),
.B(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_21),
.B(n_24),
.C(n_53),
.Y(n_198)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_23),
.A2(n_24),
.B1(n_60),
.B2(n_61),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_25),
.A2(n_70),
.B(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_26),
.B(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_31),
.B(n_206),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_32),
.B(n_207),
.Y(n_217)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_54),
.B1(n_55),
.B2(n_67),
.Y(n_37)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_38),
.B(n_77),
.C(n_78),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_38),
.B(n_55),
.C(n_68),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_38),
.A2(n_67),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_38),
.A2(n_67),
.B1(n_78),
.B2(n_295),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_51),
.B(n_52),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_39),
.A2(n_117),
.B(n_233),
.Y(n_264)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_40),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_40),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_40),
.B(n_118),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_47),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_41)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_46),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_42),
.B(n_128),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_46),
.A2(n_53),
.B(n_61),
.Y(n_169)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_47),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_47),
.B(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_47),
.B(n_132),
.Y(n_176)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_49),
.B(n_108),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_49),
.B(n_137),
.Y(n_136)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_51),
.A2(n_164),
.B(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_52),
.Y(n_132)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_63),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_57),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_62),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_62),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_58),
.B(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_58),
.A2(n_63),
.B(n_80),
.Y(n_282)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_66),
.Y(n_82)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_62),
.B(n_86),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_63),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_79),
.B(n_81),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_64),
.B(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_67),
.B(n_204),
.C(n_210),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_69),
.A2(n_77),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_70),
.B(n_217),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_72),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_74),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_75),
.A2(n_76),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_78),
.Y(n_295)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_82),
.B(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_82),
.B(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_90),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_85),
.A2(n_89),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_85),
.B(n_223),
.C(n_229),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_285),
.B(n_302),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_268),
.B(n_284),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_247),
.B(n_267),
.Y(n_95)
);

AOI321xp33_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_213),
.A3(n_240),
.B1(n_245),
.B2(n_246),
.C(n_306),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_190),
.B(n_212),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_172),
.B(n_189),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_155),
.B(n_171),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_133),
.B(n_154),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_125),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_125),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_114),
.B1(n_115),
.B2(n_124),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_104),
.B(n_151),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_111),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_106),
.A2(n_108),
.B(n_111),
.Y(n_167)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_112),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_108),
.A2(n_151),
.B(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_144),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_111),
.A2(n_200),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_117),
.B(n_131),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_119),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_122),
.C(n_124),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_126),
.A2(n_127),
.B1(n_129),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_147),
.B(n_153),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_141),
.B(n_146),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_143),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_145),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_143),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_150),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_157),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_165),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_163),
.C(n_165),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_162),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_164),
.B(n_176),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_170),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_166),
.A2(n_167),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_166),
.A2(n_167),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_168),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_167),
.B(n_264),
.Y(n_275)
);

AOI21xp33_ASAP7_75t_L g289 ( 
.A1(n_167),
.A2(n_275),
.B(n_277),
.Y(n_289)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_188),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_188),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_180),
.B1(n_181),
.B2(n_187),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_175),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_178),
.C(n_180),
.Y(n_191)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_181),
.B(n_195),
.C(n_202),
.Y(n_244)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.CI(n_184),
.CON(n_181),
.SN(n_181)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_192),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_202),
.B2(n_203),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_199),
.B2(n_201),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_201),
.Y(n_220)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_199),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_234),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_234),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_221),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_222),
.C(n_230),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.C(n_220),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_218),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_220),
.B(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_230),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_227),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_226),
.Y(n_238)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_228),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_232),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.C(n_239),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_236),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_239),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_244),
.Y(n_245)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_249),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_266),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_262),
.B2(n_263),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_263),
.C(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_255),
.C(n_260),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_260),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_264),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_270),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_273),
.C(n_280),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_279),
.B2(n_280),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B(n_283),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_282),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_283),
.A2(n_291),
.B1(n_292),
.B2(n_296),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_283),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_289),
.C(n_291),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_297),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_288),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_299),
.Y(n_304)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);


endmodule