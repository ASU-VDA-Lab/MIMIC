module real_aes_13983_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_755, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_755;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_656;
wire n_316;
wire n_153;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_598;
wire n_404;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_266;
wire n_183;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
INVx2_ASAP7_75t_SL g246 ( .A(n_0), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_1), .Y(n_178) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_2), .A2(n_38), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g192 ( .A(n_2), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_3), .B(n_131), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_4), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g138 ( .A(n_5), .B(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_6), .B(n_283), .Y(n_282) );
BUFx3_ASAP7_75t_L g541 ( .A(n_7), .Y(n_541) );
INVx3_ASAP7_75t_L g528 ( .A(n_8), .Y(n_528) );
INVx2_ASAP7_75t_L g537 ( .A(n_9), .Y(n_537) );
INVx1_ASAP7_75t_L g595 ( .A(n_9), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_10), .A2(n_719), .B1(n_720), .B2(n_721), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_10), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_11), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g96 ( .A(n_12), .Y(n_96) );
BUFx3_ASAP7_75t_L g119 ( .A(n_12), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_13), .B(n_165), .Y(n_164) );
BUFx10_ASAP7_75t_L g733 ( .A(n_14), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_15), .A2(n_711), .B1(n_712), .B2(n_713), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_15), .Y(n_712) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_16), .Y(n_215) );
NAND3xp33_ASAP7_75t_L g264 ( .A(n_17), .B(n_174), .C(n_262), .Y(n_264) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_17), .Y(n_740) );
INVx1_ASAP7_75t_L g612 ( .A(n_18), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_18), .A2(n_51), .B1(n_690), .B2(n_691), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_19), .B(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g624 ( .A(n_20), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g649 ( .A(n_20), .B(n_25), .Y(n_649) );
INVxp33_ASAP7_75t_L g682 ( .A(n_20), .Y(n_682) );
INVx1_ASAP7_75t_L g696 ( .A(n_20), .Y(n_696) );
INVx1_ASAP7_75t_L g87 ( .A(n_21), .Y(n_87) );
INVx2_ASAP7_75t_L g631 ( .A(n_22), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_23), .B(n_240), .Y(n_239) );
AOI221xp5_ASAP7_75t_L g574 ( .A1(n_24), .A2(n_70), .B1(n_575), .B2(n_577), .C(n_581), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_24), .A2(n_31), .B1(n_621), .B2(n_632), .Y(n_620) );
INVx2_ASAP7_75t_L g625 ( .A(n_25), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_25), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_26), .B(n_225), .Y(n_224) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_27), .A2(n_31), .B1(n_586), .B2(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g670 ( .A(n_27), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_28), .B(n_182), .Y(n_181) );
AOI221xp5_ASAP7_75t_L g553 ( .A1(n_29), .A2(n_55), .B1(n_554), .B2(n_560), .C(n_563), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_29), .A2(n_55), .B1(n_638), .B2(n_642), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_30), .A2(n_49), .B1(n_567), .B2(n_571), .Y(n_566) );
INVx1_ASAP7_75t_L g667 ( .A(n_30), .Y(n_667) );
AND2x4_ASAP7_75t_L g86 ( .A(n_32), .B(n_87), .Y(n_86) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_32), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_33), .B(n_165), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_34), .B(n_111), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_35), .B(n_165), .Y(n_278) );
INVx1_ASAP7_75t_L g607 ( .A(n_36), .Y(n_607) );
OAI22xp33_ASAP7_75t_SL g650 ( .A1(n_36), .A2(n_65), .B1(n_651), .B2(n_656), .Y(n_650) );
INVx1_ASAP7_75t_L g538 ( .A(n_37), .Y(n_538) );
INVx1_ASAP7_75t_L g559 ( .A(n_37), .Y(n_559) );
INVx1_ASAP7_75t_L g193 ( .A(n_38), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_39), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_40), .A2(n_130), .B(n_244), .C(n_247), .Y(n_243) );
INVx1_ASAP7_75t_L g113 ( .A(n_41), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_42), .B(n_165), .Y(n_186) );
INVx3_ASAP7_75t_L g212 ( .A(n_43), .Y(n_212) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_44), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_45), .B(n_208), .Y(n_287) );
INVx1_ASAP7_75t_L g152 ( .A(n_46), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_47), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_48), .B(n_176), .Y(n_257) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_48), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_49), .A2(n_70), .B1(n_672), .B2(n_675), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_50), .B(n_174), .Y(n_173) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_50), .Y(n_716) );
INVx1_ASAP7_75t_L g544 ( .A(n_51), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_52), .B(n_230), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_53), .Y(n_615) );
XNOR2xp5_ASAP7_75t_L g522 ( .A(n_54), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g238 ( .A(n_56), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_57), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_58), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_59), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g91 ( .A(n_60), .Y(n_91) );
INVx1_ASAP7_75t_L g136 ( .A(n_60), .Y(n_136) );
BUFx3_ASAP7_75t_L g149 ( .A(n_60), .Y(n_149) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_61), .A2(n_65), .B1(n_591), .B2(n_598), .Y(n_590) );
INVx1_ASAP7_75t_L g688 ( .A(n_61), .Y(n_688) );
INVx1_ASAP7_75t_L g711 ( .A(n_62), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_63), .B(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g210 ( .A(n_64), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_66), .Y(n_603) );
INVx2_ASAP7_75t_L g629 ( .A(n_67), .Y(n_629) );
AND2x2_ASAP7_75t_L g641 ( .A(n_67), .B(n_631), .Y(n_641) );
INVxp67_ASAP7_75t_SL g662 ( .A(n_67), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_68), .B(n_122), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_69), .B(n_139), .Y(n_231) );
INVx2_ASAP7_75t_L g543 ( .A(n_71), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_72), .B(n_93), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_73), .Y(n_203) );
INVx1_ASAP7_75t_L g198 ( .A(n_74), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_75), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_76), .B(n_208), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_97), .B(n_521), .Y(n_77) );
CKINVDCx6p67_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
CKINVDCx11_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
BUFx6f_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NOR2xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_88), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
AO31x2_ASAP7_75t_L g314 ( .A1(n_83), .A2(n_138), .A3(n_315), .B(n_316), .Y(n_314) );
AO31x2_ASAP7_75t_L g347 ( .A1(n_83), .A2(n_138), .A3(n_315), .B(n_316), .Y(n_347) );
BUFx2_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
OAI21xp33_ASAP7_75t_L g248 ( .A1(n_85), .A2(n_242), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
BUFx6f_ASAP7_75t_SL g163 ( .A(n_86), .Y(n_163) );
INVx2_ASAP7_75t_L g185 ( .A(n_86), .Y(n_185) );
INVx3_ASAP7_75t_L g201 ( .A(n_86), .Y(n_201) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_87), .Y(n_705) );
AO21x2_ASAP7_75t_L g751 ( .A1(n_88), .A2(n_704), .B(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g88 ( .A(n_89), .B(n_92), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
AOI22x1_ASAP7_75t_L g114 ( .A1(n_90), .A2(n_115), .B1(n_126), .B2(n_133), .Y(n_114) );
INVx1_ASAP7_75t_L g247 ( .A(n_90), .Y(n_247) );
AOI21x1_ASAP7_75t_L g256 ( .A1(n_90), .A2(n_257), .B(n_258), .Y(n_256) );
BUFx3_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g162 ( .A(n_91), .Y(n_162) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx2_ASAP7_75t_L g131 ( .A(n_95), .Y(n_131) );
INVx2_ASAP7_75t_L g182 ( .A(n_95), .Y(n_182) );
INVx2_ASAP7_75t_L g284 ( .A(n_95), .Y(n_284) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx2_ASAP7_75t_L g124 ( .A(n_96), .Y(n_124) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
BUFx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
NAND4xp75_ASAP7_75t_L g100 ( .A(n_101), .B(n_367), .C(n_432), .D(n_480), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
NAND3xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_325), .C(n_337), .Y(n_102) );
NOR3xp33_ASAP7_75t_L g103 ( .A(n_104), .B(n_304), .C(n_311), .Y(n_103) );
OAI221xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_216), .B1(n_266), .B2(n_272), .C(n_292), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NOR2x1_ASAP7_75t_L g483 ( .A(n_106), .B(n_484), .Y(n_483) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_166), .Y(n_106) );
INVx1_ASAP7_75t_L g267 ( .A(n_107), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_107), .B(n_383), .Y(n_463) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_141), .Y(n_107) );
INVx1_ASAP7_75t_L g303 ( .A(n_108), .Y(n_303) );
AND2x2_ASAP7_75t_L g306 ( .A(n_108), .B(n_169), .Y(n_306) );
AND2x4_ASAP7_75t_L g360 ( .A(n_108), .B(n_168), .Y(n_360) );
OAI21x1_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_114), .B(n_137), .Y(n_108) );
OAI21x1_ASAP7_75t_L g219 ( .A1(n_109), .A2(n_220), .B(n_231), .Y(n_219) );
OAI21x1_ASAP7_75t_L g353 ( .A1(n_109), .A2(n_220), .B(n_231), .Y(n_353) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NOR2x1_ASAP7_75t_SL g289 ( .A(n_110), .B(n_290), .Y(n_289) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g324 ( .A(n_111), .Y(n_324) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g140 ( .A(n_112), .Y(n_140) );
BUFx2_ASAP7_75t_L g144 ( .A(n_112), .Y(n_144) );
INVx1_ASAP7_75t_L g194 ( .A(n_113), .Y(n_194) );
INVx2_ASAP7_75t_L g315 ( .A(n_114), .Y(n_315) );
OAI22x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_120), .B1(n_121), .B2(n_125), .Y(n_115) );
INVxp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g128 ( .A(n_118), .Y(n_128) );
INVx2_ASAP7_75t_L g176 ( .A(n_118), .Y(n_176) );
INVx2_ASAP7_75t_L g180 ( .A(n_118), .Y(n_180) );
INVx2_ASAP7_75t_L g223 ( .A(n_118), .Y(n_223) );
INVx3_ASAP7_75t_L g237 ( .A(n_118), .Y(n_237) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g155 ( .A(n_119), .Y(n_155) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_119), .Y(n_160) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g225 ( .A(n_123), .Y(n_225) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_123), .Y(n_240) );
INVx2_ASAP7_75t_L g259 ( .A(n_123), .Y(n_259) );
INVx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_124), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_129), .B1(n_130), .B2(n_132), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVxp67_ASAP7_75t_L g147 ( .A(n_128), .Y(n_147) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AOI21x1_ASAP7_75t_SL g235 ( .A1(n_133), .A2(n_236), .B(n_239), .Y(n_235) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_134), .A2(n_281), .B(n_282), .Y(n_280) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g206 ( .A(n_135), .Y(n_206) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx3_ASAP7_75t_L g226 ( .A(n_136), .Y(n_226) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_139), .Y(n_165) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g296 ( .A(n_141), .Y(n_296) );
AND2x2_ASAP7_75t_L g307 ( .A(n_141), .B(n_188), .Y(n_307) );
INVx1_ASAP7_75t_L g344 ( .A(n_141), .Y(n_344) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_141), .Y(n_381) );
INVx3_ASAP7_75t_L g428 ( .A(n_141), .Y(n_428) );
INVx2_ASAP7_75t_L g441 ( .A(n_141), .Y(n_441) );
AND2x2_ASAP7_75t_L g479 ( .A(n_141), .B(n_187), .Y(n_479) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OAI21x1_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_145), .B(n_164), .Y(n_142) );
OAI21x1_ASAP7_75t_L g170 ( .A1(n_143), .A2(n_171), .B(n_186), .Y(n_170) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OAI21x1_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_156), .B(n_163), .Y(n_145) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_150), .Y(n_146) );
INVx2_ASAP7_75t_L g153 ( .A(n_149), .Y(n_153) );
INVx2_ASAP7_75t_L g183 ( .A(n_149), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_149), .B(n_201), .Y(n_200) );
NOR3xp33_ASAP7_75t_L g209 ( .A(n_149), .B(n_201), .C(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_154), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g174 ( .A(n_155), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_161), .Y(n_156) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g204 ( .A(n_160), .Y(n_204) );
INVx2_ASAP7_75t_L g245 ( .A(n_160), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_161), .A2(n_173), .B(n_175), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_161), .A2(n_228), .B(n_229), .Y(n_227) );
BUFx10_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g262 ( .A(n_162), .Y(n_262) );
OAI21x1_ASAP7_75t_L g220 ( .A1(n_163), .A2(n_221), .B(n_227), .Y(n_220) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_165), .Y(n_254) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_187), .Y(n_167) );
OR2x2_ASAP7_75t_L g397 ( .A(n_168), .B(n_347), .Y(n_397) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g269 ( .A(n_169), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g297 ( .A(n_169), .Y(n_297) );
INVx2_ASAP7_75t_L g318 ( .A(n_169), .Y(n_318) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_177), .B(n_184), .Y(n_171) );
O2A1O1Ixp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_181), .C(n_183), .Y(n_177) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_184), .A2(n_256), .B(n_260), .Y(n_255) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_SL g291 ( .A(n_185), .Y(n_291) );
BUFx2_ASAP7_75t_L g300 ( .A(n_187), .Y(n_300) );
NOR2x1_ASAP7_75t_L g317 ( .A(n_187), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_187), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g395 ( .A(n_187), .Y(n_395) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_195), .B(n_214), .Y(n_188) );
AO21x1_ASAP7_75t_L g271 ( .A1(n_189), .A2(n_195), .B(n_214), .Y(n_271) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_SL g214 ( .A(n_190), .B(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AOI21x1_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_194), .Y(n_191) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_192), .A2(n_193), .B(n_194), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_207), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_200), .B1(n_202), .B2(n_205), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
INVx1_ASAP7_75t_L g213 ( .A(n_199), .Y(n_213) );
INVx2_ASAP7_75t_L g230 ( .A(n_199), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_201), .B(n_206), .Y(n_205) );
NOR3xp33_ASAP7_75t_L g211 ( .A(n_201), .B(n_206), .C(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
INVx2_ASAP7_75t_L g208 ( .A(n_204), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B1(n_211), .B2(n_213), .Y(n_207) );
OR2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_232), .Y(n_216) );
OR2x2_ASAP7_75t_L g309 ( .A(n_217), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g326 ( .A(n_217), .B(n_276), .Y(n_326) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_218), .B(n_351), .Y(n_357) );
BUFx3_ASAP7_75t_L g363 ( .A(n_218), .Y(n_363) );
AND2x4_ASAP7_75t_L g409 ( .A(n_218), .B(n_358), .Y(n_409) );
AND2x2_ASAP7_75t_L g472 ( .A(n_218), .B(n_366), .Y(n_472) );
AND2x2_ASAP7_75t_L g520 ( .A(n_218), .B(n_274), .Y(n_520) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_219), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_224), .B(n_226), .Y(n_221) );
INVx2_ASAP7_75t_L g288 ( .A(n_226), .Y(n_288) );
INVxp67_ASAP7_75t_L g263 ( .A(n_230), .Y(n_263) );
OR2x2_ASAP7_75t_L g402 ( .A(n_232), .B(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g517 ( .A(n_232), .B(n_275), .Y(n_517) );
OR2x6_ASAP7_75t_L g232 ( .A(n_233), .B(n_251), .Y(n_232) );
OR2x2_ASAP7_75t_SL g321 ( .A(n_233), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g358 ( .A(n_233), .Y(n_358) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g274 ( .A(n_234), .Y(n_274) );
OAI21x1_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_241), .B(n_248), .Y(n_234) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVxp67_ASAP7_75t_L g316 ( .A(n_249), .Y(n_316) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g376 ( .A(n_251), .B(n_353), .Y(n_376) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g302 ( .A(n_252), .Y(n_302) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_252), .Y(n_365) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B(n_265), .Y(n_253) );
OA21x2_ASAP7_75t_L g322 ( .A1(n_255), .A2(n_265), .B(n_323), .Y(n_322) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_263), .B(n_264), .Y(n_260) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
OAI22xp33_ASAP7_75t_L g413 ( .A1(n_267), .A2(n_414), .B1(n_415), .B2(n_416), .Y(n_413) );
OR2x2_ASAP7_75t_L g426 ( .A(n_268), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g335 ( .A(n_269), .Y(n_335) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_269), .Y(n_448) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_271), .B(n_303), .Y(n_385) );
AND2x2_ASAP7_75t_L g440 ( .A(n_271), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g299 ( .A(n_274), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_274), .B(n_302), .Y(n_310) );
AND2x2_ASAP7_75t_L g328 ( .A(n_274), .B(n_322), .Y(n_328) );
AND2x4_ASAP7_75t_L g352 ( .A(n_274), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g444 ( .A(n_275), .Y(n_444) );
AND2x2_ASAP7_75t_L g476 ( .A(n_275), .B(n_358), .Y(n_476) );
NOR2xp67_ASAP7_75t_R g490 ( .A(n_275), .B(n_298), .Y(n_490) );
OR2x2_ASAP7_75t_L g496 ( .A(n_275), .B(n_296), .Y(n_496) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g295 ( .A(n_276), .Y(n_295) );
INVx2_ASAP7_75t_L g366 ( .A(n_276), .Y(n_366) );
BUFx2_ASAP7_75t_L g403 ( .A(n_276), .Y(n_403) );
AND2x2_ASAP7_75t_L g410 ( .A(n_276), .B(n_322), .Y(n_410) );
AND2x4_ASAP7_75t_L g424 ( .A(n_276), .B(n_302), .Y(n_424) );
OR2x2_ASAP7_75t_L g506 ( .A(n_276), .B(n_365), .Y(n_506) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2x1_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
OAI21x1_ASAP7_75t_SL g279 ( .A1(n_280), .A2(n_285), .B(n_289), .Y(n_279) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVxp67_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
NOR5xp2_ASAP7_75t_L g293 ( .A(n_294), .B(n_298), .C(n_300), .D(n_301), .E(n_303), .Y(n_293) );
NAND3xp33_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .C(n_297), .Y(n_294) );
INVx2_ASAP7_75t_L g320 ( .A(n_295), .Y(n_320) );
INVx2_ASAP7_75t_L g332 ( .A(n_296), .Y(n_332) );
AND2x2_ASAP7_75t_L g461 ( .A(n_296), .B(n_345), .Y(n_461) );
AND2x2_ASAP7_75t_L g345 ( .A(n_297), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g420 ( .A(n_297), .Y(n_420) );
AND2x2_ASAP7_75t_L g485 ( .A(n_297), .B(n_395), .Y(n_485) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g406 ( .A(n_299), .B(n_376), .Y(n_406) );
AND2x2_ASAP7_75t_L g437 ( .A(n_300), .B(n_360), .Y(n_437) );
AOI32xp33_ASAP7_75t_L g510 ( .A1(n_300), .A2(n_511), .A3(n_513), .B1(n_514), .B2(n_515), .Y(n_510) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g351 ( .A(n_302), .Y(n_351) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_308), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
AND2x2_ASAP7_75t_L g439 ( .A(n_306), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g359 ( .A(n_307), .B(n_360), .Y(n_359) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_307), .Y(n_492) );
AND2x2_ASAP7_75t_L g515 ( .A(n_307), .B(n_313), .Y(n_515) );
AO21x1_ASAP7_75t_L g481 ( .A1(n_308), .A2(n_482), .B(n_486), .Y(n_481) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g340 ( .A(n_310), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_319), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_317), .Y(n_312) );
INVx1_ASAP7_75t_L g513 ( .A(n_313), .Y(n_513) );
BUFx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g336 ( .A(n_314), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_317), .B(n_380), .Y(n_412) );
INVxp67_ASAP7_75t_SL g474 ( .A(n_317), .Y(n_474) );
INVx1_ASAP7_75t_L g383 ( .A(n_318), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_318), .B(n_428), .Y(n_500) );
NOR2xp67_ASAP7_75t_L g503 ( .A(n_318), .B(n_427), .Y(n_503) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x2_ASAP7_75t_L g327 ( .A(n_320), .B(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g378 ( .A(n_321), .Y(n_378) );
OR2x2_ASAP7_75t_L g450 ( .A(n_321), .B(n_353), .Y(n_450) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
OAI21xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B(n_329), .Y(n_325) );
INVx2_ASAP7_75t_L g477 ( .A(n_327), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_328), .B(n_363), .Y(n_414) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2x1p5_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_331), .A2(n_456), .B(n_517), .C(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NOR2x1p5_ASAP7_75t_L g396 ( .A(n_332), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g447 ( .A(n_332), .B(n_448), .Y(n_447) );
NAND3xp33_ASAP7_75t_L g475 ( .A(n_332), .B(n_363), .C(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g348 ( .A(n_334), .Y(n_348) );
INVx3_ASAP7_75t_L g446 ( .A(n_334), .Y(n_446) );
OR2x6_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_336), .B(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_354), .Y(n_337) );
AOI22x1_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_341), .B1(n_348), .B2(n_349), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g443 ( .A(n_340), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_340), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g508 ( .A(n_341), .Y(n_508) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_345), .Y(n_341) );
INVx1_ASAP7_75t_L g421 ( .A(n_342), .Y(n_421) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g399 ( .A(n_345), .Y(n_399) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g467 ( .A(n_347), .B(n_428), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_348), .A2(n_355), .B1(n_359), .B2(n_361), .Y(n_354) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_350), .B(n_431), .Y(n_430) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g371 ( .A(n_352), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_352), .B(n_391), .Y(n_460) );
NOR2x1_ASAP7_75t_L g511 ( .A(n_352), .B(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g514 ( .A(n_352), .B(n_410), .Y(n_514) );
INVxp67_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
OR2x2_ASAP7_75t_L g469 ( .A(n_357), .B(n_391), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_360), .B(n_380), .Y(n_415) );
INVx2_ASAP7_75t_L g456 ( .A(n_360), .Y(n_456) );
INVx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
OR2x2_ASAP7_75t_L g401 ( .A(n_363), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_363), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g431 ( .A(n_363), .Y(n_431) );
BUFx3_ASAP7_75t_L g457 ( .A(n_364), .Y(n_457) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
BUFx2_ASAP7_75t_L g372 ( .A(n_366), .Y(n_372) );
INVx1_ASAP7_75t_L g391 ( .A(n_366), .Y(n_391) );
AND4x1_ASAP7_75t_L g367 ( .A(n_368), .B(n_386), .C(n_404), .D(n_417), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI31xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_373), .A3(n_377), .B(n_379), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g501 ( .A(n_378), .B(n_472), .Y(n_501) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVxp67_ASAP7_75t_SL g407 ( .A(n_382), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g499 ( .A(n_385), .B(n_500), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_392), .B1(n_398), .B2(n_400), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
OR2x2_ASAP7_75t_L g487 ( .A(n_388), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_396), .A2(n_465), .B1(n_468), .B2(n_470), .C(n_473), .Y(n_464) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_402), .B(n_430), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_407), .B1(n_408), .B2(n_411), .C(n_413), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g416 ( .A(n_406), .Y(n_416) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx3_ASAP7_75t_R g458 ( .A(n_409), .Y(n_458) );
INVx2_ASAP7_75t_L g488 ( .A(n_410), .Y(n_488) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g417 ( .A1(n_418), .A2(n_422), .B1(n_425), .B2(n_429), .Y(n_417) );
NOR2xp67_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AOI211xp5_ASAP7_75t_L g486 ( .A1(n_420), .A2(n_487), .B(n_489), .C(n_491), .Y(n_486) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g512 ( .A(n_424), .Y(n_512) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g504 ( .A(n_431), .B(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g509 ( .A(n_431), .B(n_488), .Y(n_509) );
NOR2x1_ASAP7_75t_L g432 ( .A(n_433), .B(n_451), .Y(n_432) );
OAI21xp5_ASAP7_75t_SL g433 ( .A1(n_434), .A2(n_442), .B(n_445), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI221xp5_ASAP7_75t_L g507 ( .A1(n_438), .A2(n_469), .B1(n_508), .B2(n_509), .C(n_510), .Y(n_507) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g455 ( .A(n_440), .Y(n_455) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI21xp33_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B(n_449), .Y(n_445) );
NAND2x1_ASAP7_75t_L g494 ( .A(n_446), .B(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g465 ( .A(n_448), .B(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_464), .Y(n_451) );
AOI322xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_457), .A3(n_458), .B1(n_459), .B2(n_461), .C1(n_462), .C2(n_755), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
OAI21xp33_ASAP7_75t_L g493 ( .A1(n_458), .A2(n_494), .B(n_497), .Y(n_493) );
INVxp67_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x4_ASAP7_75t_L g484 ( .A(n_466), .B(n_485), .Y(n_484) );
INVx2_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OAI22xp33_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B1(n_477), .B2(n_478), .Y(n_473) );
NOR4xp75_ASAP7_75t_L g480 ( .A(n_481), .B(n_493), .C(n_507), .D(n_516), .Y(n_480) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVxp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_501), .B1(n_502), .B2(n_504), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g518 ( .A(n_506), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OAI221xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_698), .B2(n_708), .C(n_747), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_523), .A2(n_748), .B1(n_750), .B2(n_751), .Y(n_747) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_529), .B(n_618), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OR2x6_ASAP7_75t_L g694 ( .A(n_527), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x4_ASAP7_75t_L g623 ( .A(n_528), .B(n_624), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g648 ( .A(n_528), .B(n_649), .Y(n_648) );
AND2x4_ASAP7_75t_SL g663 ( .A(n_528), .B(n_649), .Y(n_663) );
AND3x1_ASAP7_75t_L g679 ( .A(n_528), .B(n_680), .C(n_682), .Y(n_679) );
NAND4xp25_ASAP7_75t_SL g529 ( .A(n_530), .B(n_552), .C(n_602), .D(n_611), .Y(n_529) );
AOI21xp33_ASAP7_75t_SL g530 ( .A1(n_531), .A2(n_544), .B(n_545), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_534), .B(n_539), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_536), .Y(n_570) );
INVx2_ASAP7_75t_L g576 ( .A(n_536), .Y(n_576) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
INVx2_ASAP7_75t_L g550 ( .A(n_537), .Y(n_550) );
AND2x2_ASAP7_75t_L g573 ( .A(n_537), .B(n_551), .Y(n_573) );
INVx2_ASAP7_75t_L g551 ( .A(n_538), .Y(n_551) );
AND2x4_ASAP7_75t_L g547 ( .A(n_539), .B(n_548), .Y(n_547) );
NAND2x1p5_ASAP7_75t_L g598 ( .A(n_539), .B(n_599), .Y(n_598) );
BUFx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g597 ( .A(n_540), .Y(n_597) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
OR2x2_ASAP7_75t_L g565 ( .A(n_541), .B(n_542), .Y(n_565) );
AND2x4_ASAP7_75t_L g583 ( .A(n_541), .B(n_584), .Y(n_583) );
OR2x6_ASAP7_75t_L g606 ( .A(n_541), .B(n_543), .Y(n_606) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx2_ASAP7_75t_L g584 ( .A(n_543), .Y(n_584) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x4_ASAP7_75t_L g610 ( .A(n_548), .B(n_605), .Y(n_610) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g562 ( .A(n_549), .Y(n_562) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_549), .Y(n_580) );
AND2x4_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
AND2x4_ASAP7_75t_L g558 ( .A(n_550), .B(n_559), .Y(n_558) );
AOI221xp5_ASAP7_75t_SL g552 ( .A1(n_553), .A2(n_566), .B1(n_574), .B2(n_585), .C(n_590), .Y(n_552) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx3_ASAP7_75t_L g589 ( .A(n_557), .Y(n_589) );
INVx4_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx12f_ASAP7_75t_L g617 ( .A(n_558), .Y(n_617) );
INVx1_ASAP7_75t_L g601 ( .A(n_559), .Y(n_601) );
BUFx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx4_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
BUFx6f_ASAP7_75t_L g734 ( .A(n_565), .Y(n_734) );
CKINVDCx14_ASAP7_75t_R g567 ( .A(n_568), .Y(n_567) );
CKINVDCx14_ASAP7_75t_R g568 ( .A(n_569), .Y(n_568) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x4_ASAP7_75t_L g604 ( .A(n_570), .B(n_605), .Y(n_604) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_571), .Y(n_586) );
BUFx12f_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g614 ( .A(n_572), .B(n_605), .Y(n_614) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_579), .Y(n_578) );
BUFx6f_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_582), .Y(n_581) );
BUFx6f_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_SL g739 ( .A(n_593), .Y(n_739) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g731 ( .A(n_594), .B(n_732), .C(n_734), .Y(n_731) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B1(n_607), .B2(n_608), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_603), .A2(n_684), .B1(n_686), .B2(n_688), .C(n_689), .Y(n_683) );
AND2x2_ASAP7_75t_L g616 ( .A(n_605), .B(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B1(n_615), .B2(n_616), .Y(n_611) );
BUFx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AOI211xp5_ASAP7_75t_L g645 ( .A1(n_615), .A2(n_646), .B(n_650), .C(n_664), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_645), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_637), .Y(n_619) );
OR2x6_ASAP7_75t_L g621 ( .A(n_622), .B(n_626), .Y(n_621) );
OR2x2_ASAP7_75t_L g632 ( .A(n_622), .B(n_633), .Y(n_632) );
OR2x6_ASAP7_75t_L g638 ( .A(n_622), .B(n_639), .Y(n_638) );
OR2x6_ASAP7_75t_L g642 ( .A(n_622), .B(n_643), .Y(n_642) );
INVx4_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g681 ( .A(n_625), .Y(n_681) );
OR2x6_ASAP7_75t_L g697 ( .A(n_626), .B(n_648), .Y(n_697) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
BUFx12f_ASAP7_75t_L g669 ( .A(n_627), .Y(n_669) );
NAND2x1p5_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x4_ASAP7_75t_L g635 ( .A(n_629), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_629), .B(n_631), .Y(n_644) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g636 ( .A(n_631), .Y(n_636) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx2_ASAP7_75t_L g691 ( .A(n_634), .Y(n_691) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_635), .Y(n_676) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_636), .Y(n_655) );
INVx2_ASAP7_75t_L g690 ( .A(n_639), .Y(n_690) );
INVx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
BUFx4f_ASAP7_75t_L g674 ( .A(n_641), .Y(n_674) );
OR2x4_ASAP7_75t_L g647 ( .A(n_643), .B(n_648), .Y(n_647) );
BUFx3_ASAP7_75t_L g666 ( .A(n_643), .Y(n_666) );
INVx1_ASAP7_75t_L g685 ( .A(n_643), .Y(n_685) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OR2x6_ASAP7_75t_L g653 ( .A(n_648), .B(n_654), .Y(n_653) );
INVx4_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx5_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
BUFx4f_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x4_ASAP7_75t_L g658 ( .A(n_659), .B(n_663), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_677), .B1(n_683), .B2(n_692), .C(n_697), .Y(n_664) );
OAI221xp5_ASAP7_75t_SL g665 ( .A1(n_666), .A2(n_667), .B1(n_668), .B2(n_670), .C(n_671), .Y(n_665) );
BUFx3_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_SL g687 ( .A(n_669), .Y(n_687) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
BUFx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx3_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_699), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_700), .Y(n_699) );
BUFx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
BUFx6f_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_706), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
BUFx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g729 ( .A(n_705), .Y(n_729) );
AND2x2_ASAP7_75t_L g752 ( .A(n_706), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_707), .B(n_729), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_725), .B1(n_740), .B2(n_741), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_709), .A2(n_740), .B1(n_743), .B2(n_749), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_714), .B1(n_723), .B2(n_724), .Y(n_709) );
INVx1_ASAP7_75t_L g723 ( .A(n_710), .Y(n_723) );
INVx1_ASAP7_75t_L g713 ( .A(n_711), .Y(n_713) );
INVx1_ASAP7_75t_L g724 ( .A(n_714), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_717), .B1(n_718), .B2(n_722), .Y(n_714) );
INVx1_ASAP7_75t_L g722 ( .A(n_715), .Y(n_722) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g721 ( .A(n_720), .Y(n_721) );
BUFx3_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx5_ASAP7_75t_L g749 ( .A(n_726), .Y(n_749) );
AND2x6_ASAP7_75t_L g726 ( .A(n_727), .B(n_735), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_728), .B(n_730), .Y(n_727) );
INVxp67_ASAP7_75t_L g745 ( .A(n_728), .Y(n_745) );
INVx1_ASAP7_75t_L g753 ( .A(n_729), .Y(n_753) );
INVxp67_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_731), .B(n_739), .Y(n_746) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
CKINVDCx11_ASAP7_75t_R g737 ( .A(n_733), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
CKINVDCx5p33_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx3_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
BUFx4f_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx4_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
endmodule