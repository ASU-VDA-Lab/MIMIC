module fake_jpeg_19360_n_253 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_253);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_145;
wire n_18;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx24_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_23),
.B(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_15),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_10),
.B(n_5),
.Y(n_30)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_5),
.Y(n_32)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx9p33_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx2_ASAP7_75t_SL g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_14),
.B1(n_15),
.B2(n_11),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_52),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_49),
.B(n_54),
.Y(n_63)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_41),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_26),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_14),
.B1(n_15),
.B2(n_25),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_56),
.B(n_37),
.C(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_10),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_14),
.B1(n_25),
.B2(n_27),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_27),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_41),
.C(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_41),
.C(n_38),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_69),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_37),
.B1(n_39),
.B2(n_56),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_50),
.B1(n_52),
.B2(n_44),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_61),
.B1(n_62),
.B2(n_59),
.Y(n_94)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_77),
.Y(n_98)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_85),
.Y(n_101)
);

NOR2x1_ASAP7_75t_SL g79 ( 
.A(n_72),
.B(n_50),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_31),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_45),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_82),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_73),
.B(n_50),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_84),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_48),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_61),
.B(n_53),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_60),
.B1(n_63),
.B2(n_67),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_88),
.A2(n_67),
.B1(n_65),
.B2(n_64),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_94),
.B(n_97),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_47),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_85),
.B1(n_79),
.B2(n_86),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_82),
.B1(n_78),
.B2(n_33),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_70),
.B1(n_58),
.B2(n_66),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_77),
.B1(n_49),
.B2(n_43),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_39),
.B1(n_51),
.B2(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_107),
.B(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_39),
.B1(n_51),
.B2(n_58),
.Y(n_109)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_113),
.B(n_104),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_75),
.Y(n_114)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_133),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_99),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_124),
.Y(n_136)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_36),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_125),
.B(n_126),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_91),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_36),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_127),
.B(n_128),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_36),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_78),
.C(n_38),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_68),
.C(n_104),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_10),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_12),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_36),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_132),
.B(n_119),
.Y(n_158)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_94),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_116),
.A2(n_93),
.B(n_105),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_92),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_111),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_145),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_113),
.Y(n_146)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_111),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_148),
.B(n_152),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_150),
.C(n_134),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_112),
.Y(n_151)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_19),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_19),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_154),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_121),
.A2(n_17),
.B(n_13),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_157),
.B(n_126),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_33),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_156),
.B(n_120),
.Y(n_171)
);

NAND2x1p5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_120),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_158),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_171),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_115),
.C(n_133),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_165),
.C(n_145),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_121),
.B1(n_130),
.B2(n_123),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_164),
.A2(n_166),
.B1(n_174),
.B2(n_144),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_124),
.C(n_122),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_118),
.B1(n_122),
.B2(n_112),
.Y(n_166)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_139),
.A2(n_131),
.B1(n_39),
.B2(n_17),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_176),
.B1(n_13),
.B2(n_17),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_131),
.B1(n_55),
.B2(n_34),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_157),
.B1(n_149),
.B2(n_140),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_150),
.C(n_137),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_182),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_142),
.C(n_135),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_189),
.C(n_192),
.Y(n_196)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_151),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_186),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_145),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_55),
.C(n_22),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_34),
.B1(n_12),
.B2(n_13),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_28),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_4),
.B1(n_9),
.B2(n_2),
.Y(n_192)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_161),
.A2(n_12),
.B(n_21),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_193),
.A2(n_170),
.B(n_163),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_168),
.C(n_171),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_173),
.C(n_164),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_34),
.C(n_24),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_28),
.C(n_24),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_22),
.C(n_18),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_179),
.C(n_185),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_205),
.Y(n_219)
);

BUFx12_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_209),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_174),
.C(n_169),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_206),
.A2(n_208),
.B1(n_28),
.B2(n_24),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_SL g208 ( 
.A(n_190),
.B(n_169),
.C(n_18),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_209),
.A2(n_180),
.B1(n_191),
.B2(n_18),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_197),
.A2(n_188),
.B(n_186),
.Y(n_210)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_214),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_203),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_18),
.C(n_16),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_204),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_220),
.C(n_20),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_18),
.B(n_16),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_206),
.B(n_198),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_18),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_218),
.A2(n_198),
.B1(n_1),
.B2(n_0),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_29),
.C(n_16),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_221),
.B(n_225),
.Y(n_231)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_20),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_208),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_227),
.B(n_228),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_213),
.A2(n_216),
.B(n_218),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_229),
.A2(n_220),
.B(n_6),
.Y(n_232)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_228),
.Y(n_230)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_232),
.A2(n_235),
.B(n_237),
.Y(n_238)
);

AOI322xp5_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_20),
.A3(n_7),
.B1(n_2),
.B2(n_3),
.C1(n_8),
.C2(n_9),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_226),
.A2(n_20),
.B(n_4),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_4),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_222),
.C(n_221),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_243),
.B(n_3),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_242),
.B(n_238),
.Y(n_246)
);

NOR3xp33_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_234),
.C(n_3),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_234),
.A2(n_3),
.B(n_7),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_246),
.A2(n_7),
.B(n_9),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_247),
.A2(n_7),
.B(n_9),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_248),
.B(n_0),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_250),
.A2(n_0),
.B(n_1),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_0),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_0),
.Y(n_253)
);


endmodule