module fake_jpeg_446_n_63 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_63);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_63;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx4_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_0),
.B(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_8),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_2),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_24),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_10),
.B(n_2),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_23),
.B(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_3),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_9),
.B1(n_14),
.B2(n_12),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_39),
.B1(n_26),
.B2(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_26),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

AO221x1_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_48),
.B1(n_32),
.B2(n_40),
.C(n_39),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_44),
.B(n_47),
.C(n_4),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_25),
.B(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_11),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_27),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_32),
.B1(n_31),
.B2(n_40),
.Y(n_51)
);

NAND5xp2_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_29),
.C(n_17),
.D(n_24),
.E(n_5),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_52),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_44),
.Y(n_54)
);

XNOR2x1_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_55),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_47),
.B(n_46),
.Y(n_57)
);

NAND4xp25_ASAP7_75t_SL g59 ( 
.A(n_57),
.B(n_52),
.C(n_54),
.D(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_7),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_62),
.Y(n_63)
);


endmodule