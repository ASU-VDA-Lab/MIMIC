module real_jpeg_6369_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_323;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_1),
.A2(n_39),
.B1(n_43),
.B2(n_45),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_1),
.A2(n_45),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_1),
.A2(n_45),
.B1(n_51),
.B2(n_56),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_1),
.A2(n_45),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_2),
.A2(n_242),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_2),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_2),
.A2(n_152),
.B1(n_279),
.B2(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_2),
.A2(n_279),
.B1(n_379),
.B2(n_382),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_2),
.A2(n_169),
.B1(n_279),
.B2(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_4),
.A2(n_118),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_4),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_4),
.A2(n_186),
.B1(n_228),
.B2(n_269),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_4),
.A2(n_186),
.B1(n_386),
.B2(n_388),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_4),
.A2(n_186),
.B1(n_449),
.B2(n_450),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_5),
.A2(n_49),
.B1(n_50),
.B2(n_55),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_5),
.A2(n_49),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_5),
.A2(n_49),
.B1(n_95),
.B2(n_99),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_5),
.A2(n_49),
.B1(n_258),
.B2(n_264),
.Y(n_263)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_6),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_7),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_7),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_8),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_8),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_8),
.A2(n_56),
.B1(n_132),
.B2(n_179),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_8),
.A2(n_95),
.B1(n_132),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_8),
.A2(n_132),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_9),
.A2(n_122),
.B1(n_273),
.B2(n_276),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_9),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_9),
.A2(n_194),
.B1(n_276),
.B2(n_324),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_9),
.A2(n_56),
.B1(n_276),
.B2(n_371),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_9),
.A2(n_276),
.B1(n_406),
.B2(n_408),
.Y(n_405)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_10),
.Y(n_98)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_10),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_10),
.Y(n_113)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_11),
.Y(n_106)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_12),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_12),
.Y(n_100)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_12),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_12),
.Y(n_119)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_12),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_12),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_12),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_12),
.Y(n_282)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_13),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_14),
.A2(n_82),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_14),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_14),
.A2(n_86),
.B1(n_100),
.B2(n_122),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_14),
.A2(n_86),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_14),
.A2(n_86),
.B1(n_144),
.B2(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_15),
.B(n_252),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_15),
.A2(n_99),
.B(n_251),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_15),
.B(n_188),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_15),
.B(n_355),
.C(n_359),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_L g364 ( 
.A1(n_15),
.A2(n_365),
.B1(n_366),
.B2(n_369),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_15),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_15),
.B(n_149),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_15),
.A2(n_25),
.B1(n_405),
.B2(n_413),
.Y(n_412)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_494),
.C(n_498),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_492),
.B(n_496),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_482),
.B(n_491),
.Y(n_18)
);

OAI31xp33_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_214),
.A3(n_232),
.B(n_479),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_196),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_21),
.B(n_196),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_125),
.C(n_160),
.Y(n_21)
);

FAx1_ASAP7_75t_SL g342 ( 
.A(n_22),
.B(n_125),
.CI(n_160),
.CON(n_342),
.SN(n_342)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_89),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g213 ( 
.A1(n_23),
.A2(n_24),
.B(n_91),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_46),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_24),
.A2(n_90),
.B1(n_91),
.B2(n_124),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_24),
.A2(n_46),
.B1(n_90),
.B2(n_334),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_34),
.B(n_38),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_25),
.B(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_25),
.A2(n_255),
.B1(n_261),
.B2(n_263),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_25),
.A2(n_263),
.B(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_25),
.A2(n_172),
.B(n_385),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_25),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_25),
.A2(n_395),
.B1(n_405),
.B2(n_409),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_25),
.A2(n_38),
.B(n_297),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_26),
.Y(n_396)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_28),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_30),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_30),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_31),
.B(n_298),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_31),
.A2(n_164),
.B(n_256),
.Y(n_318)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_33),
.Y(n_417)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_34),
.Y(n_399)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_37),
.Y(n_174)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_38),
.Y(n_173)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_42),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_72),
.B1(n_75),
.B2(n_77),
.Y(n_71)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_43),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_43),
.Y(n_260)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g390 ( 
.A(n_44),
.Y(n_390)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_44),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_46),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_58),
.B(n_78),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_48),
.A2(n_59),
.B1(n_79),
.B2(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_53),
.Y(n_180)
);

INVx6_ASAP7_75t_L g353 ( 
.A(n_53),
.Y(n_353)
);

INVx6_ASAP7_75t_L g368 ( 
.A(n_53),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_53),
.Y(n_451)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_54),
.Y(n_369)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_54),
.Y(n_381)
);

BUFx5_ASAP7_75t_L g382 ( 
.A(n_54),
.Y(n_382)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_54),
.Y(n_442)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_57),
.A2(n_136),
.B1(n_137),
.B2(n_140),
.Y(n_135)
);

INVx5_ASAP7_75t_L g372 ( 
.A(n_57),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_58),
.B(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_58),
.A2(n_80),
.B(n_156),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_58),
.A2(n_78),
.B(n_156),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_58),
.A2(n_80),
.B1(n_158),
.B2(n_178),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_58),
.A2(n_463),
.B(n_464),
.Y(n_462)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_59),
.A2(n_79),
.B1(n_364),
.B2(n_370),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_59),
.A2(n_79),
.B1(n_370),
.B2(n_378),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_59),
.A2(n_79),
.B1(n_378),
.B2(n_448),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_71),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B1(n_66),
.B2(n_69),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g358 ( 
.A(n_68),
.Y(n_358)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_80),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_80),
.B(n_365),
.Y(n_403)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_88),
.Y(n_431)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_114),
.B(n_120),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_92),
.B(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_92),
.A2(n_188),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_92),
.A2(n_188),
.B1(n_272),
.B2(n_277),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_92),
.A2(n_114),
.B(n_188),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_93),
.A2(n_183),
.B(n_187),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_93),
.A2(n_123),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_93),
.A2(n_123),
.B1(n_183),
.B2(n_278),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_93),
.A2(n_488),
.B(n_489),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_97),
.B1(n_99),
.B2(n_101),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_107),
.B1(n_109),
.B2(n_112),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_106),
.Y(n_241)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_111),
.Y(n_270)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_112),
.Y(n_245)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_113),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_114),
.B(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_119),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_120),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_121),
.Y(n_211)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_122),
.Y(n_243)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_123),
.A2(n_207),
.B(n_210),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_154),
.B(n_159),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_154),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_134),
.B1(n_149),
.B2(n_150),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_128),
.A2(n_135),
.B(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_131),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_131),
.Y(n_435)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_134),
.B(n_192),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_134),
.A2(n_150),
.B(n_202),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_134),
.A2(n_225),
.B(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_134),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_134),
.A2(n_149),
.B1(n_323),
.B2(n_446),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_134),
.A2(n_149),
.B(n_486),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_143),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_135),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_135),
.A2(n_289),
.B1(n_293),
.B2(n_294),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_135),
.A2(n_289),
.B1(n_293),
.B2(n_322),
.Y(n_321)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_139),
.Y(n_438)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_142),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_145),
.Y(n_227)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_147),
.Y(n_247)
);

INVx6_ASAP7_75t_L g432 ( 
.A(n_148),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_149),
.B(n_192),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_SL g446 ( 
.A1(n_151),
.A2(n_365),
.B(n_433),
.Y(n_446)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_153),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_155),
.Y(n_464)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_159),
.B(n_197),
.CI(n_213),
.CON(n_196),
.SN(n_196)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_181),
.C(n_189),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_161),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_175),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_162),
.A2(n_175),
.B1(n_176),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_162),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_172),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_165),
.Y(n_298)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_171),
.Y(n_265)
);

INVx5_ASAP7_75t_L g362 ( 
.A(n_171),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_181),
.A2(n_182),
.B1(n_189),
.B2(n_190),
.Y(n_336)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_187),
.B(n_210),
.Y(n_494)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI32xp33_ASAP7_75t_L g429 ( 
.A1(n_194),
.A2(n_430),
.A3(n_432),
.B1(n_433),
.B2(n_436),
.Y(n_429)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_196),
.B(n_216),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_206),
.B2(n_212),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_199)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_200),
.A2(n_205),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_200),
.B(n_222),
.C(n_229),
.Y(n_490)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_205),
.C(n_206),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_203),
.A2(n_226),
.B(n_293),
.Y(n_308)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_206),
.A2(n_212),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_206),
.B(n_217),
.C(n_220),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_215),
.A2(n_480),
.B(n_481),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_226),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_231),
.Y(n_488)
);

OA21x2_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_343),
.B(n_473),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_328),
.C(n_340),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_312),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_235),
.A2(n_475),
.B(n_476),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_300),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_236),
.B(n_300),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_283),
.C(n_295),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_237),
.B(n_327),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_266),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_238),
.B(n_267),
.C(n_271),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_254),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_239),
.B(n_254),
.Y(n_315)
);

OAI32xp33_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_242),
.A3(n_244),
.B1(n_246),
.B2(n_250),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.Y(n_266)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx8_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_283),
.B(n_295),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.C(n_288),
.Y(n_283)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_284),
.B(n_285),
.CI(n_288),
.CON(n_314),
.SN(n_314)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_299),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_299),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_303),
.C(n_305),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_311),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_310),
.C(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_311),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_326),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_313),
.B(n_326),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.C(n_316),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_314),
.B(n_471),
.Y(n_470)
);

BUFx24_ASAP7_75t_SL g500 ( 
.A(n_314),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_315),
.B(n_316),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.C(n_321),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_317),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_458)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_321),
.B(n_458),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx5_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

A2O1A1O1Ixp25_ASAP7_75t_L g473 ( 
.A1(n_328),
.A2(n_340),
.B(n_474),
.C(n_477),
.D(n_478),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_339),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_329),
.B(n_339),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_332),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_333),
.C(n_338),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_335),
.B1(n_337),
.B2(n_338),
.Y(n_332)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_333),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_335),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_341),
.B(n_342),
.Y(n_478)
);

BUFx24_ASAP7_75t_SL g501 ( 
.A(n_342),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_468),
.B(n_472),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_345),
.A2(n_453),
.B(n_467),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_425),
.B(n_452),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_347),
.A2(n_391),
.B(n_424),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_373),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_348),
.B(n_373),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_363),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_349),
.B(n_363),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_354),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_365),
.B(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_365),
.B(n_434),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_384),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_376),
.B1(n_377),
.B2(n_383),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_375),
.B(n_383),
.C(n_384),
.Y(n_426)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_377),
.Y(n_383)
);

INVx4_ASAP7_75t_SL g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_385),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx8_ASAP7_75t_L g408 ( 
.A(n_387),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_392),
.A2(n_401),
.B(n_423),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_400),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_393),
.B(n_400),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_394),
.A2(n_397),
.B1(n_398),
.B2(n_399),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_402),
.A2(n_411),
.B(n_422),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_403),
.B(n_404),
.Y(n_422)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_409),
.Y(n_414)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_415),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_414),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_418),
.Y(n_415)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_427),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_444),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_445),
.C(n_447),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_443),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_429),
.B(n_443),
.Y(n_461)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_439),
.Y(n_436)
);

INVx6_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_441),
.Y(n_449)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_447),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_448),
.Y(n_463)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_454),
.B(n_455),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_456),
.A2(n_457),
.B1(n_459),
.B2(n_460),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_456),
.B(n_462),
.C(n_465),
.Y(n_469)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_461),
.A2(n_462),
.B1(n_465),
.B2(n_466),
.Y(n_460)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_461),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_462),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_469),
.B(n_470),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_483),
.B(n_484),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_483),
.B(n_484),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_484),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_484),
.B(n_494),
.Y(n_497)
);

FAx1_ASAP7_75t_SL g484 ( 
.A(n_485),
.B(n_487),
.CI(n_490),
.CON(n_484),
.SN(n_484)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_495),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_494),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);


endmodule