module fake_jpeg_28904_n_209 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_209);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_8),
.B(n_11),
.Y(n_14)
);

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_3),
.B(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_13),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_42),
.Y(n_69)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_10),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_51),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_29),
.B(n_10),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_5),
.Y(n_91)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_34),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_75),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_25),
.B1(n_16),
.B2(n_31),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_61),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_25),
.B1(n_16),
.B2(n_31),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_16),
.B1(n_24),
.B2(n_28),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_16),
.B1(n_33),
.B2(n_28),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_39),
.B(n_33),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_22),
.B1(n_20),
.B2(n_18),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_38),
.A2(n_22),
.B1(n_20),
.B2(n_18),
.Y(n_82)
);

OR2x2_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_47),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_83),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_9),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_9),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_36),
.B(n_0),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_37),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_5),
.Y(n_96)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_96),
.B(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_45),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_78),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_59),
.Y(n_134)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_65),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_107),
.A2(n_59),
.B1(n_68),
.B2(n_118),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_50),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_58),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_7),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_69),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_48),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_115),
.Y(n_139)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_48),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_71),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_64),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_72),
.Y(n_128)
);

AOI32xp33_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_80),
.A3(n_61),
.B1(n_63),
.B2(n_90),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_94),
.B(n_119),
.C(n_109),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_118),
.A2(n_77),
.B1(n_67),
.B2(n_92),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_103),
.B1(n_117),
.B2(n_137),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_133),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_71),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_65),
.B1(n_80),
.B2(n_85),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_135),
.A2(n_107),
.B1(n_106),
.B2(n_98),
.Y(n_152)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_94),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_68),
.C(n_99),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_141),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_93),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_104),
.Y(n_142)
);

FAx1_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_124),
.CI(n_126),
.CON(n_162),
.SN(n_162)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_142),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_144),
.B(n_145),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_148),
.B(n_150),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_141),
.B(n_112),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_132),
.B(n_105),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_154),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_153),
.B1(n_156),
.B2(n_142),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_100),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_95),
.B1(n_116),
.B2(n_114),
.Y(n_155)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_133),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_159),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_124),
.Y(n_160)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_135),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_164),
.A2(n_156),
.B1(n_144),
.B2(n_158),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_143),
.C(n_131),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_166),
.B(n_167),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_143),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_149),
.C(n_153),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_158),
.Y(n_172)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_176),
.B(n_182),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_167),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_183),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_162),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_181),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_153),
.C(n_152),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_121),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_164),
.B(n_172),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_SL g193 ( 
.A1(n_186),
.A2(n_179),
.B(n_180),
.C(n_181),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_163),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_130),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_174),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_168),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_188),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_195),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_186),
.A2(n_173),
.B1(n_179),
.B2(n_165),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_123),
.C(n_130),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_196),
.B(n_197),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_199),
.B(n_200),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_187),
.B(n_192),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_201),
.B(n_190),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_204),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g204 ( 
.A1(n_198),
.A2(n_193),
.B(n_123),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_199),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_205),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_206),
.C(n_129),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_129),
.Y(n_209)
);


endmodule