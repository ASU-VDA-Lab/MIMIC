module fake_jpeg_20306_n_186 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_186);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_35),
.B(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx2_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_16),
.Y(n_62)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_1),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_17),
.A2(n_2),
.B(n_3),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_51),
.A2(n_19),
.B(n_17),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_57),
.Y(n_78)
);

FAx1_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_24),
.CI(n_19),
.CON(n_56),
.SN(n_56)
);

NOR2xp33_ASAP7_75t_R g81 ( 
.A(n_56),
.B(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_21),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_27),
.B1(n_16),
.B2(n_29),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_2),
.B(n_3),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_71),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_32),
.B1(n_23),
.B2(n_20),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_66),
.A2(n_47),
.B1(n_50),
.B2(n_43),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_32),
.B1(n_29),
.B2(n_27),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_42),
.B1(n_38),
.B2(n_37),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_32),
.B1(n_21),
.B2(n_25),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_80),
.Y(n_101)
);

OR2x2_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_19),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_81),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_43),
.B1(n_42),
.B2(n_39),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_82),
.A2(n_88),
.B1(n_96),
.B2(n_68),
.Y(n_108)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_90),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_37),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_25),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_92),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_49),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_94),
.Y(n_111)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_24),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_98),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_31),
.B1(n_18),
.B2(n_17),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_3),
.C(n_4),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_72),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_60),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_93),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_69),
.A3(n_58),
.B1(n_51),
.B2(n_64),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_92),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_112),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_108),
.A2(n_89),
.B1(n_76),
.B2(n_90),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_69),
.B1(n_58),
.B2(n_64),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

BUFx24_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_123),
.B1(n_125),
.B2(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_75),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_118),
.B(n_122),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_119),
.A2(n_124),
.B(n_99),
.Y(n_136)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_76),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_85),
.B1(n_80),
.B2(n_98),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_68),
.B1(n_59),
.B2(n_93),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_126),
.B(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_128),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_79),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_100),
.C(n_99),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_130),
.B(n_131),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_133),
.A2(n_59),
.B1(n_87),
.B2(n_84),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_134),
.B(n_138),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_103),
.B(n_51),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_124),
.B(n_128),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_137),
.A2(n_132),
.B(n_136),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_115),
.Y(n_138)
);

NOR4xp25_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_104),
.C(n_106),
.D(n_78),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_109),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_142),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_121),
.B1(n_118),
.B2(n_117),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_147),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_140),
.B(n_127),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_146),
.B(n_15),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_148),
.A2(n_152),
.B1(n_154),
.B2(n_110),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_131),
.C(n_130),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_114),
.B(n_112),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_156),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_147),
.C(n_141),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_133),
.C(n_114),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_148),
.Y(n_167)
);

AO221x1_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_114),
.B1(n_107),
.B2(n_86),
.C(n_74),
.Y(n_158)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_161),
.A2(n_152),
.B1(n_153),
.B2(n_24),
.Y(n_170)
);

AO221x1_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_107),
.B1(n_86),
.B2(n_110),
.C(n_61),
.Y(n_162)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_153),
.B(n_12),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_157),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_174),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_156),
.C(n_155),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_163),
.B(n_160),
.C(n_7),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_175),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_31),
.C(n_12),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_173),
.C(n_168),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_166),
.C(n_169),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_179),
.B(n_175),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_181),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_180),
.A2(n_177),
.B(n_178),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_171),
.B(n_13),
.Y(n_184)
);

AOI221xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_183),
.B1(n_13),
.B2(n_8),
.C(n_5),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_8),
.Y(n_186)
);


endmodule