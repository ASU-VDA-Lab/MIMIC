module real_aes_10109_n_360 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_360);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_360;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_1929;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1694;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1583;
wire n_1250;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_1926;
wire n_898;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1940;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1914;
wire n_724;
wire n_1648;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_676;
wire n_658;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_367;
wire n_1017;
wire n_1942;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1939;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1592;
wire n_1056;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_1672;
wire n_747;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1457;
wire n_465;
wire n_719;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1931;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_1049;
wire n_466;
wire n_1584;
wire n_1277;
wire n_559;
wire n_1950;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1257;
wire n_1082;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1647;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1352;
wire n_729;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
AOI221xp5_ASAP7_75t_L g1539 ( .A1(n_0), .A2(n_257), .B1(n_836), .B2(n_903), .C(n_1141), .Y(n_1539) );
INVx1_ASAP7_75t_L g1552 ( .A(n_0), .Y(n_1552) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_1), .A2(n_108), .B1(n_451), .B2(n_459), .Y(n_450) );
INVx1_ASAP7_75t_L g552 ( .A(n_1), .Y(n_552) );
INVx1_ASAP7_75t_L g1717 ( .A(n_2), .Y(n_1717) );
OAI22xp5_ASAP7_75t_L g1500 ( .A1(n_3), .A2(n_321), .B1(n_678), .B2(n_681), .Y(n_1500) );
INVx1_ASAP7_75t_L g1520 ( .A(n_3), .Y(n_1520) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_4), .A2(n_222), .B1(n_902), .B2(n_903), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_4), .A2(n_222), .B1(n_918), .B2(n_920), .Y(n_917) );
AOI221xp5_ASAP7_75t_L g1646 ( .A1(n_5), .A2(n_213), .B1(n_713), .B2(n_714), .C(n_836), .Y(n_1646) );
OAI22xp33_ASAP7_75t_L g1651 ( .A1(n_5), .A2(n_324), .B1(n_681), .B2(n_1104), .Y(n_1651) );
INVx1_ASAP7_75t_L g700 ( .A(n_6), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_6), .A2(n_116), .B1(n_733), .B2(n_734), .Y(n_732) );
AOI221xp5_ASAP7_75t_L g1390 ( .A1(n_7), .A2(n_34), .B1(n_1391), .B2(n_1392), .C(n_1394), .Y(n_1390) );
INVx1_ASAP7_75t_L g1429 ( .A(n_7), .Y(n_1429) );
OAI22xp33_ASAP7_75t_L g618 ( .A1(n_8), .A2(n_107), .B1(n_619), .B2(n_621), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g639 ( .A1(n_8), .A2(n_107), .B1(n_628), .B2(n_640), .C(n_642), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g1295 ( .A1(n_9), .A2(n_21), .B1(n_1293), .B2(n_1296), .Y(n_1295) );
INVxp67_ASAP7_75t_SL g1301 ( .A(n_9), .Y(n_1301) );
AOI221xp5_ASAP7_75t_L g1608 ( .A1(n_10), .A2(n_284), .B1(n_593), .B2(n_596), .C(n_1174), .Y(n_1608) );
OAI22xp33_ASAP7_75t_L g1614 ( .A1(n_10), .A2(n_114), .B1(n_1106), .B2(n_1108), .Y(n_1614) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_11), .A2(n_123), .B1(n_716), .B2(n_718), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g726 ( .A1(n_11), .A2(n_123), .B1(n_727), .B2(n_728), .Y(n_726) );
AOI221xp5_ASAP7_75t_L g850 ( .A1(n_12), .A2(n_310), .B1(n_530), .B2(n_596), .C(n_703), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_12), .A2(n_310), .B1(n_733), .B2(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g1925 ( .A(n_13), .Y(n_1925) );
AOI22xp33_ASAP7_75t_SL g1938 ( .A1(n_13), .A2(n_300), .B1(n_730), .B2(n_1939), .Y(n_1938) );
INVx1_ASAP7_75t_L g1495 ( .A(n_14), .Y(n_1495) );
AO221x2_ASAP7_75t_L g1715 ( .A1(n_15), .A2(n_293), .B1(n_1672), .B2(n_1694), .C(n_1716), .Y(n_1715) );
OAI22xp33_ASAP7_75t_L g1005 ( .A1(n_16), .A2(n_79), .B1(n_451), .B2(n_459), .Y(n_1005) );
OAI22xp33_ASAP7_75t_L g1010 ( .A1(n_16), .A2(n_197), .B1(n_376), .B2(n_698), .Y(n_1010) );
AOI22xp33_ASAP7_75t_SL g1281 ( .A1(n_17), .A2(n_40), .B1(n_703), .B2(n_1282), .Y(n_1281) );
AOI22xp33_ASAP7_75t_L g1292 ( .A1(n_17), .A2(n_40), .B1(n_1293), .B2(n_1294), .Y(n_1292) );
CKINVDCx20_ASAP7_75t_R g1340 ( .A(n_18), .Y(n_1340) );
AO22x2_ASAP7_75t_L g880 ( .A1(n_19), .A2(n_881), .B1(n_941), .B2(n_942), .Y(n_880) );
INVxp67_ASAP7_75t_SL g941 ( .A(n_19), .Y(n_941) );
CKINVDCx16_ASAP7_75t_R g1534 ( .A(n_20), .Y(n_1534) );
INVxp33_ASAP7_75t_L g1307 ( .A(n_21), .Y(n_1307) );
CKINVDCx5p33_ASAP7_75t_R g1130 ( .A(n_22), .Y(n_1130) );
INVx1_ASAP7_75t_L g1168 ( .A(n_23), .Y(n_1168) );
AOI221xp5_ASAP7_75t_L g1228 ( .A1(n_23), .A2(n_232), .B1(n_923), .B2(n_1229), .C(n_1231), .Y(n_1228) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_24), .A2(n_95), .B1(n_925), .B2(n_998), .Y(n_1120) );
INVx1_ASAP7_75t_L g1148 ( .A(n_24), .Y(n_1148) );
XNOR2xp5_ASAP7_75t_L g1319 ( .A(n_25), .B(n_1320), .Y(n_1319) );
AOI22xp33_ASAP7_75t_SL g719 ( .A1(n_26), .A2(n_102), .B1(n_716), .B2(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_SL g754 ( .A(n_26), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g1626 ( .A1(n_27), .A2(n_358), .B1(n_927), .B2(n_1029), .Y(n_1626) );
INVxp67_ASAP7_75t_SL g1641 ( .A(n_27), .Y(n_1641) );
AOI22xp33_ASAP7_75t_L g1380 ( .A1(n_28), .A2(n_140), .B1(n_1381), .B2(n_1382), .Y(n_1380) );
INVx1_ASAP7_75t_L g1408 ( .A(n_28), .Y(n_1408) );
INVx1_ASAP7_75t_L g1002 ( .A(n_29), .Y(n_1002) );
OAI222xp33_ASAP7_75t_L g1008 ( .A1(n_29), .A2(n_244), .B1(n_335), .B2(n_590), .C1(n_934), .C2(n_1009), .Y(n_1008) );
CKINVDCx5p33_ASAP7_75t_R g1384 ( .A(n_30), .Y(n_1384) );
AOI22xp33_ASAP7_75t_SL g963 ( .A1(n_31), .A2(n_137), .B1(n_964), .B2(n_965), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_31), .A2(n_137), .B1(n_972), .B2(n_973), .Y(n_971) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_32), .A2(n_220), .B1(n_657), .B2(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1082 ( .A(n_32), .Y(n_1082) );
INVx1_ASAP7_75t_L g1544 ( .A(n_33), .Y(n_1544) );
AOI22xp33_ASAP7_75t_SL g1574 ( .A1(n_33), .A2(n_314), .B1(n_923), .B2(n_1022), .Y(n_1574) );
INVx1_ASAP7_75t_L g1424 ( .A(n_34), .Y(n_1424) );
AOI22xp33_ASAP7_75t_L g1538 ( .A1(n_35), .A2(n_81), .B1(n_972), .B2(n_1284), .Y(n_1538) );
INVx1_ASAP7_75t_L g1555 ( .A(n_35), .Y(n_1555) );
AOI221xp5_ASAP7_75t_L g832 ( .A1(n_36), .A2(n_214), .B1(n_833), .B2(n_834), .C(n_836), .Y(n_832) );
INVx1_ASAP7_75t_L g868 ( .A(n_36), .Y(n_868) );
INVx1_ASAP7_75t_L g950 ( .A(n_37), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_37), .A2(n_337), .B1(n_703), .B2(n_713), .Y(n_969) );
INVx1_ASAP7_75t_L g1540 ( .A(n_38), .Y(n_1540) );
AOI22xp33_ASAP7_75t_L g1572 ( .A1(n_38), .A2(n_178), .B1(n_1569), .B2(n_1573), .Y(n_1572) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_39), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g550 ( .A(n_39), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g1909 ( .A(n_41), .Y(n_1909) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_42), .A2(n_273), .B1(n_905), .B2(n_906), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_42), .A2(n_273), .B1(n_802), .B2(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g367 ( .A(n_43), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g1541 ( .A1(n_44), .A2(n_122), .B1(n_840), .B2(n_844), .Y(n_1541) );
INVx1_ASAP7_75t_L g1565 ( .A(n_44), .Y(n_1565) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_45), .A2(n_124), .B1(n_441), .B2(n_1004), .Y(n_1003) );
AOI22xp33_ASAP7_75t_SL g1017 ( .A1(n_45), .A2(n_124), .B1(n_968), .B2(n_972), .Y(n_1017) );
CKINVDCx5p33_ASAP7_75t_R g1217 ( .A(n_46), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_47), .A2(n_168), .B1(n_830), .B2(n_831), .Y(n_829) );
INVx1_ASAP7_75t_L g869 ( .A(n_47), .Y(n_869) );
CKINVDCx5p33_ASAP7_75t_R g1205 ( .A(n_48), .Y(n_1205) );
XOR2xp5_ASAP7_75t_L g1491 ( .A(n_49), .B(n_1492), .Y(n_1491) );
INVxp67_ASAP7_75t_SL g704 ( .A(n_50), .Y(n_704) );
OAI22xp33_ASAP7_75t_L g742 ( .A1(n_50), .A2(n_191), .B1(n_743), .B2(n_746), .Y(n_742) );
INVx1_ASAP7_75t_L g762 ( .A(n_51), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_51), .A2(n_231), .B1(n_713), .B2(n_793), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_52), .A2(n_306), .B1(n_927), .B2(n_1029), .Y(n_1050) );
INVx1_ASAP7_75t_L g1096 ( .A(n_52), .Y(n_1096) );
INVx1_ASAP7_75t_L g1012 ( .A(n_53), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_53), .A2(n_240), .B1(n_927), .B2(n_1029), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_54), .A2(n_157), .B1(n_792), .B2(n_793), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_54), .A2(n_157), .B1(n_628), .B2(n_730), .Y(n_804) );
AOI22x1_ASAP7_75t_SL g992 ( .A1(n_55), .A2(n_993), .B1(n_1030), .B2(n_1031), .Y(n_992) );
INVx1_ASAP7_75t_L g1030 ( .A(n_55), .Y(n_1030) );
INVx1_ASAP7_75t_L g1132 ( .A(n_56), .Y(n_1132) );
INVx1_ASAP7_75t_L g1370 ( .A(n_57), .Y(n_1370) );
INVx1_ASAP7_75t_L g1591 ( .A(n_58), .Y(n_1591) );
OAI221xp5_ASAP7_75t_L g1597 ( .A1(n_58), .A2(n_619), .B1(n_854), .B2(n_1598), .C(n_1602), .Y(n_1597) );
INVx1_ASAP7_75t_L g1451 ( .A(n_59), .Y(n_1451) );
OAI221xp5_ASAP7_75t_L g1470 ( .A1(n_59), .A2(n_621), .B1(n_1471), .B2(n_1475), .C(n_1479), .Y(n_1470) );
INVx1_ASAP7_75t_L g1129 ( .A(n_60), .Y(n_1129) );
AOI221xp5_ASAP7_75t_L g1140 ( .A1(n_60), .A2(n_212), .B1(n_723), .B2(n_1077), .C(n_1141), .Y(n_1140) );
AOI22xp5_ASAP7_75t_L g1730 ( .A1(n_61), .A2(n_336), .B1(n_1672), .B2(n_1694), .Y(n_1730) );
AOI22xp33_ASAP7_75t_L g1276 ( .A1(n_62), .A2(n_72), .B1(n_1277), .B2(n_1279), .Y(n_1276) );
AOI22xp33_ASAP7_75t_L g1287 ( .A1(n_62), .A2(n_72), .B1(n_1288), .B2(n_1290), .Y(n_1287) );
INVx1_ASAP7_75t_L g1511 ( .A(n_63), .Y(n_1511) );
AOI22xp33_ASAP7_75t_L g1525 ( .A1(n_63), .A2(n_242), .B1(n_918), .B2(n_1526), .Y(n_1525) );
INVx1_ASAP7_75t_L g1625 ( .A(n_64), .Y(n_1625) );
INVx1_ASAP7_75t_L g958 ( .A(n_65), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_65), .A2(n_195), .B1(n_716), .B2(n_968), .Y(n_967) );
INVx1_ASAP7_75t_L g1198 ( .A(n_66), .Y(n_1198) );
AOI221xp5_ASAP7_75t_L g1240 ( .A1(n_66), .A2(n_183), .B1(n_923), .B2(n_1241), .C(n_1243), .Y(n_1240) );
INVx1_ASAP7_75t_L g1358 ( .A(n_67), .Y(n_1358) );
OAI22xp33_ASAP7_75t_L g1365 ( .A1(n_67), .A2(n_138), .B1(n_681), .B2(n_1104), .Y(n_1365) );
AOI22xp33_ASAP7_75t_L g1548 ( .A1(n_68), .A2(n_247), .B1(n_905), .B2(n_906), .Y(n_1548) );
AOI22xp33_ASAP7_75t_L g1567 ( .A1(n_68), .A2(n_247), .B1(n_802), .B2(n_1391), .Y(n_1567) );
INVxp33_ASAP7_75t_L g1265 ( .A(n_69), .Y(n_1265) );
AOI22xp33_ASAP7_75t_SL g1283 ( .A1(n_69), .A2(n_147), .B1(n_1277), .B2(n_1284), .Y(n_1283) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_70), .A2(n_347), .B1(n_1061), .B2(n_1063), .Y(n_1060) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_70), .A2(n_347), .B1(n_1099), .B2(n_1100), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1326 ( .A1(n_71), .A2(n_359), .B1(n_927), .B2(n_1327), .Y(n_1326) );
INVx1_ASAP7_75t_L g1346 ( .A(n_71), .Y(n_1346) );
INVx1_ASAP7_75t_L g1506 ( .A(n_73), .Y(n_1506) );
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_73), .A2(n_208), .B1(n_1327), .B2(n_1528), .Y(n_1527) );
INVx1_ASAP7_75t_L g579 ( .A(n_74), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_74), .A2(n_266), .B1(n_628), .B2(n_630), .C(n_633), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_75), .B(n_822), .Y(n_821) );
OAI22xp33_ASAP7_75t_L g1905 ( .A1(n_76), .A2(n_326), .B1(n_1099), .B2(n_1100), .Y(n_1905) );
AOI22xp33_ASAP7_75t_L g1941 ( .A1(n_76), .A2(n_326), .B1(n_501), .B2(n_728), .Y(n_1941) );
INVx1_ASAP7_75t_L g1059 ( .A(n_77), .Y(n_1059) );
OAI211xp5_ASAP7_75t_SL g1068 ( .A1(n_77), .A2(n_621), .B(n_1069), .C(n_1078), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_78), .A2(n_207), .B1(n_716), .B2(n_790), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_78), .A2(n_207), .B1(n_727), .B2(n_802), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_79), .A2(n_152), .B1(n_793), .B2(n_902), .Y(n_1018) );
CKINVDCx5p33_ASAP7_75t_R g1445 ( .A(n_80), .Y(n_1445) );
INVx1_ASAP7_75t_L g1553 ( .A(n_81), .Y(n_1553) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_82), .A2(n_309), .B1(n_666), .B2(n_1024), .Y(n_1121) );
OAI221xp5_ASAP7_75t_L g1145 ( .A1(n_82), .A2(n_619), .B1(n_1097), .B2(n_1146), .C(n_1152), .Y(n_1145) );
INVx1_ASAP7_75t_L g1264 ( .A(n_83), .Y(n_1264) );
INVx1_ASAP7_75t_L g1502 ( .A(n_84), .Y(n_1502) );
AOI22xp33_ASAP7_75t_SL g1015 ( .A1(n_85), .A2(n_161), .B1(n_596), .B2(n_793), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_85), .A2(n_161), .B1(n_925), .B2(n_1024), .Y(n_1023) );
CKINVDCx5p33_ASAP7_75t_R g1399 ( .A(n_86), .Y(n_1399) );
CKINVDCx5p33_ASAP7_75t_R g1049 ( .A(n_87), .Y(n_1049) );
CKINVDCx5p33_ASAP7_75t_R g1207 ( .A(n_88), .Y(n_1207) );
OAI22xp5_ASAP7_75t_L g1385 ( .A1(n_89), .A2(n_261), .B1(n_1386), .B2(n_1387), .Y(n_1385) );
OAI221xp5_ASAP7_75t_L g1415 ( .A1(n_89), .A2(n_261), .B1(n_1186), .B2(n_1188), .C(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1472 ( .A(n_90), .Y(n_1472) );
OAI22xp33_ASAP7_75t_L g1485 ( .A1(n_90), .A2(n_181), .B1(n_678), .B2(n_681), .Y(n_1485) );
INVx1_ASAP7_75t_L g763 ( .A(n_91), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_91), .A2(n_179), .B1(n_716), .B2(n_797), .Y(n_796) );
XNOR2xp5_ASAP7_75t_L g1957 ( .A(n_92), .B(n_1958), .Y(n_1957) );
CKINVDCx5p33_ASAP7_75t_R g1126 ( .A(n_93), .Y(n_1126) );
CKINVDCx5p33_ASAP7_75t_R g1325 ( .A(n_94), .Y(n_1325) );
INVx1_ASAP7_75t_L g1151 ( .A(n_95), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_96), .A2(n_268), .B1(n_802), .B2(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g936 ( .A(n_96), .Y(n_936) );
INVx1_ASAP7_75t_L g890 ( .A(n_97), .Y(n_890) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_97), .A2(n_205), .B1(n_933), .B2(n_934), .Y(n_932) );
CKINVDCx20_ASAP7_75t_R g1620 ( .A(n_98), .Y(n_1620) );
XNOR2x2_ASAP7_75t_L g567 ( .A(n_99), .B(n_568), .Y(n_567) );
INVxp67_ASAP7_75t_SL g692 ( .A(n_100), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_100), .A2(n_274), .B1(n_727), .B2(n_737), .Y(n_736) );
CKINVDCx5p33_ASAP7_75t_R g595 ( .A(n_101), .Y(n_595) );
INVxp33_ASAP7_75t_L g753 ( .A(n_102), .Y(n_753) );
BUFx2_ASAP7_75t_L g393 ( .A(n_103), .Y(n_393) );
BUFx2_ASAP7_75t_L g491 ( .A(n_103), .Y(n_491) );
INVx1_ASAP7_75t_L g562 ( .A(n_103), .Y(n_562) );
OR2x2_ASAP7_75t_L g1185 ( .A(n_103), .B(n_606), .Y(n_1185) );
AOI22xp33_ASAP7_75t_SL g1016 ( .A1(n_104), .A2(n_250), .B1(n_905), .B2(n_968), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_104), .A2(n_250), .B1(n_1021), .B2(n_1022), .Y(n_1020) );
INVx1_ASAP7_75t_L g1073 ( .A(n_105), .Y(n_1073) );
OAI22xp5_ASAP7_75t_L g1105 ( .A1(n_105), .A2(n_203), .B1(n_1106), .B2(n_1108), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_106), .A2(n_343), .B1(n_628), .B2(n_730), .Y(n_962) );
AOI22xp33_ASAP7_75t_SL g974 ( .A1(n_106), .A2(n_343), .B1(n_713), .B2(n_975), .Y(n_974) );
INVx1_ASAP7_75t_L g430 ( .A(n_108), .Y(n_430) );
INVx1_ASAP7_75t_L g1476 ( .A(n_109), .Y(n_1476) );
OAI22xp33_ASAP7_75t_L g1486 ( .A1(n_109), .A2(n_209), .B1(n_1106), .B2(n_1108), .Y(n_1486) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_110), .A2(n_170), .B1(n_746), .B2(n_953), .Y(n_952) );
OAI22xp33_ASAP7_75t_L g985 ( .A1(n_110), .A2(n_170), .B1(n_706), .B2(n_986), .Y(n_985) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_111), .Y(n_577) );
INVx1_ASAP7_75t_L g1455 ( .A(n_112), .Y(n_1455) );
OAI22xp5_ASAP7_75t_L g1462 ( .A1(n_112), .A2(n_117), .B1(n_608), .B2(n_614), .Y(n_1462) );
AOI221xp5_ASAP7_75t_L g1546 ( .A1(n_113), .A2(n_198), .B1(n_530), .B2(n_701), .C(n_1547), .Y(n_1546) );
AOI22xp33_ASAP7_75t_L g1568 ( .A1(n_113), .A2(n_198), .B1(n_998), .B2(n_1569), .Y(n_1568) );
INVx1_ASAP7_75t_L g1606 ( .A(n_114), .Y(n_1606) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_115), .A2(n_217), .B1(n_713), .B2(n_722), .Y(n_721) );
INVxp67_ASAP7_75t_SL g741 ( .A(n_115), .Y(n_741) );
INVxp33_ASAP7_75t_L g695 ( .A(n_116), .Y(n_695) );
INVx1_ASAP7_75t_L g1454 ( .A(n_117), .Y(n_1454) );
OAI221xp5_ASAP7_75t_L g1504 ( .A1(n_118), .A2(n_619), .B1(n_854), .B2(n_1505), .C(n_1509), .Y(n_1504) );
AOI22xp33_ASAP7_75t_SL g1529 ( .A1(n_118), .A2(n_282), .B1(n_925), .B2(n_1024), .Y(n_1529) );
AOI22xp33_ASAP7_75t_L g1396 ( .A1(n_119), .A2(n_288), .B1(n_925), .B2(n_1397), .Y(n_1396) );
INVx1_ASAP7_75t_L g1430 ( .A(n_119), .Y(n_1430) );
AOI221xp5_ASAP7_75t_L g1076 ( .A1(n_120), .A2(n_203), .B1(n_713), .B2(n_722), .C(n_1077), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g1103 ( .A1(n_120), .A2(n_252), .B1(n_681), .B2(n_1104), .Y(n_1103) );
INVxp67_ASAP7_75t_SL g1267 ( .A(n_121), .Y(n_1267) );
AOI22xp33_ASAP7_75t_SL g1285 ( .A1(n_121), .A2(n_225), .B1(n_903), .B2(n_1282), .Y(n_1285) );
INVx1_ASAP7_75t_L g1564 ( .A(n_122), .Y(n_1564) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_125), .A2(n_228), .B1(n_927), .B2(n_1029), .Y(n_1298) );
INVxp33_ASAP7_75t_SL g1304 ( .A(n_125), .Y(n_1304) );
CKINVDCx16_ASAP7_75t_R g1727 ( .A(n_126), .Y(n_1727) );
CKINVDCx5p33_ASAP7_75t_R g1116 ( .A(n_127), .Y(n_1116) );
CKINVDCx5p33_ASAP7_75t_R g1115 ( .A(n_128), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_129), .A2(n_155), .B1(n_1021), .B2(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1153 ( .A(n_129), .Y(n_1153) );
OAI22xp33_ASAP7_75t_L g1337 ( .A1(n_130), .A2(n_206), .B1(n_657), .B2(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g1363 ( .A(n_130), .Y(n_1363) );
INVx1_ASAP7_75t_L g1448 ( .A(n_131), .Y(n_1448) );
CKINVDCx5p33_ASAP7_75t_R g1587 ( .A(n_132), .Y(n_1587) );
OA22x2_ASAP7_75t_L g390 ( .A1(n_133), .A2(n_391), .B1(n_565), .B2(n_566), .Y(n_390) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_133), .Y(n_566) );
INVx1_ASAP7_75t_L g1644 ( .A(n_134), .Y(n_1644) );
OAI22xp33_ASAP7_75t_L g1652 ( .A1(n_134), .A2(n_213), .B1(n_1106), .B2(n_1108), .Y(n_1652) );
AOI22xp5_ASAP7_75t_L g1714 ( .A1(n_135), .A2(n_331), .B1(n_1672), .B2(n_1694), .Y(n_1714) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_136), .A2(n_176), .B1(n_920), .B2(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g939 ( .A(n_136), .Y(n_939) );
AOI221xp5_ASAP7_75t_L g1359 ( .A1(n_138), .A2(n_315), .B1(n_593), .B2(n_713), .C(n_714), .Y(n_1359) );
CKINVDCx5p33_ASAP7_75t_R g1914 ( .A(n_139), .Y(n_1914) );
INVx1_ASAP7_75t_L g1413 ( .A(n_140), .Y(n_1413) );
INVx1_ASAP7_75t_L g1628 ( .A(n_141), .Y(n_1628) );
OAI221xp5_ASAP7_75t_L g1634 ( .A1(n_141), .A2(n_619), .B1(n_1097), .B2(n_1635), .C(n_1639), .Y(n_1634) );
INVx1_ASAP7_75t_L g1499 ( .A(n_142), .Y(n_1499) );
INVx1_ASAP7_75t_L g781 ( .A(n_143), .Y(n_781) );
AOI22xp33_ASAP7_75t_SL g809 ( .A1(n_143), .A2(n_323), .B1(n_628), .B2(n_810), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_144), .A2(n_171), .B1(n_980), .B2(n_981), .Y(n_979) );
INVx1_ASAP7_75t_L g988 ( .A(n_144), .Y(n_988) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_145), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g1703 ( .A1(n_146), .A2(n_150), .B1(n_1704), .B2(n_1707), .Y(n_1703) );
INVxp33_ASAP7_75t_SL g1262 ( .A(n_147), .Y(n_1262) );
OAI22xp5_ASAP7_75t_L g1522 ( .A1(n_148), .A2(n_303), .B1(n_1099), .B2(n_1100), .Y(n_1522) );
AOI22xp33_ASAP7_75t_L g1530 ( .A1(n_148), .A2(n_303), .B1(n_1063), .B2(n_1531), .Y(n_1530) );
INVx1_ASAP7_75t_L g1923 ( .A(n_149), .Y(n_1923) );
AOI22xp33_ASAP7_75t_L g1936 ( .A1(n_149), .A2(n_304), .B1(n_964), .B2(n_1937), .Y(n_1936) );
INVx1_ASAP7_75t_L g1357 ( .A(n_151), .Y(n_1357) );
OAI22xp33_ASAP7_75t_L g1366 ( .A1(n_151), .A2(n_315), .B1(n_1106), .B2(n_1108), .Y(n_1366) );
INVx1_ASAP7_75t_L g997 ( .A(n_152), .Y(n_997) );
AOI22xp5_ASAP7_75t_L g1709 ( .A1(n_153), .A2(n_341), .B1(n_1664), .B2(n_1710), .Y(n_1709) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_154), .Y(n_431) );
INVx1_ASAP7_75t_L g1155 ( .A(n_155), .Y(n_1155) );
AO221x2_ASAP7_75t_L g1738 ( .A1(n_156), .A2(n_227), .B1(n_1664), .B2(n_1672), .C(n_1739), .Y(n_1738) );
INVx1_ASAP7_75t_L g1669 ( .A(n_158), .Y(n_1669) );
INVx1_ASAP7_75t_L g1670 ( .A(n_159), .Y(n_1670) );
OAI22xp33_ASAP7_75t_L g1594 ( .A1(n_160), .A2(n_338), .B1(n_1457), .B2(n_1458), .Y(n_1594) );
INVx1_ASAP7_75t_L g1610 ( .A(n_160), .Y(n_1610) );
AOI22xp5_ASAP7_75t_L g1729 ( .A1(n_162), .A2(n_349), .B1(n_1704), .B2(n_1707), .Y(n_1729) );
INVx1_ASAP7_75t_L g776 ( .A(n_163), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_163), .A2(n_204), .B1(n_673), .B2(n_802), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g1588 ( .A1(n_164), .A2(n_356), .B1(n_1062), .B2(n_1589), .Y(n_1588) );
INVx1_ASAP7_75t_L g1599 ( .A(n_164), .Y(n_1599) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_165), .A2(n_296), .B1(n_927), .B2(n_1029), .Y(n_1122) );
OAI22xp5_ASAP7_75t_L g1157 ( .A1(n_165), .A2(n_296), .B1(n_614), .B2(n_1099), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_166), .A2(n_318), .B1(n_830), .B2(n_852), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_166), .A2(n_318), .B1(n_635), .B2(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g1930 ( .A(n_167), .Y(n_1930) );
INVx1_ASAP7_75t_L g865 ( .A(n_168), .Y(n_865) );
INVx1_ASAP7_75t_L g696 ( .A(n_169), .Y(n_696) );
INVx1_ASAP7_75t_L g989 ( .A(n_171), .Y(n_989) );
INVx1_ASAP7_75t_L g1667 ( .A(n_172), .Y(n_1667) );
NAND2xp5_ASAP7_75t_L g1686 ( .A(n_172), .B(n_1680), .Y(n_1686) );
INVx1_ASAP7_75t_L g1268 ( .A(n_173), .Y(n_1268) );
OAI22xp5_ASAP7_75t_L g1302 ( .A1(n_173), .A2(n_352), .B1(n_706), .B2(n_934), .Y(n_1302) );
INVx1_ASAP7_75t_L g1592 ( .A(n_174), .Y(n_1592) );
OAI211xp5_ASAP7_75t_SL g1604 ( .A1(n_174), .A2(n_621), .B(n_1605), .C(n_1609), .Y(n_1604) );
INVx1_ASAP7_75t_L g886 ( .A(n_175), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_175), .A2(n_201), .B1(n_910), .B2(n_913), .Y(n_909) );
INVx1_ASAP7_75t_L g931 ( .A(n_176), .Y(n_931) );
INVx2_ASAP7_75t_L g379 ( .A(n_177), .Y(n_379) );
INVx1_ASAP7_75t_L g1549 ( .A(n_178), .Y(n_1549) );
INVx1_ASAP7_75t_L g766 ( .A(n_179), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g1631 ( .A1(n_180), .A2(n_219), .B1(n_1041), .B2(n_1458), .Y(n_1631) );
INVx1_ASAP7_75t_L g1648 ( .A(n_180), .Y(n_1648) );
INVx1_ASAP7_75t_L g1477 ( .A(n_181), .Y(n_1477) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_182), .Y(n_503) );
INVx1_ASAP7_75t_L g1200 ( .A(n_183), .Y(n_1200) );
AOI22xp33_ASAP7_75t_L g1334 ( .A1(n_184), .A2(n_353), .B1(n_802), .B2(n_1335), .Y(n_1334) );
OAI22xp5_ASAP7_75t_L g1342 ( .A1(n_184), .A2(n_353), .B1(n_1099), .B2(n_1100), .Y(n_1342) );
INVx1_ASAP7_75t_L g449 ( .A(n_185), .Y(n_449) );
BUFx3_ASAP7_75t_L g465 ( .A(n_185), .Y(n_465) );
INVx1_ASAP7_75t_L g1202 ( .A(n_186), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_186), .A2(n_215), .B1(n_859), .B2(n_1245), .Y(n_1244) );
INVx1_ASAP7_75t_L g1607 ( .A(n_187), .Y(n_1607) );
OAI22xp33_ASAP7_75t_L g1613 ( .A1(n_187), .A2(n_284), .B1(n_681), .B2(n_1104), .Y(n_1613) );
INVx1_ASAP7_75t_L g849 ( .A(n_188), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_188), .A2(n_278), .B1(n_661), .B2(n_666), .Y(n_862) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_189), .Y(n_477) );
INVx1_ASAP7_75t_L g1740 ( .A(n_190), .Y(n_1740) );
INVx1_ASAP7_75t_L g707 ( .A(n_191), .Y(n_707) );
CKINVDCx5p33_ASAP7_75t_R g438 ( .A(n_192), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g1176 ( .A(n_193), .Y(n_1176) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_194), .A2(n_328), .B1(n_608), .B2(n_614), .Y(n_607) );
INVx1_ASAP7_75t_L g646 ( .A(n_194), .Y(n_646) );
INVx1_ASAP7_75t_L g959 ( .A(n_195), .Y(n_959) );
OAI221xp5_ASAP7_75t_L g767 ( .A1(n_196), .A2(n_265), .B1(n_746), .B2(n_768), .C(n_769), .Y(n_767) );
INVx1_ASAP7_75t_L g779 ( .A(n_196), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_197), .A2(n_244), .B1(n_1026), .B2(n_1027), .Y(n_1025) );
INVx1_ASAP7_75t_L g1629 ( .A(n_199), .Y(n_1629) );
OAI211xp5_ASAP7_75t_SL g1642 ( .A1(n_199), .A2(n_621), .B(n_1643), .C(n_1647), .Y(n_1642) );
XNOR2xp5_ASAP7_75t_L g1110 ( .A(n_200), .B(n_1111), .Y(n_1110) );
INVx1_ASAP7_75t_L g1662 ( .A(n_200), .Y(n_1662) );
INVx1_ASAP7_75t_L g896 ( .A(n_201), .Y(n_896) );
AOI221xp5_ASAP7_75t_L g1376 ( .A1(n_202), .A2(n_216), .B1(n_1377), .B2(n_1378), .C(n_1379), .Y(n_1376) );
INVx1_ASAP7_75t_L g1412 ( .A(n_202), .Y(n_1412) );
INVx1_ASAP7_75t_L g777 ( .A(n_204), .Y(n_777) );
INVx1_ASAP7_75t_L g893 ( .A(n_205), .Y(n_893) );
INVx1_ASAP7_75t_L g1361 ( .A(n_206), .Y(n_1361) );
INVx1_ASAP7_75t_L g1508 ( .A(n_208), .Y(n_1508) );
INVx1_ASAP7_75t_L g1473 ( .A(n_209), .Y(n_1473) );
INVx1_ASAP7_75t_L g1741 ( .A(n_210), .Y(n_1741) );
CKINVDCx5p33_ASAP7_75t_R g1910 ( .A(n_211), .Y(n_1910) );
INVx1_ASAP7_75t_L g1127 ( .A(n_212), .Y(n_1127) );
INVx1_ASAP7_75t_L g866 ( .A(n_214), .Y(n_866) );
INVx1_ASAP7_75t_L g1195 ( .A(n_215), .Y(n_1195) );
INVx1_ASAP7_75t_L g1410 ( .A(n_216), .Y(n_1410) );
INVxp33_ASAP7_75t_L g748 ( .A(n_217), .Y(n_748) );
INVx1_ASAP7_75t_L g489 ( .A(n_218), .Y(n_489) );
INVx1_ASAP7_75t_L g655 ( .A(n_218), .Y(n_655) );
INVx1_ASAP7_75t_L g1649 ( .A(n_219), .Y(n_1649) );
INVx1_ASAP7_75t_L g1079 ( .A(n_220), .Y(n_1079) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_221), .Y(n_508) );
INVx1_ASAP7_75t_L g1698 ( .A(n_223), .Y(n_1698) );
INVx1_ASAP7_75t_L g846 ( .A(n_224), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_224), .A2(n_270), .B1(n_635), .B2(n_803), .Y(n_863) );
INVxp33_ASAP7_75t_SL g1261 ( .A(n_225), .Y(n_1261) );
CKINVDCx5p33_ASAP7_75t_R g1916 ( .A(n_226), .Y(n_1916) );
XOR2x2_ASAP7_75t_L g1902 ( .A(n_227), .B(n_1903), .Y(n_1902) );
AOI22xp33_ASAP7_75t_L g1952 ( .A1(n_227), .A2(n_1953), .B1(n_1956), .B2(n_1960), .Y(n_1952) );
INVxp67_ASAP7_75t_SL g1305 ( .A(n_228), .Y(n_1305) );
CKINVDCx5p33_ASAP7_75t_R g956 ( .A(n_229), .Y(n_956) );
CKINVDCx5p33_ASAP7_75t_R g885 ( .A(n_230), .Y(n_885) );
INVx1_ASAP7_75t_L g770 ( .A(n_231), .Y(n_770) );
INVx1_ASAP7_75t_L g1178 ( .A(n_232), .Y(n_1178) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_233), .Y(n_600) );
OAI221xp5_ASAP7_75t_L g647 ( .A1(n_233), .A2(n_648), .B1(n_656), .B2(n_657), .C(n_660), .Y(n_647) );
CKINVDCx5p33_ASAP7_75t_R g1209 ( .A(n_234), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_235), .A2(n_259), .B1(n_840), .B2(n_844), .Y(n_839) );
INVx1_ASAP7_75t_L g874 ( .A(n_235), .Y(n_874) );
INVx1_ASAP7_75t_L g1460 ( .A(n_236), .Y(n_1460) );
AOI22xp5_ASAP7_75t_L g1713 ( .A1(n_237), .A2(n_311), .B1(n_1704), .B2(n_1707), .Y(n_1713) );
INVx1_ASAP7_75t_L g1498 ( .A(n_238), .Y(n_1498) );
INVx1_ASAP7_75t_L g878 ( .A(n_239), .Y(n_878) );
INVx1_ASAP7_75t_L g1013 ( .A(n_240), .Y(n_1013) );
CKINVDCx5p33_ASAP7_75t_R g1913 ( .A(n_241), .Y(n_1913) );
INVx1_ASAP7_75t_L g1510 ( .A(n_242), .Y(n_1510) );
CKINVDCx5p33_ASAP7_75t_R g1172 ( .A(n_243), .Y(n_1172) );
CKINVDCx5p33_ASAP7_75t_R g765 ( .A(n_245), .Y(n_765) );
OAI22xp33_ASAP7_75t_L g1456 ( .A1(n_246), .A2(n_333), .B1(n_1457), .B2(n_1458), .Y(n_1456) );
INVx1_ASAP7_75t_L g1481 ( .A(n_246), .Y(n_1481) );
INVx1_ASAP7_75t_L g1333 ( .A(n_248), .Y(n_1333) );
OAI211xp5_ASAP7_75t_SL g1354 ( .A1(n_248), .A2(n_621), .B(n_1355), .C(n_1360), .Y(n_1354) );
CKINVDCx16_ASAP7_75t_R g684 ( .A(n_249), .Y(n_684) );
INVx1_ASAP7_75t_L g1066 ( .A(n_251), .Y(n_1066) );
INVx1_ASAP7_75t_L g1075 ( .A(n_252), .Y(n_1075) );
INVx1_ASAP7_75t_L g1581 ( .A(n_253), .Y(n_1581) );
INVx1_ASAP7_75t_L g1330 ( .A(n_254), .Y(n_1330) );
OAI221xp5_ASAP7_75t_L g1343 ( .A1(n_254), .A2(n_619), .B1(n_854), .B2(n_1344), .C(n_1351), .Y(n_1343) );
CKINVDCx5p33_ASAP7_75t_R g1048 ( .A(n_255), .Y(n_1048) );
INVx1_ASAP7_75t_L g1450 ( .A(n_256), .Y(n_1450) );
OAI221xp5_ASAP7_75t_L g1463 ( .A1(n_256), .A2(n_619), .B1(n_854), .B2(n_1464), .C(n_1469), .Y(n_1463) );
INVx1_ASAP7_75t_L g1556 ( .A(n_257), .Y(n_1556) );
XNOR2xp5_ASAP7_75t_L g1163 ( .A(n_258), .B(n_1164), .Y(n_1163) );
XNOR2x1_ASAP7_75t_L g1311 ( .A(n_258), .B(n_1164), .Y(n_1311) );
INVx1_ASAP7_75t_L g872 ( .A(n_259), .Y(n_872) );
INVx1_ASAP7_75t_L g895 ( .A(n_260), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_260), .A2(n_344), .B1(n_902), .B2(n_903), .Y(n_914) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_262), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_263), .A2(n_286), .B1(n_398), .B2(n_406), .Y(n_397) );
INVx1_ASAP7_75t_L g522 ( .A(n_263), .Y(n_522) );
INVx1_ASAP7_75t_L g1585 ( .A(n_264), .Y(n_1585) );
AOI21xp33_ASAP7_75t_L g1603 ( .A1(n_264), .A2(n_530), .B(n_1143), .Y(n_1603) );
INVx1_ASAP7_75t_L g780 ( .A(n_265), .Y(n_780) );
AOI21xp33_ASAP7_75t_L g581 ( .A1(n_266), .A2(n_530), .B(n_582), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g1324 ( .A(n_267), .Y(n_1324) );
INVx1_ASAP7_75t_L g937 ( .A(n_268), .Y(n_937) );
OAI221xp5_ASAP7_75t_L g1906 ( .A1(n_269), .A2(n_621), .B1(n_1907), .B2(n_1911), .C(n_1915), .Y(n_1906) );
AOI22xp33_ASAP7_75t_SL g1940 ( .A1(n_269), .A2(n_334), .B1(n_640), .B2(n_1939), .Y(n_1940) );
INVx1_ASAP7_75t_L g847 ( .A(n_270), .Y(n_847) );
INVx1_ASAP7_75t_L g1403 ( .A(n_271), .Y(n_1403) );
OAI211xp5_ASAP7_75t_L g412 ( .A1(n_272), .A2(n_413), .B(n_418), .C(n_425), .Y(n_412) );
INVx1_ASAP7_75t_L g518 ( .A(n_272), .Y(n_518) );
INVx1_ASAP7_75t_L g690 ( .A(n_274), .Y(n_690) );
CKINVDCx5p33_ASAP7_75t_R g1401 ( .A(n_275), .Y(n_1401) );
XNOR2xp5_ASAP7_75t_L g1578 ( .A(n_276), .B(n_1579), .Y(n_1578) );
OAI221xp5_ASAP7_75t_L g1180 ( .A1(n_277), .A2(n_351), .B1(n_1181), .B2(n_1186), .C(n_1188), .Y(n_1180) );
OAI22xp5_ASAP7_75t_L g1222 ( .A1(n_277), .A2(n_351), .B1(n_1223), .B2(n_1226), .Y(n_1222) );
INVx1_ASAP7_75t_L g838 ( .A(n_278), .Y(n_838) );
INVx1_ASAP7_75t_L g1444 ( .A(n_279), .Y(n_1444) );
AOI22xp33_ASAP7_75t_SL g1593 ( .A1(n_280), .A2(n_305), .B1(n_737), .B2(n_1289), .Y(n_1593) );
OAI22xp5_ASAP7_75t_L g1596 ( .A1(n_280), .A2(n_305), .B1(n_1099), .B2(n_1100), .Y(n_1596) );
BUFx3_ASAP7_75t_L g448 ( .A(n_281), .Y(n_448) );
INVx1_ASAP7_75t_L g458 ( .A(n_281), .Y(n_458) );
OAI221xp5_ASAP7_75t_L g1512 ( .A1(n_282), .A2(n_621), .B1(n_1513), .B2(n_1515), .C(n_1521), .Y(n_1512) );
XNOR2xp5_ASAP7_75t_L g1036 ( .A(n_283), .B(n_1037), .Y(n_1036) );
AO22x2_ASAP7_75t_L g757 ( .A1(n_285), .A2(n_758), .B1(n_812), .B2(n_813), .Y(n_757) );
INVxp67_ASAP7_75t_L g812 ( .A(n_285), .Y(n_812) );
INVx1_ASAP7_75t_L g520 ( .A(n_286), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g1211 ( .A(n_287), .Y(n_1211) );
INVx1_ASAP7_75t_L g1422 ( .A(n_288), .Y(n_1422) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_289), .Y(n_375) );
INVx1_ASAP7_75t_L g564 ( .A(n_289), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_289), .B(n_339), .Y(n_606) );
AND2x2_ASAP7_75t_L g610 ( .A(n_289), .B(n_402), .Y(n_610) );
INVx1_ASAP7_75t_L g1681 ( .A(n_290), .Y(n_1681) );
AOI21xp33_ASAP7_75t_L g591 ( .A1(n_291), .A2(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g671 ( .A(n_291), .Y(n_671) );
AO22x2_ASAP7_75t_L g1256 ( .A1(n_292), .A2(n_1257), .B1(n_1258), .B2(n_1308), .Y(n_1256) );
INVxp67_ASAP7_75t_SL g1257 ( .A(n_292), .Y(n_1257) );
XNOR2xp5_ASAP7_75t_L g946 ( .A(n_293), .B(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g1699 ( .A(n_294), .Y(n_1699) );
INVx2_ASAP7_75t_L g445 ( .A(n_295), .Y(n_445) );
OR2x2_ASAP7_75t_L g670 ( .A(n_295), .B(n_655), .Y(n_670) );
INVx1_ASAP7_75t_L g1674 ( .A(n_297), .Y(n_1674) );
CKINVDCx5p33_ASAP7_75t_R g1402 ( .A(n_298), .Y(n_1402) );
CKINVDCx16_ASAP7_75t_R g1696 ( .A(n_299), .Y(n_1696) );
INVx1_ASAP7_75t_L g1928 ( .A(n_300), .Y(n_1928) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_301), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_302), .Y(n_499) );
INVx1_ASAP7_75t_L g1920 ( .A(n_304), .Y(n_1920) );
INVx1_ASAP7_75t_L g1092 ( .A(n_306), .Y(n_1092) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_307), .Y(n_585) );
INVx1_ASAP7_75t_L g1723 ( .A(n_308), .Y(n_1723) );
OAI211xp5_ASAP7_75t_SL g1134 ( .A1(n_309), .A2(n_621), .B(n_1135), .C(n_1144), .Y(n_1134) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_312), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_313), .A2(n_327), .B1(n_628), .B2(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g991 ( .A(n_313), .Y(n_991) );
INVx1_ASAP7_75t_L g1543 ( .A(n_314), .Y(n_1543) );
AOI22xp5_ASAP7_75t_L g1630 ( .A1(n_316), .A2(n_340), .B1(n_1063), .B2(n_1288), .Y(n_1630) );
OAI22xp5_ASAP7_75t_L g1633 ( .A1(n_316), .A2(n_340), .B1(n_608), .B2(n_614), .Y(n_1633) );
INVx1_ASAP7_75t_L g1617 ( .A(n_317), .Y(n_1617) );
INVx1_ASAP7_75t_L g1055 ( .A(n_319), .Y(n_1055) );
OAI221xp5_ASAP7_75t_L g1084 ( .A1(n_319), .A2(n_619), .B1(n_1085), .B2(n_1088), .C(n_1097), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_320), .A2(n_354), .B1(n_713), .B2(n_714), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_320), .A2(n_354), .B1(n_470), .B2(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g1514 ( .A(n_321), .Y(n_1514) );
INVx1_ASAP7_75t_L g1718 ( .A(n_322), .Y(n_1718) );
INVx1_ASAP7_75t_L g786 ( .A(n_323), .Y(n_786) );
INVx1_ASAP7_75t_L g1645 ( .A(n_324), .Y(n_1645) );
INVx1_ASAP7_75t_L g1496 ( .A(n_325), .Y(n_1496) );
INVx1_ASAP7_75t_L g984 ( .A(n_327), .Y(n_984) );
INVx1_ASAP7_75t_L g643 ( .A(n_328), .Y(n_643) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_329), .Y(n_369) );
AND3x2_ASAP7_75t_L g1668 ( .A(n_329), .B(n_367), .C(n_1669), .Y(n_1668) );
NAND2xp5_ASAP7_75t_L g1678 ( .A(n_329), .B(n_367), .Y(n_1678) );
INVx2_ASAP7_75t_L g380 ( .A(n_330), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g1447 ( .A(n_332), .Y(n_1447) );
INVx1_ASAP7_75t_L g1480 ( .A(n_333), .Y(n_1480) );
OAI221xp5_ASAP7_75t_L g1918 ( .A1(n_334), .A2(n_619), .B1(n_854), .B2(n_1919), .C(n_1924), .Y(n_1918) );
CKINVDCx5p33_ASAP7_75t_R g1001 ( .A(n_335), .Y(n_1001) );
XNOR2xp5_ASAP7_75t_L g1438 ( .A(n_336), .B(n_1439), .Y(n_1438) );
INVx1_ASAP7_75t_L g955 ( .A(n_337), .Y(n_955) );
INVx1_ASAP7_75t_L g1611 ( .A(n_338), .Y(n_1611) );
INVx1_ASAP7_75t_L g382 ( .A(n_339), .Y(n_382) );
INVx2_ASAP7_75t_L g402 ( .A(n_339), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_342), .Y(n_396) );
INVx1_ASAP7_75t_L g888 ( .A(n_344), .Y(n_888) );
INVx1_ASAP7_75t_L g599 ( .A(n_345), .Y(n_599) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_345), .Y(n_656) );
OAI211xp5_ASAP7_75t_L g467 ( .A1(n_346), .A2(n_468), .B(n_473), .C(n_484), .Y(n_467) );
INVx1_ASAP7_75t_L g557 ( .A(n_346), .Y(n_557) );
INVx1_ASAP7_75t_L g1724 ( .A(n_348), .Y(n_1724) );
NOR2xp33_ASAP7_75t_L g1557 ( .A(n_350), .B(n_1558), .Y(n_1557) );
INVx1_ASAP7_75t_L g1269 ( .A(n_352), .Y(n_1269) );
INVx1_ASAP7_75t_L g1624 ( .A(n_355), .Y(n_1624) );
INVx1_ASAP7_75t_L g1601 ( .A(n_356), .Y(n_1601) );
CKINVDCx5p33_ASAP7_75t_R g1917 ( .A(n_357), .Y(n_1917) );
INVxp33_ASAP7_75t_SL g1640 ( .A(n_358), .Y(n_1640) );
INVx1_ASAP7_75t_L g1350 ( .A(n_359), .Y(n_1350) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_383), .B(n_1656), .Y(n_360) );
BUFx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx3_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_365), .B(n_370), .Y(n_364) );
AND2x4_ASAP7_75t_L g1951 ( .A(n_365), .B(n_371), .Y(n_1951) );
NOR2xp33_ASAP7_75t_SL g365 ( .A(n_366), .B(n_368), .Y(n_365) );
INVx1_ASAP7_75t_SL g1955 ( .A(n_366), .Y(n_1955) );
NAND2xp5_ASAP7_75t_L g1965 ( .A(n_366), .B(n_368), .Y(n_1965) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g1954 ( .A(n_368), .B(n_1955), .Y(n_1954) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_372), .B(n_376), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g392 ( .A(n_373), .B(n_393), .Y(n_392) );
OR2x6_ASAP7_75t_L g687 ( .A(n_373), .B(n_393), .Y(n_687) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g711 ( .A(n_374), .B(n_382), .Y(n_711) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g530 ( .A(n_375), .B(n_401), .Y(n_530) );
INVx8_ASAP7_75t_L g395 ( .A(n_376), .Y(n_395) );
OR2x6_ASAP7_75t_L g376 ( .A(n_377), .B(n_381), .Y(n_376) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_377), .Y(n_532) );
OR2x6_ASAP7_75t_L g698 ( .A(n_377), .B(n_400), .Y(n_698) );
INVx1_ASAP7_75t_L g1150 ( .A(n_377), .Y(n_1150) );
INVx2_ASAP7_75t_SL g1194 ( .A(n_377), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1215 ( .A(n_377), .B(n_1185), .Y(n_1215) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx2_ASAP7_75t_L g405 ( .A(n_379), .Y(n_405) );
AND2x4_ASAP7_75t_L g410 ( .A(n_379), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g417 ( .A(n_379), .Y(n_417) );
INVx1_ASAP7_75t_L g424 ( .A(n_379), .Y(n_424) );
AND2x2_ASAP7_75t_L g429 ( .A(n_379), .B(n_380), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_380), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g411 ( .A(n_380), .Y(n_411) );
INVx1_ASAP7_75t_L g416 ( .A(n_380), .Y(n_416) );
INVx1_ASAP7_75t_L g433 ( .A(n_380), .Y(n_433) );
INVx1_ASAP7_75t_L g613 ( .A(n_380), .Y(n_613) );
AND2x4_ASAP7_75t_L g432 ( .A(n_381), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g934 ( .A(n_382), .B(n_436), .Y(n_934) );
OR2x2_ASAP7_75t_L g986 ( .A(n_382), .B(n_436), .Y(n_986) );
XNOR2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_1315), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_1033), .B1(n_1313), .B2(n_1314), .Y(n_384) );
INVx2_ASAP7_75t_L g1313 ( .A(n_385), .Y(n_1313) );
XNOR2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_815), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
XNOR2x1_ASAP7_75t_L g388 ( .A(n_389), .B(n_682), .Y(n_388) );
XNOR2x1_ASAP7_75t_L g389 ( .A(n_390), .B(n_567), .Y(n_389) );
INVx1_ASAP7_75t_L g565 ( .A(n_391), .Y(n_565) );
OAI211xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B(n_439), .C(n_492), .Y(n_391) );
AOI31xp33_ASAP7_75t_L g929 ( .A1(n_392), .A2(n_930), .A3(n_935), .B(n_938), .Y(n_929) );
AOI31xp33_ASAP7_75t_L g1299 ( .A1(n_392), .A2(n_1300), .A3(n_1303), .B(n_1306), .Y(n_1299) );
AND2x4_ASAP7_75t_L g525 ( .A(n_393), .B(n_526), .Y(n_525) );
AND2x4_ASAP7_75t_L g674 ( .A(n_393), .B(n_675), .Y(n_674) );
AND2x4_ASAP7_75t_L g738 ( .A(n_393), .B(n_526), .Y(n_738) );
AOI211xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B(n_397), .C(n_412), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_395), .A2(n_695), .B1(n_696), .B2(n_697), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_395), .A2(n_697), .B1(n_765), .B2(n_786), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_395), .A2(n_885), .B1(n_939), .B2(n_940), .Y(n_938) );
AOI22xp33_ASAP7_75t_SL g990 ( .A1(n_395), .A2(n_940), .B1(n_956), .B2(n_991), .Y(n_990) );
AOI22xp33_ASAP7_75t_SL g1306 ( .A1(n_395), .A2(n_940), .B1(n_1264), .B2(n_1307), .Y(n_1306) );
OAI22xp33_ASAP7_75t_L g515 ( .A1(n_396), .A2(n_509), .B1(n_516), .B2(n_518), .Y(n_515) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_403), .Y(n_398) );
AOI322xp5_ASAP7_75t_L g425 ( .A1(n_399), .A2(n_426), .A3(n_430), .B1(n_431), .B2(n_432), .C1(n_434), .C2(n_438), .Y(n_425) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g407 ( .A(n_400), .B(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g691 ( .A(n_400), .B(n_611), .Y(n_691) );
AND2x4_ASAP7_75t_L g693 ( .A(n_400), .B(n_408), .Y(n_693) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g422 ( .A(n_402), .Y(n_422) );
INVx2_ASAP7_75t_L g538 ( .A(n_403), .Y(n_538) );
BUFx2_ASAP7_75t_L g1201 ( .A(n_403), .Y(n_1201) );
BUFx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g545 ( .A(n_404), .Y(n_545) );
INVx1_ASAP7_75t_L g573 ( .A(n_404), .Y(n_573) );
INVx1_ASAP7_75t_L g602 ( .A(n_405), .Y(n_602) );
AND2x4_ASAP7_75t_L g611 ( .A(n_405), .B(n_612), .Y(n_611) );
INVx5_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_407), .A2(n_691), .B1(n_936), .B2(n_937), .Y(n_935) );
AOI22xp33_ASAP7_75t_SL g987 ( .A1(n_407), .A2(n_691), .B1(n_988), .B2(n_989), .Y(n_987) );
AOI22xp5_ASAP7_75t_L g1011 ( .A1(n_407), .A2(n_691), .B1(n_1012), .B2(n_1013), .Y(n_1011) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
HB1xp67_ASAP7_75t_L g1468 ( .A(n_409), .Y(n_1468) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g541 ( .A(n_410), .Y(n_541) );
INVx3_ASAP7_75t_L g549 ( .A(n_410), .Y(n_549) );
BUFx6f_ASAP7_75t_L g908 ( .A(n_410), .Y(n_908) );
AND2x4_ASAP7_75t_L g423 ( .A(n_411), .B(n_424), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g1085 ( .A1(n_413), .A2(n_1048), .B1(n_1049), .B2(n_1086), .C(n_1087), .Y(n_1085) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g1636 ( .A(n_414), .Y(n_1636) );
BUFx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g535 ( .A(n_415), .Y(n_535) );
INVx3_ASAP7_75t_L g580 ( .A(n_415), .Y(n_580) );
INVx2_ASAP7_75t_L g590 ( .A(n_415), .Y(n_590) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_416), .B(n_417), .Y(n_556) );
INVx1_ASAP7_75t_L g436 ( .A(n_417), .Y(n_436) );
NAND4xp25_ASAP7_75t_SL g688 ( .A(n_418), .B(n_689), .C(n_694), .D(n_699), .Y(n_688) );
NAND4xp25_ASAP7_75t_SL g774 ( .A(n_418), .B(n_775), .C(n_778), .D(n_785), .Y(n_774) );
CKINVDCx11_ASAP7_75t_R g418 ( .A(n_419), .Y(n_418) );
AOI211xp5_ASAP7_75t_L g930 ( .A1(n_419), .A2(n_834), .B(n_931), .C(n_932), .Y(n_930) );
AOI211xp5_ASAP7_75t_L g983 ( .A1(n_419), .A2(n_903), .B(n_984), .C(n_985), .Y(n_983) );
NOR3xp33_ASAP7_75t_L g1007 ( .A(n_419), .B(n_1008), .C(n_1010), .Y(n_1007) );
AOI211xp5_ASAP7_75t_L g1300 ( .A1(n_419), .A2(n_834), .B(n_1301), .C(n_1302), .Y(n_1300) );
AND2x4_ASAP7_75t_L g419 ( .A(n_420), .B(n_423), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g437 ( .A(n_421), .Y(n_437) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND2x1p5_ASAP7_75t_L g563 ( .A(n_422), .B(n_564), .Y(n_563) );
BUFx3_ASAP7_75t_L g623 ( .A(n_423), .Y(n_623) );
BUFx6f_ASAP7_75t_L g703 ( .A(n_423), .Y(n_703) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_423), .Y(n_723) );
BUFx2_ASAP7_75t_L g784 ( .A(n_423), .Y(n_784) );
BUFx3_ASAP7_75t_L g1174 ( .A(n_423), .Y(n_1174) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g792 ( .A(n_427), .Y(n_792) );
INVx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_428), .Y(n_596) );
AND2x4_ASAP7_75t_L g620 ( .A(n_428), .B(n_610), .Y(n_620) );
BUFx2_ASAP7_75t_L g833 ( .A(n_428), .Y(n_833) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx3_ASAP7_75t_L g583 ( .A(n_429), .Y(n_583) );
AOI322xp5_ASAP7_75t_L g473 ( .A1(n_431), .A2(n_438), .A3(n_474), .B1(n_476), .B2(n_477), .C1(n_478), .C2(n_482), .Y(n_473) );
INVx2_ASAP7_75t_L g706 ( .A(n_432), .Y(n_706) );
AOI222xp33_ASAP7_75t_L g778 ( .A1(n_432), .A2(n_434), .B1(n_779), .B2(n_780), .C1(n_781), .C2(n_782), .Y(n_778) );
INVx2_ASAP7_75t_L g933 ( .A(n_432), .Y(n_933) );
INVx2_ASAP7_75t_L g1009 ( .A(n_432), .Y(n_1009) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_433), .A2(n_599), .B1(n_600), .B2(n_601), .Y(n_598) );
INVx1_ASAP7_75t_L g842 ( .A(n_433), .Y(n_842) );
HB1xp67_ASAP7_75t_L g1081 ( .A(n_433), .Y(n_1081) );
AOI222xp33_ASAP7_75t_L g699 ( .A1(n_434), .A2(n_700), .B1(n_701), .B2(n_704), .C1(n_705), .C2(n_707), .Y(n_699) );
AND2x4_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI31xp33_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_450), .A3(n_467), .B(n_487), .Y(n_439) );
INVx4_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_442), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_442), .A2(n_761), .B1(n_762), .B2(n_763), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_442), .A2(n_460), .B1(n_885), .B2(n_886), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_442), .A2(n_752), .B1(n_958), .B2(n_959), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g1263 ( .A1(n_442), .A2(n_460), .B1(n_1264), .B2(n_1265), .Y(n_1263) );
AND2x6_ASAP7_75t_L g442 ( .A(n_443), .B(n_446), .Y(n_442) );
AND2x4_ASAP7_75t_L g749 ( .A(n_443), .B(n_750), .Y(n_749) );
AND2x4_ASAP7_75t_L g761 ( .A(n_443), .B(n_750), .Y(n_761) );
INVx1_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g744 ( .A(n_444), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g454 ( .A(n_445), .Y(n_454) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_445), .Y(n_462) );
AND2x2_ASAP7_75t_L g496 ( .A(n_445), .B(n_489), .Y(n_496) );
INVx2_ASAP7_75t_L g527 ( .A(n_445), .Y(n_527) );
INVx1_ASAP7_75t_L g523 ( .A(n_446), .Y(n_523) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_446), .Y(n_728) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_446), .Y(n_737) );
INVx2_ASAP7_75t_L g1064 ( .A(n_446), .Y(n_1064) );
INVx1_ASAP7_75t_L g1291 ( .A(n_446), .Y(n_1291) );
BUFx6f_ASAP7_75t_L g1589 ( .A(n_446), .Y(n_1589) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g506 ( .A(n_447), .Y(n_506) );
INVx1_ASAP7_75t_L g636 ( .A(n_447), .Y(n_636) );
INVx1_ASAP7_75t_L g679 ( .A(n_447), .Y(n_679) );
BUFx6f_ASAP7_75t_L g803 ( .A(n_447), .Y(n_803) );
AND2x4_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
INVx2_ASAP7_75t_L g466 ( .A(n_448), .Y(n_466) );
AND2x2_ASAP7_75t_L g472 ( .A(n_448), .B(n_465), .Y(n_472) );
INVx1_ASAP7_75t_L g456 ( .A(n_449), .Y(n_456) );
OR2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_455), .Y(n_451) );
INVx1_ASAP7_75t_L g476 ( .A(n_452), .Y(n_476) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g469 ( .A(n_453), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g486 ( .A(n_453), .Y(n_486) );
AND2x6_ASAP7_75t_L g752 ( .A(n_453), .B(n_475), .Y(n_752) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x6_ASAP7_75t_L g482 ( .A(n_454), .B(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g510 ( .A(n_455), .Y(n_510) );
INVx1_ASAP7_75t_L g1047 ( .A(n_455), .Y(n_1047) );
BUFx2_ASAP7_75t_L g1233 ( .A(n_455), .Y(n_1233) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_455), .B(n_670), .Y(n_1251) );
OR2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
AND2x2_ASAP7_75t_L g514 ( .A(n_456), .B(n_457), .Y(n_514) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g475 ( .A(n_458), .B(n_465), .Y(n_475) );
INVx4_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_460), .A2(n_696), .B1(n_748), .B2(n_749), .Y(n_747) );
AOI221xp5_ASAP7_75t_L g764 ( .A1(n_460), .A2(n_752), .B1(n_765), .B2(n_766), .C(n_767), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_460), .A2(n_761), .B1(n_955), .B2(n_956), .Y(n_954) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_463), .Y(n_460) );
AND2x2_ASAP7_75t_SL g478 ( .A(n_461), .B(n_479), .Y(n_478) );
AND2x4_ASAP7_75t_L g892 ( .A(n_461), .B(n_479), .Y(n_892) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx6_ASAP7_75t_L g632 ( .A(n_463), .Y(n_632) );
INVx2_ASAP7_75t_L g667 ( .A(n_463), .Y(n_667) );
AND2x2_ASAP7_75t_L g675 ( .A(n_463), .B(n_653), .Y(n_675) );
BUFx2_ASAP7_75t_L g733 ( .A(n_463), .Y(n_733) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g483 ( .A(n_464), .Y(n_483) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g481 ( .A(n_466), .Y(n_481) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AOI211xp5_ASAP7_75t_L g740 ( .A1(n_469), .A2(n_485), .B(n_741), .C(n_742), .Y(n_740) );
HB1xp67_ASAP7_75t_L g889 ( .A(n_470), .Y(n_889) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_470), .Y(n_951) );
HB1xp67_ASAP7_75t_L g1294 ( .A(n_470), .Y(n_1294) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x4_ASAP7_75t_L g485 ( .A(n_471), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g629 ( .A(n_471), .Y(n_629) );
BUFx6f_ASAP7_75t_L g771 ( .A(n_471), .Y(n_771) );
INVx1_ASAP7_75t_L g877 ( .A(n_471), .Y(n_877) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_472), .Y(n_662) );
INVx2_ASAP7_75t_L g502 ( .A(n_474), .Y(n_502) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_SL g521 ( .A(n_475), .Y(n_521) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_475), .Y(n_635) );
BUFx2_ASAP7_75t_L g727 ( .A(n_475), .Y(n_727) );
BUFx6f_ASAP7_75t_L g928 ( .A(n_475), .Y(n_928) );
BUFx6f_ASAP7_75t_L g1062 ( .A(n_475), .Y(n_1062) );
BUFx3_ASAP7_75t_L g1289 ( .A(n_475), .Y(n_1289) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_477), .A2(n_543), .B1(n_546), .B2(n_550), .Y(n_542) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g745 ( .A(n_480), .Y(n_745) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g650 ( .A(n_481), .Y(n_650) );
INVx3_ASAP7_75t_L g746 ( .A(n_482), .Y(n_746) );
AOI222xp33_ASAP7_75t_L g887 ( .A1(n_482), .A2(n_888), .B1(n_889), .B2(n_890), .C1(n_891), .C2(n_893), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_482), .A2(n_892), .B1(n_1001), .B2(n_1002), .Y(n_1000) );
AOI222xp33_ASAP7_75t_L g1266 ( .A1(n_482), .A2(n_892), .B1(n_1024), .B2(n_1267), .C1(n_1268), .C2(n_1269), .Y(n_1266) );
BUFx3_ASAP7_75t_L g659 ( .A(n_483), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g995 ( .A(n_484), .B(n_996), .C(n_1000), .Y(n_995) );
CKINVDCx8_ASAP7_75t_R g484 ( .A(n_485), .Y(n_484) );
INVx5_ASAP7_75t_L g883 ( .A(n_485), .Y(n_883) );
AOI211xp5_ASAP7_75t_L g949 ( .A1(n_485), .A2(n_950), .B(n_951), .C(n_952), .Y(n_949) );
OAI21xp33_ASAP7_75t_L g769 ( .A1(n_486), .A2(n_770), .B(n_771), .Y(n_769) );
INVx1_ASAP7_75t_SL g755 ( .A(n_487), .Y(n_755) );
OAI31xp33_ASAP7_75t_L g994 ( .A1(n_487), .A2(n_995), .A3(n_1003), .B(n_1005), .Y(n_994) );
AND2x4_ASAP7_75t_L g487 ( .A(n_488), .B(n_490), .Y(n_487) );
AND2x4_ASAP7_75t_L g773 ( .A(n_488), .B(n_490), .Y(n_773) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x4_ASAP7_75t_L g526 ( .A(n_489), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g1159 ( .A(n_490), .Y(n_1159) );
BUFx2_ASAP7_75t_L g1255 ( .A(n_490), .Y(n_1255) );
BUFx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g497 ( .A(n_491), .Y(n_497) );
OR2x6_ASAP7_75t_L g529 ( .A(n_491), .B(n_530), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_528), .Y(n_492) );
OAI33xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_498), .A3(n_507), .B1(n_515), .B2(n_519), .B3(n_524), .Y(n_493) );
INVx1_ASAP7_75t_SL g725 ( .A(n_494), .Y(n_725) );
OAI33xp33_ASAP7_75t_L g1442 ( .A1(n_494), .A2(n_524), .A3(n_1443), .B1(n_1446), .B2(n_1449), .B3(n_1452), .Y(n_1442) );
OAI22xp5_ASAP7_75t_L g1583 ( .A1(n_494), .A2(n_1051), .B1(n_1584), .B2(n_1590), .Y(n_1583) );
OR2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_497), .Y(n_494) );
OR2x6_ASAP7_75t_L g638 ( .A(n_495), .B(n_497), .Y(n_638) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g807 ( .A(n_496), .Y(n_807) );
INVx2_ASAP7_75t_SL g1243 ( .A(n_496), .Y(n_1243) );
INVx2_ASAP7_75t_L g625 ( .A(n_497), .Y(n_625) );
AND2x4_ASAP7_75t_L g710 ( .A(n_497), .B(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g806 ( .A(n_497), .B(n_807), .Y(n_806) );
AND2x4_ASAP7_75t_L g900 ( .A(n_497), .B(n_711), .Y(n_900) );
BUFx2_ASAP7_75t_L g1101 ( .A(n_497), .Y(n_1101) );
OAI31xp33_ASAP7_75t_L g1904 ( .A1(n_497), .A2(n_1905), .A3(n_1906), .B(n_1918), .Y(n_1904) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B1(n_503), .B2(n_504), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_499), .A2(n_503), .B1(n_537), .B2(n_539), .Y(n_536) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_502), .A2(n_643), .B1(n_644), .B2(n_646), .Y(n_642) );
INVx2_ASAP7_75t_SL g1531 ( .A(n_502), .Y(n_1531) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g645 ( .A(n_506), .Y(n_645) );
OR2x2_ASAP7_75t_L g1253 ( .A(n_506), .B(n_670), .Y(n_1253) );
OAI22xp33_ASAP7_75t_SL g507 ( .A1(n_508), .A2(n_509), .B1(n_511), .B2(n_512), .Y(n_507) );
OAI22xp33_ASAP7_75t_L g531 ( .A1(n_508), .A2(n_511), .B1(n_532), .B2(n_533), .Y(n_531) );
OAI22xp33_ASAP7_75t_L g1449 ( .A1(n_509), .A2(n_516), .B1(n_1450), .B2(n_1451), .Y(n_1449) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g1054 ( .A(n_510), .Y(n_1054) );
INVx1_ASAP7_75t_L g1107 ( .A(n_510), .Y(n_1107) );
OAI221xp5_ASAP7_75t_L g1590 ( .A1(n_512), .A2(n_1233), .B1(n_1591), .B2(n_1592), .C(n_1593), .Y(n_1590) );
BUFx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g1332 ( .A(n_513), .Y(n_1332) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g517 ( .A(n_514), .Y(n_517) );
BUFx4f_ASAP7_75t_L g1058 ( .A(n_514), .Y(n_1058) );
OAI22xp33_ASAP7_75t_L g1446 ( .A1(n_516), .A2(n_1233), .B1(n_1447), .B2(n_1448), .Y(n_1446) );
BUFx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
OR2x6_ASAP7_75t_L g681 ( .A(n_517), .B(n_669), .Y(n_681) );
OAI221xp5_ASAP7_75t_L g1044 ( .A1(n_517), .A2(n_1045), .B1(n_1048), .B2(n_1049), .C(n_1050), .Y(n_1044) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B1(n_522), .B2(n_523), .Y(n_519) );
INVx2_ASAP7_75t_L g673 ( .A(n_521), .Y(n_673) );
INVx1_ASAP7_75t_L g980 ( .A(n_521), .Y(n_980) );
OAI22xp5_ASAP7_75t_SL g1322 ( .A1(n_524), .A2(n_638), .B1(n_1323), .B2(n_1329), .Y(n_1322) );
INVx4_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_525), .A2(n_627), .B1(n_637), .B2(n_639), .C(n_647), .Y(n_626) );
AOI33xp33_ASAP7_75t_L g915 ( .A1(n_525), .A2(n_916), .A3(n_917), .B1(n_922), .B2(n_924), .B3(n_926), .Y(n_915) );
AOI33xp33_ASAP7_75t_L g1019 ( .A1(n_525), .A2(n_916), .A3(n_1020), .B1(n_1023), .B2(n_1025), .B3(n_1028), .Y(n_1019) );
BUFx4f_ASAP7_75t_L g1052 ( .A(n_525), .Y(n_1052) );
BUFx4f_ASAP7_75t_L g1123 ( .A(n_525), .Y(n_1123) );
AOI33xp33_ASAP7_75t_L g1286 ( .A1(n_525), .A2(n_916), .A3(n_1287), .B1(n_1292), .B2(n_1295), .B3(n_1298), .Y(n_1286) );
INVx2_ASAP7_75t_L g1235 ( .A(n_526), .Y(n_1235) );
AND2x4_ASAP7_75t_L g653 ( .A(n_527), .B(n_654), .Y(n_653) );
OAI33xp33_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_531), .A3(n_536), .B1(n_542), .B2(n_551), .B3(n_558), .Y(n_528) );
OAI33xp33_ASAP7_75t_L g1190 ( .A1(n_529), .A2(n_558), .A3(n_1191), .B1(n_1199), .B2(n_1204), .B3(n_1208), .Y(n_1190) );
INVx1_ASAP7_75t_L g1419 ( .A(n_529), .Y(n_1419) );
OAI22xp33_ASAP7_75t_L g551 ( .A1(n_532), .A2(n_552), .B1(n_553), .B2(n_557), .Y(n_551) );
BUFx2_ASAP7_75t_L g1086 ( .A(n_532), .Y(n_1086) );
OAI221xp5_ASAP7_75t_L g1509 ( .A1(n_532), .A2(n_555), .B1(n_1087), .B2(n_1510), .C(n_1511), .Y(n_1509) );
OAI221xp5_ASAP7_75t_L g1513 ( .A1(n_532), .A2(n_580), .B1(n_1474), .B2(n_1499), .C(n_1514), .Y(n_1513) );
INVx1_ASAP7_75t_L g1638 ( .A(n_532), .Y(n_1638) );
INVx1_ASAP7_75t_L g1927 ( .A(n_532), .Y(n_1927) );
OAI221xp5_ASAP7_75t_L g1924 ( .A1(n_533), .A2(n_1352), .B1(n_1925), .B2(n_1926), .C(n_1928), .Y(n_1924) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_535), .B(n_598), .Y(n_597) );
OR2x6_ASAP7_75t_L g854 ( .A(n_535), .B(n_604), .Y(n_854) );
OR2x2_ASAP7_75t_L g1097 ( .A(n_535), .B(n_604), .Y(n_1097) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g973 ( .A(n_539), .Y(n_973) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x4_ASAP7_75t_L g615 ( .A(n_540), .B(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g852 ( .A(n_541), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g1505 ( .A1(n_543), .A2(n_1506), .B1(n_1507), .B2(n_1508), .Y(n_1505) );
INVx2_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g1154 ( .A(n_544), .Y(n_1154) );
INVx2_ASAP7_75t_L g1428 ( .A(n_544), .Y(n_1428) );
INVx2_ASAP7_75t_L g1465 ( .A(n_544), .Y(n_1465) );
BUFx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g1072 ( .A(n_545), .Y(n_1072) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g797 ( .A(n_548), .Y(n_797) );
INVx2_ASAP7_75t_L g1280 ( .A(n_548), .Y(n_1280) );
INVx3_ASAP7_75t_L g1519 ( .A(n_548), .Y(n_1519) );
INVx2_ASAP7_75t_L g1922 ( .A(n_548), .Y(n_1922) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx3_ASAP7_75t_L g576 ( .A(n_549), .Y(n_576) );
INVx3_ASAP7_75t_L g1095 ( .A(n_549), .Y(n_1095) );
OAI221xp5_ASAP7_75t_L g1471 ( .A1(n_553), .A2(n_1421), .B1(n_1472), .B2(n_1473), .C(n_1474), .Y(n_1471) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g1423 ( .A(n_554), .Y(n_1423) );
INVx2_ASAP7_75t_L g1908 ( .A(n_554), .Y(n_1908) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx3_ASAP7_75t_L g1433 ( .A(n_555), .Y(n_1433) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AOI33xp33_ASAP7_75t_L g709 ( .A1(n_559), .A2(n_710), .A3(n_712), .B1(n_715), .B2(n_719), .B3(n_721), .Y(n_709) );
AOI33xp33_ASAP7_75t_L g898 ( .A1(n_559), .A2(n_899), .A3(n_901), .B1(n_904), .B2(n_909), .B3(n_914), .Y(n_898) );
AOI33xp33_ASAP7_75t_L g1014 ( .A1(n_559), .A2(n_710), .A3(n_1015), .B1(n_1016), .B2(n_1017), .B3(n_1018), .Y(n_1014) );
INVx6_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx5_ASAP7_75t_L g799 ( .A(n_560), .Y(n_799) );
OR2x6_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
NAND2x1p5_ASAP7_75t_L g652 ( .A(n_561), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g669 ( .A(n_562), .B(n_670), .Y(n_669) );
AND2x4_ASAP7_75t_L g1171 ( .A(n_562), .B(n_610), .Y(n_1171) );
BUFx2_ASAP7_75t_L g593 ( .A(n_563), .Y(n_593) );
INVx2_ASAP7_75t_L g837 ( .A(n_563), .Y(n_837) );
NAND4xp25_ASAP7_75t_L g568 ( .A(n_569), .B(n_626), .C(n_664), .D(n_676), .Y(n_568) );
OAI31xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_607), .A3(n_618), .B(n_624), .Y(n_569) );
OAI221xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_578), .B1(n_584), .B2(n_588), .C(n_594), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_574), .B1(n_575), .B2(n_577), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_572), .A2(n_585), .B1(n_586), .B2(n_587), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g1639 ( .A1(n_572), .A2(n_907), .B1(n_1640), .B2(n_1641), .Y(n_1639) );
BUFx2_ASAP7_75t_L g1912 ( .A(n_572), .Y(n_1912) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g1091 ( .A(n_573), .Y(n_1091) );
INVx1_ASAP7_75t_L g1517 ( .A(n_573), .Y(n_1517) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_574), .A2(n_577), .B1(n_634), .B2(n_636), .Y(n_633) );
INVx2_ASAP7_75t_L g720 ( .A(n_575), .Y(n_720) );
INVx2_ASAP7_75t_SL g790 ( .A(n_575), .Y(n_790) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g586 ( .A(n_576), .Y(n_586) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_576), .Y(n_831) );
INVx1_ASAP7_75t_L g1349 ( .A(n_576), .Y(n_1349) );
OAI21xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_580), .B(n_581), .Y(n_578) );
BUFx2_ASAP7_75t_L g1147 ( .A(n_580), .Y(n_1147) );
INVx1_ASAP7_75t_L g1197 ( .A(n_580), .Y(n_1197) );
OAI221xp5_ASAP7_75t_L g1469 ( .A1(n_580), .A2(n_1193), .B1(n_1352), .B2(n_1447), .C(n_1448), .Y(n_1469) );
BUFx2_ASAP7_75t_L g713 ( .A(n_582), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_582), .B(n_826), .Y(n_825) );
INVx2_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g592 ( .A(n_583), .Y(n_592) );
INVx2_ASAP7_75t_SL g1143 ( .A(n_583), .Y(n_1143) );
AOI222xp33_ASAP7_75t_L g664 ( .A1(n_585), .A2(n_595), .B1(n_665), .B2(n_671), .C1(n_672), .C2(n_674), .Y(n_664) );
INVx1_ASAP7_75t_L g718 ( .A(n_586), .Y(n_718) );
INVx2_ASAP7_75t_L g968 ( .A(n_586), .Y(n_968) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_587), .A2(n_589), .B1(n_677), .B2(n_680), .Y(n_676) );
OAI21xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B(n_591), .Y(n_588) );
OAI221xp5_ASAP7_75t_L g1351 ( .A1(n_590), .A2(n_1086), .B1(n_1324), .B2(n_1325), .C(n_1352), .Y(n_1351) );
BUFx3_ASAP7_75t_L g902 ( .A(n_592), .Y(n_902) );
A2O1A1Ixp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B(n_597), .C(n_603), .Y(n_594) );
NAND2x1p5_ASAP7_75t_L g1187 ( .A(n_601), .B(n_1184), .Y(n_1187) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OR2x6_ASAP7_75t_L g844 ( .A(n_602), .B(n_604), .Y(n_844) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g826 ( .A(n_604), .Y(n_826) );
INVx1_ASAP7_75t_L g843 ( .A(n_604), .Y(n_843) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx3_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_609), .A2(n_615), .B1(n_846), .B2(n_847), .Y(n_845) );
INVx3_ASAP7_75t_L g1099 ( .A(n_609), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1542 ( .A1(n_609), .A2(n_615), .B1(n_1543), .B2(n_1544), .Y(n_1542) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx2_ASAP7_75t_L g617 ( .A(n_610), .Y(n_617) );
INVx1_ASAP7_75t_L g717 ( .A(n_611), .Y(n_717) );
BUFx6f_ASAP7_75t_L g830 ( .A(n_611), .Y(n_830) );
BUFx2_ASAP7_75t_L g905 ( .A(n_611), .Y(n_905) );
BUFx6f_ASAP7_75t_L g912 ( .A(n_611), .Y(n_912) );
BUFx2_ASAP7_75t_L g972 ( .A(n_611), .Y(n_972) );
BUFx6f_ASAP7_75t_L g1278 ( .A(n_611), .Y(n_1278) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx3_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx3_ASAP7_75t_L g1100 ( .A(n_615), .Y(n_1100) );
AND2x4_ASAP7_75t_L g622 ( .A(n_616), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
CKINVDCx6p67_ASAP7_75t_R g619 ( .A(n_620), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g848 ( .A1(n_620), .A2(n_849), .B1(n_850), .B2(n_851), .C(n_853), .Y(n_848) );
AOI221xp5_ASAP7_75t_L g1545 ( .A1(n_620), .A2(n_853), .B1(n_1546), .B2(n_1548), .C(n_1549), .Y(n_1545) );
INVx8_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AOI221xp5_ASAP7_75t_SL g828 ( .A1(n_622), .A2(n_829), .B1(n_832), .B2(n_838), .C(n_839), .Y(n_828) );
AOI221xp5_ASAP7_75t_L g1537 ( .A1(n_622), .A2(n_1538), .B1(n_1539), .B2(n_1540), .C(n_1541), .Y(n_1537) );
INVx1_ASAP7_75t_L g835 ( .A(n_623), .Y(n_835) );
INVx1_ASAP7_75t_L g855 ( .A(n_624), .Y(n_855) );
OAI31xp33_ASAP7_75t_L g1632 ( .A1(n_624), .A2(n_1633), .A3(n_1634), .B(n_1642), .Y(n_1632) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NOR2xp67_ASAP7_75t_L g824 ( .A(n_625), .B(n_825), .Y(n_824) );
INVx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g861 ( .A(n_629), .Y(n_861) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_632), .Y(n_641) );
INVx2_ASAP7_75t_L g731 ( .A(n_632), .Y(n_731) );
INVx2_ASAP7_75t_L g750 ( .A(n_632), .Y(n_750) );
INVx1_ASAP7_75t_L g810 ( .A(n_632), .Y(n_810) );
INVx2_ASAP7_75t_L g919 ( .A(n_632), .Y(n_919) );
INVx1_ASAP7_75t_L g1571 ( .A(n_632), .Y(n_1571) );
INVx1_ASAP7_75t_L g1021 ( .A(n_634), .Y(n_1021) );
INVx1_ASAP7_75t_L g1381 ( .A(n_634), .Y(n_1381) );
INVx1_ASAP7_75t_L g1528 ( .A(n_634), .Y(n_1528) );
INVx2_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
BUFx3_ASAP7_75t_L g923 ( .A(n_635), .Y(n_923) );
AND2x4_ASAP7_75t_L g1220 ( .A(n_635), .B(n_1221), .Y(n_1220) );
INVx1_ASAP7_75t_L g1022 ( .A(n_636), .Y(n_1022) );
INVx1_ASAP7_75t_L g1029 ( .A(n_636), .Y(n_1029) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g916 ( .A(n_638), .Y(n_916) );
OAI22xp5_ASAP7_75t_SL g1043 ( .A1(n_638), .A2(n_1044), .B1(n_1051), .B2(n_1053), .Y(n_1043) );
CKINVDCx5p33_ASAP7_75t_R g1524 ( .A(n_638), .Y(n_1524) );
OAI22xp5_ASAP7_75t_SL g1622 ( .A1(n_638), .A2(n_1051), .B1(n_1623), .B2(n_1627), .Y(n_1622) );
INVx4_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g978 ( .A(n_641), .Y(n_978) );
INVx1_ASAP7_75t_L g1378 ( .A(n_641), .Y(n_1378) );
INVx1_ASAP7_75t_L g965 ( .A(n_644), .Y(n_965) );
INVx1_ASAP7_75t_L g981 ( .A(n_644), .Y(n_981) );
INVx2_ASAP7_75t_SL g1937 ( .A(n_644), .Y(n_1937) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx2_ASAP7_75t_L g1383 ( .A(n_645), .Y(n_1383) );
INVx2_ASAP7_75t_L g873 ( .A(n_648), .Y(n_873) );
INVx1_ASAP7_75t_L g1042 ( .A(n_648), .Y(n_1042) );
HB1xp67_ASAP7_75t_L g1338 ( .A(n_648), .Y(n_1338) );
INVx2_ASAP7_75t_L g1563 ( .A(n_648), .Y(n_1563) );
INVx1_ASAP7_75t_L g1934 ( .A(n_648), .Y(n_1934) );
NAND2x1p5_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g1225 ( .A(n_650), .Y(n_1225) );
INVx2_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
OR2x6_ASAP7_75t_L g657 ( .A(n_652), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g663 ( .A(n_652), .Y(n_663) );
OR2x2_ASAP7_75t_L g1458 ( .A(n_652), .B(n_658), .Y(n_1458) );
AND2x4_ASAP7_75t_L g1224 ( .A(n_653), .B(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1227 ( .A(n_653), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_653), .B(n_659), .Y(n_1388) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g871 ( .A(n_657), .Y(n_871) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_658), .B(n_1227), .Y(n_1226) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND3xp33_ASAP7_75t_SL g1113 ( .A(n_660), .B(n_1114), .C(n_1117), .Y(n_1113) );
INVx1_ASAP7_75t_L g1561 ( .A(n_660), .Y(n_1561) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
INVx1_ASAP7_75t_L g1297 ( .A(n_661), .Y(n_1297) );
HB1xp67_ASAP7_75t_L g1573 ( .A(n_661), .Y(n_1573) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g735 ( .A(n_662), .Y(n_735) );
INVx2_ASAP7_75t_SL g999 ( .A(n_662), .Y(n_999) );
BUFx3_ASAP7_75t_L g1024 ( .A(n_662), .Y(n_1024) );
AND2x4_ASAP7_75t_L g1239 ( .A(n_662), .B(n_1221), .Y(n_1239) );
INVx1_ASAP7_75t_L g1242 ( .A(n_662), .Y(n_1242) );
BUFx4f_ASAP7_75t_L g1526 ( .A(n_662), .Y(n_1526) );
AND2x2_ASAP7_75t_L g875 ( .A(n_663), .B(n_876), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_665), .A2(n_672), .B1(n_868), .B2(n_869), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g1128 ( .A1(n_665), .A2(n_672), .B1(n_1129), .B2(n_1130), .Y(n_1128) );
AOI221xp5_ASAP7_75t_L g1497 ( .A1(n_665), .A2(n_672), .B1(n_1498), .B2(n_1499), .C(n_1500), .Y(n_1497) );
AOI22xp33_ASAP7_75t_L g1551 ( .A1(n_665), .A2(n_672), .B1(n_1552), .B2(n_1553), .Y(n_1551) );
AOI22xp33_ASAP7_75t_L g1946 ( .A1(n_665), .A2(n_672), .B1(n_1910), .B2(n_1913), .Y(n_1946) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
BUFx2_ASAP7_75t_L g1293 ( .A(n_666), .Y(n_1293) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g925 ( .A(n_667), .Y(n_925) );
AND2x2_ASAP7_75t_L g672 ( .A(n_668), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OR2x6_ASAP7_75t_L g678 ( .A(n_669), .B(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_669), .B(n_679), .Y(n_1104) );
OR2x2_ASAP7_75t_L g1106 ( .A(n_669), .B(n_1107), .Y(n_1106) );
OR2x2_ASAP7_75t_L g1108 ( .A(n_669), .B(n_1109), .Y(n_1108) );
INVx2_ASAP7_75t_L g1221 ( .A(n_670), .Y(n_1221) );
OR2x6_ASAP7_75t_L g823 ( .A(n_674), .B(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g1216 ( .A(n_674), .Y(n_1216) );
AOI22xp5_ASAP7_75t_L g864 ( .A1(n_677), .A2(n_680), .B1(n_865), .B2(n_866), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_677), .A2(n_680), .B1(n_1126), .B2(n_1127), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g1554 ( .A1(n_677), .A2(n_680), .B1(n_1555), .B2(n_1556), .Y(n_1554) );
AOI22xp33_ASAP7_75t_L g1945 ( .A1(n_677), .A2(n_680), .B1(n_1909), .B2(n_1914), .Y(n_1945) );
CKINVDCx6p67_ASAP7_75t_R g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g859 ( .A(n_679), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g1452 ( .A1(n_679), .A2(n_1453), .B1(n_1454), .B2(n_1455), .Y(n_1452) );
CKINVDCx6p67_ASAP7_75t_R g680 ( .A(n_681), .Y(n_680) );
OA22x2_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_756), .B1(n_757), .B2(n_814), .Y(n_682) );
INVx1_ASAP7_75t_L g814 ( .A(n_683), .Y(n_814) );
XNOR2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g1692 ( .A1(n_684), .A2(n_1693), .B1(n_1695), .B2(n_1696), .Y(n_1692) );
AOI211xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B(n_708), .C(n_739), .Y(n_685) );
AOI221x1_ASAP7_75t_L g758 ( .A1(n_686), .A2(n_759), .B1(n_772), .B2(n_774), .C(n_787), .Y(n_758) );
CKINVDCx16_ASAP7_75t_R g686 ( .A(n_687), .Y(n_686) );
AOI31xp33_ASAP7_75t_L g982 ( .A1(n_687), .A2(n_983), .A3(n_987), .B(n_990), .Y(n_982) );
AO21x1_ASAP7_75t_SL g1006 ( .A1(n_687), .A2(n_1007), .B(n_1011), .Y(n_1006) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B1(n_692), .B2(n_693), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_691), .A2(n_693), .B1(n_776), .B2(n_777), .Y(n_775) );
AOI22xp33_ASAP7_75t_SL g1303 ( .A1(n_691), .A2(n_693), .B1(n_1304), .B2(n_1305), .Y(n_1303) );
INVx4_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx5_ASAP7_75t_L g940 ( .A(n_698), .Y(n_940) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_SL g903 ( .A(n_702), .Y(n_903) );
INVx2_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_703), .Y(n_714) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_709), .B(n_724), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g788 ( .A(n_710), .B(n_789), .C(n_791), .Y(n_788) );
BUFx2_ASAP7_75t_SL g1087 ( .A(n_711), .Y(n_1087) );
INVx1_ASAP7_75t_L g1353 ( .A(n_711), .Y(n_1353) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
BUFx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_SL g794 ( .A(n_723), .Y(n_794) );
HB1xp67_ASAP7_75t_L g975 ( .A(n_723), .Y(n_975) );
AOI33xp33_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .A3(n_729), .B1(n_732), .B2(n_736), .B3(n_738), .Y(n_724) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g1246 ( .A(n_731), .Y(n_1246) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g808 ( .A(n_738), .B(n_809), .C(n_811), .Y(n_808) );
AOI33xp33_ASAP7_75t_L g857 ( .A1(n_738), .A2(n_805), .A3(n_858), .B1(n_860), .B2(n_862), .B3(n_863), .Y(n_857) );
NAND3xp33_ASAP7_75t_L g976 ( .A(n_738), .B(n_977), .C(n_979), .Y(n_976) );
INVx1_ASAP7_75t_L g1943 ( .A(n_738), .Y(n_1943) );
AOI31xp33_ASAP7_75t_SL g739 ( .A1(n_740), .A2(n_747), .A3(n_751), .B(n_755), .Y(n_739) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g768 ( .A(n_744), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g1260 ( .A1(n_749), .A2(n_752), .B1(n_1261), .B2(n_1262), .Y(n_1260) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_752), .A2(n_761), .B1(n_895), .B2(n_896), .Y(n_894) );
CKINVDCx6p67_ASAP7_75t_R g1004 ( .A(n_752), .Y(n_1004) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g813 ( .A(n_758), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_764), .Y(n_759) );
INVx1_ASAP7_75t_L g921 ( .A(n_771), .Y(n_921) );
BUFx6f_ASAP7_75t_L g1027 ( .A(n_771), .Y(n_1027) );
AND2x4_ASAP7_75t_L g1247 ( .A(n_771), .B(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1393 ( .A(n_771), .Y(n_1393) );
BUFx6f_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
AOI211x1_ASAP7_75t_SL g881 ( .A1(n_773), .A2(n_882), .B(n_897), .C(n_929), .Y(n_881) );
AO211x2_ASAP7_75t_L g947 ( .A1(n_773), .A2(n_948), .B(n_960), .C(n_982), .Y(n_947) );
INVx1_ASAP7_75t_L g1271 ( .A(n_773), .Y(n_1271) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NAND4xp25_ASAP7_75t_L g787 ( .A(n_788), .B(n_795), .C(n_800), .D(n_808), .Y(n_787) );
INVx1_ASAP7_75t_L g1478 ( .A(n_790), .Y(n_1478) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NAND3xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_798), .C(n_799), .Y(n_795) );
INVx1_ASAP7_75t_L g1600 ( .A(n_797), .Y(n_1600) );
NAND3xp33_ASAP7_75t_L g966 ( .A(n_799), .B(n_967), .C(n_969), .Y(n_966) );
AOI33xp33_ASAP7_75t_L g1273 ( .A1(n_799), .A2(n_1274), .A3(n_1276), .B1(n_1281), .B2(n_1283), .B3(n_1285), .Y(n_1273) );
CKINVDCx8_ASAP7_75t_R g1434 ( .A(n_799), .Y(n_1434) );
NAND3xp33_ASAP7_75t_L g800 ( .A(n_801), .B(n_804), .C(n_805), .Y(n_800) );
BUFx6f_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g1230 ( .A(n_803), .Y(n_1230) );
INVx1_ASAP7_75t_L g1328 ( .A(n_803), .Y(n_1328) );
BUFx3_ASAP7_75t_L g1397 ( .A(n_803), .Y(n_1397) );
NAND3xp33_ASAP7_75t_L g961 ( .A(n_805), .B(n_962), .C(n_963), .Y(n_961) );
INVx3_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_817), .B1(n_944), .B2(n_1032), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
AOI21x1_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_879), .B(n_943), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
AND2x2_ASAP7_75t_L g943 ( .A(n_819), .B(n_880), .Y(n_943) );
XOR2x2_ASAP7_75t_L g819 ( .A(n_820), .B(n_878), .Y(n_819) );
NOR3xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_827), .C(n_856), .Y(n_820) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_823), .B(n_1066), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_823), .B(n_1132), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_823), .B(n_1340), .Y(n_1339) );
NAND2xp5_ASAP7_75t_L g1459 ( .A(n_823), .B(n_1460), .Y(n_1459) );
NAND2xp5_ASAP7_75t_L g1501 ( .A(n_823), .B(n_1502), .Y(n_1501) );
INVx1_ASAP7_75t_L g1558 ( .A(n_823), .Y(n_1558) );
NAND2xp5_ASAP7_75t_L g1580 ( .A(n_823), .B(n_1581), .Y(n_1580) );
NAND2xp5_ASAP7_75t_L g1619 ( .A(n_823), .B(n_1620), .Y(n_1619) );
NAND2xp5_ASAP7_75t_L g1929 ( .A(n_823), .B(n_1930), .Y(n_1929) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_826), .B(n_1081), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_826), .B(n_1081), .Y(n_1362) );
AOI31xp33_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_845), .A3(n_848), .B(n_855), .Y(n_827) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g1474 ( .A(n_836), .Y(n_1474) );
INVx2_ASAP7_75t_SL g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g1077 ( .A(n_837), .Y(n_1077) );
NAND2x1p5_ASAP7_75t_L g840 ( .A(n_841), .B(n_843), .Y(n_840) );
NAND2x1_ASAP7_75t_SL g1183 ( .A(n_841), .B(n_1184), .Y(n_1183) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
CKINVDCx11_ASAP7_75t_R g1083 ( .A(n_844), .Y(n_1083) );
INVx1_ASAP7_75t_L g1139 ( .A(n_852), .Y(n_1139) );
INVx2_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
NAND4xp25_ASAP7_75t_L g856 ( .A(n_857), .B(n_864), .C(n_867), .D(n_870), .Y(n_856) );
AOI221xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B1(n_873), .B2(n_874), .C(n_875), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_871), .A2(n_1042), .B1(n_1115), .B2(n_1116), .Y(n_1114) );
AOI221xp5_ASAP7_75t_L g1494 ( .A1(n_871), .A2(n_875), .B1(n_1042), .B2(n_1495), .C(n_1496), .Y(n_1494) );
AOI22xp5_ASAP7_75t_L g1562 ( .A1(n_871), .A2(n_1563), .B1(n_1564), .B2(n_1565), .Y(n_1562) );
AOI22xp5_ASAP7_75t_L g1933 ( .A1(n_871), .A2(n_1916), .B1(n_1917), .B2(n_1934), .Y(n_1933) );
INVx2_ASAP7_75t_L g1457 ( .A(n_873), .Y(n_1457) );
BUFx2_ASAP7_75t_L g1039 ( .A(n_875), .Y(n_1039) );
HB1xp67_ASAP7_75t_L g1441 ( .A(n_875), .Y(n_1441) );
NOR3xp33_ASAP7_75t_SL g1582 ( .A(n_875), .B(n_1583), .C(n_1594), .Y(n_1582) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g1377 ( .A(n_877), .Y(n_1377) );
INVx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g942 ( .A(n_881), .Y(n_942) );
NAND4xp25_ASAP7_75t_L g882 ( .A(n_883), .B(n_884), .C(n_887), .D(n_894), .Y(n_882) );
NAND4xp25_ASAP7_75t_L g1259 ( .A(n_883), .B(n_1260), .C(n_1263), .D(n_1266), .Y(n_1259) );
BUFx4f_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g953 ( .A(n_892), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_898), .B(n_915), .Y(n_897) );
BUFx3_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
NAND3xp33_ASAP7_75t_L g970 ( .A(n_900), .B(n_971), .C(n_974), .Y(n_970) );
INVx2_ASAP7_75t_L g1275 ( .A(n_900), .Y(n_1275) );
INVx2_ASAP7_75t_SL g906 ( .A(n_907), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g1431 ( .A1(n_907), .A2(n_1384), .B1(n_1402), .B2(n_1426), .Y(n_1431) );
OAI221xp5_ASAP7_75t_L g1605 ( .A1(n_907), .A2(n_1428), .B1(n_1606), .B2(n_1607), .C(n_1608), .Y(n_1605) );
INVx4_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
BUFx3_ASAP7_75t_L g913 ( .A(n_908), .Y(n_913) );
INVx2_ASAP7_75t_SL g1203 ( .A(n_908), .Y(n_1203) );
INVx2_ASAP7_75t_SL g1206 ( .A(n_908), .Y(n_1206) );
INVx2_ASAP7_75t_SL g1507 ( .A(n_908), .Y(n_1507) );
INVx3_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx2_ASAP7_75t_SL g911 ( .A(n_912), .Y(n_911) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_912), .B(n_1171), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_912), .B(n_1171), .Y(n_1414) );
INVx1_ASAP7_75t_L g1156 ( .A(n_913), .Y(n_1156) );
AOI33xp33_ASAP7_75t_L g1117 ( .A1(n_916), .A2(n_1118), .A3(n_1120), .B1(n_1121), .B2(n_1122), .B3(n_1123), .Y(n_1117) );
AOI33xp33_ASAP7_75t_L g1566 ( .A1(n_916), .A2(n_1123), .A3(n_1567), .B1(n_1568), .B2(n_1572), .B3(n_1574), .Y(n_1566) );
BUFx3_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
HB1xp67_ASAP7_75t_L g1026 ( .A(n_919), .Y(n_1026) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
BUFx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
BUFx4f_ASAP7_75t_L g964 ( .A(n_928), .Y(n_964) );
INVx1_ASAP7_75t_L g1109 ( .A(n_928), .Y(n_1109) );
INVx1_ASAP7_75t_L g1032 ( .A(n_944), .Y(n_1032) );
INVx1_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
XNOR2x1_ASAP7_75t_L g945 ( .A(n_946), .B(n_992), .Y(n_945) );
NAND3xp33_ASAP7_75t_L g948 ( .A(n_949), .B(n_954), .C(n_957), .Y(n_948) );
NAND4xp25_ASAP7_75t_L g960 ( .A(n_961), .B(n_966), .C(n_970), .D(n_976), .Y(n_960) );
INVx1_ASAP7_75t_L g1074 ( .A(n_973), .Y(n_1074) );
AND4x1_ASAP7_75t_L g993 ( .A(n_994), .B(n_1006), .C(n_1014), .D(n_1019), .Y(n_993) );
NAND4xp25_ASAP7_75t_L g1031 ( .A(n_994), .B(n_1006), .C(n_1014), .D(n_1019), .Y(n_1031) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_997), .B(n_998), .Y(n_996) );
INVx2_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1939 ( .A(n_999), .Y(n_1939) );
INVx2_ASAP7_75t_SL g1314 ( .A(n_1033), .Y(n_1314) );
AO22x2_ASAP7_75t_L g1033 ( .A1(n_1034), .A2(n_1035), .B1(n_1162), .B2(n_1312), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
AO22x1_ASAP7_75t_L g1035 ( .A1(n_1036), .A2(n_1110), .B1(n_1160), .B2(n_1161), .Y(n_1035) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1036), .Y(n_1161) );
AND4x1_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1065), .C(n_1067), .D(n_1102), .Y(n_1037) );
NOR3xp33_ASAP7_75t_SL g1038 ( .A(n_1039), .B(n_1040), .C(n_1043), .Y(n_1038) );
NOR3xp33_ASAP7_75t_SL g1321 ( .A(n_1039), .B(n_1322), .C(n_1337), .Y(n_1321) );
NOR3xp33_ASAP7_75t_SL g1621 ( .A(n_1039), .B(n_1622), .C(n_1631), .Y(n_1621) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
OAI221xp5_ASAP7_75t_L g1323 ( .A1(n_1045), .A2(n_1056), .B1(n_1324), .B2(n_1325), .C(n_1326), .Y(n_1323) );
OAI221xp5_ASAP7_75t_L g1623 ( .A1(n_1045), .A2(n_1056), .B1(n_1624), .B2(n_1625), .C(n_1626), .Y(n_1623) );
BUFx2_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
INVx2_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
CKINVDCx5p33_ASAP7_75t_R g1051 ( .A(n_1052), .Y(n_1051) );
AOI33xp33_ASAP7_75t_L g1523 ( .A1(n_1052), .A2(n_1524), .A3(n_1525), .B1(n_1527), .B2(n_1529), .B3(n_1530), .Y(n_1523) );
OAI221xp5_ASAP7_75t_L g1053 ( .A1(n_1054), .A2(n_1055), .B1(n_1056), .B2(n_1059), .C(n_1060), .Y(n_1053) );
OAI221xp5_ASAP7_75t_L g1329 ( .A1(n_1054), .A2(n_1330), .B1(n_1331), .B2(n_1333), .C(n_1334), .Y(n_1329) );
OAI221xp5_ASAP7_75t_L g1627 ( .A1(n_1054), .A2(n_1586), .B1(n_1628), .B2(n_1629), .C(n_1630), .Y(n_1627) );
BUFx2_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1058), .Y(n_1232) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1058), .Y(n_1586) );
BUFx3_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1062), .Y(n_1336) );
BUFx2_ASAP7_75t_L g1391 ( .A(n_1062), .Y(n_1391) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1064), .Y(n_1119) );
OAI31xp33_ASAP7_75t_L g1067 ( .A1(n_1068), .A2(n_1084), .A3(n_1098), .B(n_1101), .Y(n_1067) );
OAI221xp5_ASAP7_75t_L g1069 ( .A1(n_1070), .A2(n_1073), .B1(n_1074), .B2(n_1075), .C(n_1076), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
INVx2_ASAP7_75t_L g1345 ( .A(n_1071), .Y(n_1345) );
INVx2_ASAP7_75t_L g1356 ( .A(n_1071), .Y(n_1356) );
INVx2_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
BUFx2_ASAP7_75t_L g1136 ( .A(n_1072), .Y(n_1136) );
OAI221xp5_ASAP7_75t_L g1643 ( .A1(n_1074), .A2(n_1356), .B1(n_1644), .B2(n_1645), .C(n_1646), .Y(n_1643) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_1079), .A2(n_1080), .B1(n_1082), .B2(n_1083), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1144 ( .A1(n_1080), .A2(n_1083), .B1(n_1115), .B2(n_1116), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g1479 ( .A1(n_1080), .A2(n_1083), .B1(n_1480), .B2(n_1481), .Y(n_1479) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_1083), .A2(n_1361), .B1(n_1362), .B2(n_1363), .Y(n_1360) );
AOI22xp5_ASAP7_75t_L g1521 ( .A1(n_1083), .A2(n_1362), .B1(n_1495), .B2(n_1496), .Y(n_1521) );
AOI22xp33_ASAP7_75t_L g1609 ( .A1(n_1083), .A2(n_1362), .B1(n_1610), .B2(n_1611), .Y(n_1609) );
AOI22xp33_ASAP7_75t_L g1647 ( .A1(n_1083), .A2(n_1362), .B1(n_1648), .B2(n_1649), .Y(n_1647) );
AOI22xp33_ASAP7_75t_L g1915 ( .A1(n_1083), .A2(n_1362), .B1(n_1916), .B2(n_1917), .Y(n_1915) );
OAI221xp5_ASAP7_75t_L g1146 ( .A1(n_1087), .A2(n_1147), .B1(n_1148), .B2(n_1149), .C(n_1151), .Y(n_1146) );
OAI22xp5_ASAP7_75t_L g1088 ( .A1(n_1089), .A2(n_1092), .B1(n_1093), .B2(n_1096), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
CKINVDCx5p33_ASAP7_75t_R g1093 ( .A(n_1094), .Y(n_1093) );
BUFx3_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
AND2x4_ASAP7_75t_L g1170 ( .A(n_1095), .B(n_1171), .Y(n_1170) );
OAI31xp33_ASAP7_75t_SL g1341 ( .A1(n_1101), .A2(n_1342), .A3(n_1343), .B(n_1354), .Y(n_1341) );
CKINVDCx8_ASAP7_75t_R g1483 ( .A(n_1101), .Y(n_1483) );
NOR2xp33_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1105), .Y(n_1102) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1110), .Y(n_1160) );
AND3x1_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1131), .C(n_1133), .Y(n_1111) );
NOR2xp33_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1124), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1128), .Y(n_1124) );
OAI221xp5_ASAP7_75t_L g1135 ( .A1(n_1126), .A2(n_1130), .B1(n_1136), .B2(n_1137), .C(n_1140), .Y(n_1135) );
OAI31xp33_ASAP7_75t_L g1133 ( .A1(n_1134), .A2(n_1145), .A3(n_1157), .B(n_1158), .Y(n_1133) );
OAI22xp5_ASAP7_75t_L g1919 ( .A1(n_1136), .A2(n_1920), .B1(n_1921), .B2(n_1923), .Y(n_1919) );
OAI221xp5_ASAP7_75t_L g1355 ( .A1(n_1137), .A2(n_1356), .B1(n_1357), .B2(n_1358), .C(n_1359), .Y(n_1355) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
AND2x4_ASAP7_75t_L g1177 ( .A(n_1143), .B(n_1171), .Y(n_1177) );
BUFx3_ASAP7_75t_L g1282 ( .A(n_1143), .Y(n_1282) );
BUFx2_ASAP7_75t_L g1547 ( .A(n_1143), .Y(n_1547) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
INVx2_ASAP7_75t_L g1421 ( .A(n_1150), .Y(n_1421) );
OAI22xp5_ASAP7_75t_L g1152 ( .A1(n_1153), .A2(n_1154), .B1(n_1155), .B2(n_1156), .Y(n_1152) );
OAI31xp33_ASAP7_75t_L g1503 ( .A1(n_1158), .A2(n_1504), .A3(n_1512), .B(n_1522), .Y(n_1503) );
OAI31xp33_ASAP7_75t_L g1595 ( .A1(n_1158), .A2(n_1596), .A3(n_1597), .B(n_1604), .Y(n_1595) );
BUFx8_ASAP7_75t_SL g1158 ( .A(n_1159), .Y(n_1158) );
INVx2_ASAP7_75t_L g1373 ( .A(n_1159), .Y(n_1373) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1162), .Y(n_1312) );
AOI22x1_ASAP7_75t_L g1162 ( .A1(n_1163), .A2(n_1256), .B1(n_1309), .B2(n_1310), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1165), .B(n_1212), .Y(n_1164) );
NOR3xp33_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1180), .C(n_1190), .Y(n_1165) );
NAND2xp5_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1175), .Y(n_1166) );
AOI22xp33_ASAP7_75t_L g1167 ( .A1(n_1168), .A2(n_1169), .B1(n_1172), .B2(n_1173), .Y(n_1167) );
BUFx2_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
BUFx2_ASAP7_75t_L g1409 ( .A(n_1170), .Y(n_1409) );
AND2x6_ASAP7_75t_L g1173 ( .A(n_1171), .B(n_1174), .Y(n_1173) );
OAI221xp5_ASAP7_75t_L g1231 ( .A1(n_1172), .A2(n_1176), .B1(n_1232), .B2(n_1233), .C(n_1234), .Y(n_1231) );
AOI22xp33_ASAP7_75t_L g1407 ( .A1(n_1173), .A2(n_1408), .B1(n_1409), .B2(n_1410), .Y(n_1407) );
NAND2x1p5_ASAP7_75t_L g1189 ( .A(n_1174), .B(n_1184), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_1176), .A2(n_1177), .B1(n_1178), .B2(n_1179), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g1411 ( .A1(n_1177), .A2(n_1412), .B1(n_1413), .B2(n_1414), .Y(n_1411) );
INVx2_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
INVx2_ASAP7_75t_SL g1416 ( .A(n_1182), .Y(n_1416) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
INVx3_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
BUFx4f_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
BUFx2_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
OAI22xp33_ASAP7_75t_L g1191 ( .A1(n_1192), .A2(n_1195), .B1(n_1196), .B2(n_1198), .Y(n_1191) );
OAI22xp33_ASAP7_75t_L g1208 ( .A1(n_1192), .A2(n_1209), .B1(n_1210), .B2(n_1211), .Y(n_1208) );
OAI22xp33_ASAP7_75t_L g1432 ( .A1(n_1192), .A2(n_1399), .B1(n_1401), .B2(n_1433), .Y(n_1432) );
BUFx2_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
INVx2_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1197), .Y(n_1210) );
OAI22xp5_ASAP7_75t_L g1199 ( .A1(n_1200), .A2(n_1201), .B1(n_1202), .B2(n_1203), .Y(n_1199) );
OAI22xp5_ASAP7_75t_L g1204 ( .A1(n_1201), .A2(n_1205), .B1(n_1206), .B2(n_1207), .Y(n_1204) );
OAI22xp5_ASAP7_75t_L g1425 ( .A1(n_1203), .A2(n_1426), .B1(n_1429), .B2(n_1430), .Y(n_1425) );
OAI22xp5_ASAP7_75t_L g1911 ( .A1(n_1203), .A2(n_1912), .B1(n_1913), .B2(n_1914), .Y(n_1911) );
AOI211xp5_ASAP7_75t_L g1219 ( .A1(n_1205), .A2(n_1220), .B(n_1222), .C(n_1228), .Y(n_1219) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1206), .Y(n_1284) );
AOI22xp33_ASAP7_75t_L g1249 ( .A1(n_1207), .A2(n_1209), .B1(n_1250), .B2(n_1252), .Y(n_1249) );
AOI221xp5_ASAP7_75t_L g1236 ( .A1(n_1211), .A2(n_1237), .B1(n_1240), .B2(n_1244), .C(n_1247), .Y(n_1236) );
AOI21xp5_ASAP7_75t_L g1212 ( .A1(n_1213), .A2(n_1217), .B(n_1218), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
INVx5_ASAP7_75t_L g1404 ( .A(n_1214), .Y(n_1404) );
AND2x4_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1216), .Y(n_1214) );
AOI31xp33_ASAP7_75t_L g1218 ( .A1(n_1219), .A2(n_1236), .A3(n_1249), .B(n_1254), .Y(n_1218) );
AOI221xp5_ASAP7_75t_L g1375 ( .A1(n_1220), .A2(n_1376), .B1(n_1380), .B2(n_1384), .C(n_1385), .Y(n_1375) );
INVx2_ASAP7_75t_SL g1223 ( .A(n_1224), .Y(n_1223) );
INVx2_ASAP7_75t_L g1386 ( .A(n_1224), .Y(n_1386) );
INVx1_ASAP7_75t_SL g1248 ( .A(n_1227), .Y(n_1248) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
OAI221xp5_ASAP7_75t_L g1584 ( .A1(n_1233), .A2(n_1585), .B1(n_1586), .B2(n_1587), .C(n_1588), .Y(n_1584) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
BUFx2_ASAP7_75t_L g1379 ( .A(n_1235), .Y(n_1379) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
BUFx6f_ASAP7_75t_L g1398 ( .A(n_1239), .Y(n_1398) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1243), .Y(n_1395) );
INVx2_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
AOI221xp5_ASAP7_75t_L g1389 ( .A1(n_1247), .A2(n_1390), .B1(n_1396), .B2(n_1398), .C(n_1399), .Y(n_1389) );
AOI22xp33_ASAP7_75t_L g1400 ( .A1(n_1250), .A2(n_1252), .B1(n_1401), .B2(n_1402), .Y(n_1400) );
INVx6_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
INVx4_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
INVx2_ASAP7_75t_L g1309 ( .A(n_1256), .Y(n_1309) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1258), .Y(n_1308) );
AOI211x1_ASAP7_75t_L g1258 ( .A1(n_1259), .A2(n_1270), .B(n_1272), .C(n_1299), .Y(n_1258) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1272 ( .A(n_1273), .B(n_1286), .Y(n_1272) );
INVx2_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
BUFx3_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
HB1xp67_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
BUFx3_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
INVx2_ASAP7_75t_SL g1453 ( .A(n_1289), .Y(n_1453) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
INVx3_ASAP7_75t_SL g1310 ( .A(n_1311), .Y(n_1310) );
AOI22xp5_ASAP7_75t_L g1315 ( .A1(n_1316), .A2(n_1575), .B1(n_1576), .B2(n_1655), .Y(n_1315) );
INVx1_ASAP7_75t_SL g1655 ( .A(n_1316), .Y(n_1655) );
XNOR2xp5_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1488), .Y(n_1316) );
XOR2xp5_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1367), .Y(n_1317) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
AND4x1_ASAP7_75t_L g1320 ( .A(n_1321), .B(n_1339), .C(n_1341), .D(n_1364), .Y(n_1320) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
OAI22xp33_ASAP7_75t_L g1443 ( .A1(n_1328), .A2(n_1336), .B1(n_1444), .B2(n_1445), .Y(n_1443) );
INVx2_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
OAI22xp5_ASAP7_75t_L g1344 ( .A1(n_1345), .A2(n_1346), .B1(n_1347), .B2(n_1350), .Y(n_1344) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
OAI221xp5_ASAP7_75t_L g1635 ( .A1(n_1352), .A2(n_1624), .B1(n_1625), .B2(n_1636), .C(n_1637), .Y(n_1635) );
INVx2_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
NOR2xp33_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1366), .Y(n_1364) );
AOI22xp5_ASAP7_75t_L g1367 ( .A1(n_1368), .A2(n_1435), .B1(n_1436), .B2(n_1487), .Y(n_1367) );
INVx2_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
HB1xp67_ASAP7_75t_L g1487 ( .A(n_1369), .Y(n_1487) );
XNOR2x1_ASAP7_75t_L g1369 ( .A(n_1370), .B(n_1371), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1372), .B(n_1405), .Y(n_1371) );
AOI22xp33_ASAP7_75t_L g1372 ( .A1(n_1373), .A2(n_1374), .B1(n_1403), .B2(n_1404), .Y(n_1372) );
NAND3xp33_ASAP7_75t_L g1374 ( .A(n_1375), .B(n_1389), .C(n_1400), .Y(n_1374) );
HB1xp67_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
INVx2_ASAP7_75t_SL g1387 ( .A(n_1388), .Y(n_1387) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
NOR3xp33_ASAP7_75t_SL g1405 ( .A(n_1406), .B(n_1415), .C(n_1417), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1411), .Y(n_1406) );
OAI33xp33_ASAP7_75t_L g1417 ( .A1(n_1418), .A2(n_1420), .A3(n_1425), .B1(n_1431), .B2(n_1432), .B3(n_1434), .Y(n_1417) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
OAI22xp33_ASAP7_75t_L g1420 ( .A1(n_1421), .A2(n_1422), .B1(n_1423), .B2(n_1424), .Y(n_1420) );
INVx2_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
INVx2_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
OAI21xp33_ASAP7_75t_L g1602 ( .A1(n_1433), .A2(n_1587), .B(n_1603), .Y(n_1602) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
AND4x1_ASAP7_75t_L g1439 ( .A(n_1440), .B(n_1459), .C(n_1461), .D(n_1484), .Y(n_1439) );
NOR3xp33_ASAP7_75t_SL g1440 ( .A(n_1441), .B(n_1442), .C(n_1456), .Y(n_1440) );
OAI22xp5_ASAP7_75t_L g1464 ( .A1(n_1444), .A2(n_1445), .B1(n_1465), .B2(n_1466), .Y(n_1464) );
OAI31xp33_ASAP7_75t_L g1461 ( .A1(n_1462), .A2(n_1463), .A3(n_1470), .B(n_1482), .Y(n_1461) );
OAI22xp5_ASAP7_75t_SL g1475 ( .A1(n_1465), .A2(n_1476), .B1(n_1477), .B2(n_1478), .Y(n_1475) );
OAI22xp5_ASAP7_75t_L g1598 ( .A1(n_1465), .A2(n_1599), .B1(n_1600), .B2(n_1601), .Y(n_1598) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
OAI221xp5_ASAP7_75t_L g1907 ( .A1(n_1474), .A2(n_1637), .B1(n_1908), .B2(n_1909), .C(n_1910), .Y(n_1907) );
INVx2_ASAP7_75t_L g1482 ( .A(n_1483), .Y(n_1482) );
AOI31xp33_ASAP7_75t_SL g1536 ( .A1(n_1483), .A2(n_1537), .A3(n_1542), .B(n_1545), .Y(n_1536) );
NOR2xp33_ASAP7_75t_L g1484 ( .A(n_1485), .B(n_1486), .Y(n_1484) );
HB1xp67_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
AOI22xp5_ASAP7_75t_L g1489 ( .A1(n_1490), .A2(n_1491), .B1(n_1532), .B2(n_1533), .Y(n_1489) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
NAND4xp75_ASAP7_75t_SL g1492 ( .A(n_1493), .B(n_1501), .C(n_1503), .D(n_1523), .Y(n_1492) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1494), .B(n_1497), .Y(n_1493) );
OAI22xp5_ASAP7_75t_L g1515 ( .A1(n_1498), .A2(n_1516), .B1(n_1518), .B2(n_1520), .Y(n_1515) );
BUFx2_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
AOI33xp33_ASAP7_75t_L g1935 ( .A1(n_1524), .A2(n_1936), .A3(n_1938), .B1(n_1940), .B2(n_1941), .B3(n_1942), .Y(n_1935) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
XNOR2xp5_ASAP7_75t_L g1533 ( .A(n_1534), .B(n_1535), .Y(n_1533) );
OAI22xp5_ASAP7_75t_L g1725 ( .A1(n_1534), .A2(n_1695), .B1(n_1726), .B2(n_1727), .Y(n_1725) );
NOR4xp75_ASAP7_75t_L g1535 ( .A(n_1536), .B(n_1550), .C(n_1557), .D(n_1559), .Y(n_1535) );
NAND2xp5_ASAP7_75t_L g1550 ( .A(n_1551), .B(n_1554), .Y(n_1550) );
NAND3xp33_ASAP7_75t_SL g1559 ( .A(n_1560), .B(n_1562), .C(n_1566), .Y(n_1559) );
NAND3xp33_ASAP7_75t_SL g1932 ( .A(n_1560), .B(n_1933), .C(n_1935), .Y(n_1932) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
AOI22xp5_ASAP7_75t_L g1576 ( .A1(n_1577), .A2(n_1615), .B1(n_1653), .B2(n_1654), .Y(n_1576) );
INVx1_ASAP7_75t_L g1653 ( .A(n_1577), .Y(n_1653) );
HB1xp67_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
AND4x1_ASAP7_75t_L g1579 ( .A(n_1580), .B(n_1582), .C(n_1595), .D(n_1612), .Y(n_1579) );
NOR2xp33_ASAP7_75t_L g1612 ( .A(n_1613), .B(n_1614), .Y(n_1612) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1615), .Y(n_1654) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1616), .Y(n_1615) );
XNOR2xp5_ASAP7_75t_L g1616 ( .A(n_1617), .B(n_1618), .Y(n_1616) );
AND4x1_ASAP7_75t_L g1618 ( .A(n_1619), .B(n_1621), .C(n_1632), .D(n_1650), .Y(n_1618) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
NOR2xp33_ASAP7_75t_L g1650 ( .A(n_1651), .B(n_1652), .Y(n_1650) );
OAI221xp5_ASAP7_75t_SL g1656 ( .A1(n_1657), .A2(n_1899), .B1(n_1902), .B2(n_1947), .C(n_1952), .Y(n_1656) );
AND4x1_ASAP7_75t_L g1657 ( .A(n_1658), .B(n_1826), .C(n_1840), .D(n_1872), .Y(n_1657) );
AOI211xp5_ASAP7_75t_L g1658 ( .A1(n_1659), .A2(n_1687), .B(n_1788), .C(n_1802), .Y(n_1658) );
NAND2xp5_ASAP7_75t_L g1803 ( .A(n_1659), .B(n_1804), .Y(n_1803) );
NAND2xp5_ASAP7_75t_L g1849 ( .A(n_1659), .B(n_1761), .Y(n_1849) );
AOI221xp5_ASAP7_75t_L g1867 ( .A1(n_1659), .A2(n_1737), .B1(n_1765), .B2(n_1868), .C(n_1869), .Y(n_1867) );
OAI333xp33_ASAP7_75t_L g1891 ( .A1(n_1659), .A2(n_1735), .A3(n_1793), .B1(n_1828), .B2(n_1892), .B3(n_1894), .C1(n_1895), .C2(n_1897), .C3(n_1898), .Y(n_1891) );
CKINVDCx5p33_ASAP7_75t_R g1659 ( .A(n_1660), .Y(n_1659) );
NAND2xp5_ASAP7_75t_L g1828 ( .A(n_1660), .B(n_1795), .Y(n_1828) );
OAI32xp33_ASAP7_75t_L g1848 ( .A1(n_1660), .A2(n_1700), .A3(n_1761), .B1(n_1820), .B2(n_1849), .Y(n_1848) );
INVx1_ASAP7_75t_L g1882 ( .A(n_1660), .Y(n_1882) );
NAND2xp5_ASAP7_75t_L g1897 ( .A(n_1660), .B(n_1720), .Y(n_1897) );
OR2x6_ASAP7_75t_SL g1660 ( .A(n_1661), .B(n_1673), .Y(n_1660) );
OAI22xp5_ASAP7_75t_L g1661 ( .A1(n_1662), .A2(n_1663), .B1(n_1670), .B2(n_1671), .Y(n_1661) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
INVx1_ASAP7_75t_L g1726 ( .A(n_1664), .Y(n_1726) );
BUFx3_ASAP7_75t_L g1901 ( .A(n_1664), .Y(n_1901) );
AND2x4_ASAP7_75t_L g1664 ( .A(n_1665), .B(n_1668), .Y(n_1664) );
AND2x2_ASAP7_75t_L g1694 ( .A(n_1665), .B(n_1668), .Y(n_1694) );
HB1xp67_ASAP7_75t_L g1964 ( .A(n_1665), .Y(n_1964) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1666), .Y(n_1665) );
AND2x4_ASAP7_75t_L g1672 ( .A(n_1666), .B(n_1668), .Y(n_1672) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
NAND2xp5_ASAP7_75t_L g1679 ( .A(n_1667), .B(n_1680), .Y(n_1679) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1669), .Y(n_1680) );
INVx2_ASAP7_75t_L g1710 ( .A(n_1671), .Y(n_1710) );
INVx2_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
INVx1_ASAP7_75t_SL g1695 ( .A(n_1672), .Y(n_1695) );
OAI22xp5_ASAP7_75t_L g1673 ( .A1(n_1674), .A2(n_1675), .B1(n_1681), .B2(n_1682), .Y(n_1673) );
BUFx3_ASAP7_75t_L g1675 ( .A(n_1676), .Y(n_1675) );
OAI22xp5_ASAP7_75t_L g1697 ( .A1(n_1676), .A2(n_1685), .B1(n_1698), .B2(n_1699), .Y(n_1697) );
OAI22xp33_ASAP7_75t_L g1722 ( .A1(n_1676), .A2(n_1683), .B1(n_1723), .B2(n_1724), .Y(n_1722) );
OAI22xp33_ASAP7_75t_L g1739 ( .A1(n_1676), .A2(n_1685), .B1(n_1740), .B2(n_1741), .Y(n_1739) );
BUFx6f_ASAP7_75t_L g1676 ( .A(n_1677), .Y(n_1676) );
OAI22xp5_ASAP7_75t_L g1716 ( .A1(n_1677), .A2(n_1685), .B1(n_1717), .B2(n_1718), .Y(n_1716) );
OR2x2_ASAP7_75t_L g1677 ( .A(n_1678), .B(n_1679), .Y(n_1677) );
OR2x2_ASAP7_75t_L g1685 ( .A(n_1678), .B(n_1686), .Y(n_1685) );
INVx1_ASAP7_75t_L g1706 ( .A(n_1678), .Y(n_1706) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1679), .Y(n_1705) );
HB1xp67_ASAP7_75t_L g1963 ( .A(n_1680), .Y(n_1963) );
HB1xp67_ASAP7_75t_L g1682 ( .A(n_1683), .Y(n_1682) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1686), .Y(n_1708) );
NAND5xp2_ASAP7_75t_L g1687 ( .A(n_1688), .B(n_1756), .C(n_1769), .D(n_1777), .E(n_1781), .Y(n_1687) );
AOI211xp5_ASAP7_75t_SL g1688 ( .A1(n_1689), .A2(n_1719), .B(n_1731), .C(n_1752), .Y(n_1688) );
INVx1_ASAP7_75t_L g1838 ( .A(n_1689), .Y(n_1838) );
AND2x2_ASAP7_75t_L g1689 ( .A(n_1690), .B(n_1700), .Y(n_1689) );
AND2x2_ASAP7_75t_L g1733 ( .A(n_1690), .B(n_1734), .Y(n_1733) );
AND2x2_ASAP7_75t_L g1751 ( .A(n_1690), .B(n_1735), .Y(n_1751) );
AND2x2_ASAP7_75t_L g1768 ( .A(n_1690), .B(n_1702), .Y(n_1768) );
NOR2xp33_ASAP7_75t_L g1780 ( .A(n_1690), .B(n_1702), .Y(n_1780) );
NAND2xp5_ASAP7_75t_L g1811 ( .A(n_1690), .B(n_1812), .Y(n_1811) );
AND2x2_ASAP7_75t_L g1823 ( .A(n_1690), .B(n_1746), .Y(n_1823) );
OR2x2_ASAP7_75t_L g1825 ( .A(n_1690), .B(n_1746), .Y(n_1825) );
AND2x2_ASAP7_75t_L g1847 ( .A(n_1690), .B(n_1745), .Y(n_1847) );
AND2x2_ASAP7_75t_L g1852 ( .A(n_1690), .B(n_1711), .Y(n_1852) );
NOR2xp33_ASAP7_75t_L g1863 ( .A(n_1690), .B(n_1763), .Y(n_1863) );
NOR2xp33_ASAP7_75t_L g1893 ( .A(n_1690), .B(n_1715), .Y(n_1893) );
CKINVDCx6p67_ASAP7_75t_R g1690 ( .A(n_1691), .Y(n_1690) );
OR2x2_ASAP7_75t_L g1783 ( .A(n_1691), .B(n_1735), .Y(n_1783) );
AND2x2_ASAP7_75t_L g1806 ( .A(n_1691), .B(n_1770), .Y(n_1806) );
AND2x2_ASAP7_75t_L g1818 ( .A(n_1691), .B(n_1735), .Y(n_1818) );
AND2x2_ASAP7_75t_L g1820 ( .A(n_1691), .B(n_1711), .Y(n_1820) );
NAND2xp5_ASAP7_75t_L g1832 ( .A(n_1691), .B(n_1833), .Y(n_1832) );
AND2x2_ASAP7_75t_L g1836 ( .A(n_1691), .B(n_1734), .Y(n_1836) );
AND2x2_ASAP7_75t_L g1866 ( .A(n_1691), .B(n_1745), .Y(n_1866) );
OR2x2_ASAP7_75t_L g1875 ( .A(n_1691), .B(n_1771), .Y(n_1875) );
OR2x6_ASAP7_75t_SL g1691 ( .A(n_1692), .B(n_1697), .Y(n_1691) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1694), .Y(n_1693) );
AND2x2_ASAP7_75t_L g1700 ( .A(n_1701), .B(n_1711), .Y(n_1700) );
NAND2xp5_ASAP7_75t_L g1732 ( .A(n_1701), .B(n_1733), .Y(n_1732) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1701), .Y(n_1744) );
NOR2xp33_ASAP7_75t_L g1796 ( .A(n_1701), .B(n_1797), .Y(n_1796) );
NOR2xp33_ASAP7_75t_L g1833 ( .A(n_1701), .B(n_1771), .Y(n_1833) );
INVx4_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1750 ( .A(n_1702), .B(n_1751), .Y(n_1750) );
NAND2xp5_ASAP7_75t_L g1763 ( .A(n_1702), .B(n_1711), .Y(n_1763) );
INVx2_ASAP7_75t_L g1775 ( .A(n_1702), .Y(n_1775) );
AND2x2_ASAP7_75t_L g1812 ( .A(n_1702), .B(n_1721), .Y(n_1812) );
OR2x2_ASAP7_75t_L g1859 ( .A(n_1702), .B(n_1786), .Y(n_1859) );
NAND2xp5_ASAP7_75t_L g1865 ( .A(n_1702), .B(n_1866), .Y(n_1865) );
OR2x2_ASAP7_75t_L g1870 ( .A(n_1702), .B(n_1771), .Y(n_1870) );
OR2x2_ASAP7_75t_L g1874 ( .A(n_1702), .B(n_1875), .Y(n_1874) );
NAND2xp5_ASAP7_75t_L g1894 ( .A(n_1702), .B(n_1787), .Y(n_1894) );
AND2x2_ASAP7_75t_L g1896 ( .A(n_1702), .B(n_1765), .Y(n_1896) );
AND2x6_ASAP7_75t_L g1702 ( .A(n_1703), .B(n_1709), .Y(n_1702) );
AND2x4_ASAP7_75t_L g1704 ( .A(n_1705), .B(n_1706), .Y(n_1704) );
AND2x4_ASAP7_75t_L g1707 ( .A(n_1706), .B(n_1708), .Y(n_1707) );
AND2x2_ASAP7_75t_L g1711 ( .A(n_1712), .B(n_1715), .Y(n_1711) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1712), .Y(n_1735) );
AND2x2_ASAP7_75t_L g1745 ( .A(n_1712), .B(n_1746), .Y(n_1745) );
OR2x2_ASAP7_75t_L g1771 ( .A(n_1712), .B(n_1715), .Y(n_1771) );
AND2x2_ASAP7_75t_L g1712 ( .A(n_1713), .B(n_1714), .Y(n_1712) );
AND2x2_ASAP7_75t_L g1734 ( .A(n_1715), .B(n_1735), .Y(n_1734) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1715), .Y(n_1746) );
NAND2xp5_ASAP7_75t_L g1800 ( .A(n_1719), .B(n_1801), .Y(n_1800) );
AND2x2_ASAP7_75t_L g1879 ( .A(n_1719), .B(n_1868), .Y(n_1879) );
AND2x2_ASAP7_75t_L g1719 ( .A(n_1720), .B(n_1728), .Y(n_1719) );
AND2x2_ASAP7_75t_L g1747 ( .A(n_1720), .B(n_1737), .Y(n_1747) );
AND2x2_ASAP7_75t_L g1748 ( .A(n_1720), .B(n_1749), .Y(n_1748) );
AND2x2_ASAP7_75t_L g1760 ( .A(n_1720), .B(n_1761), .Y(n_1760) );
OR2x2_ASAP7_75t_L g1793 ( .A(n_1720), .B(n_1728), .Y(n_1793) );
INVx3_ASAP7_75t_L g1795 ( .A(n_1720), .Y(n_1795) );
AOI21xp5_ASAP7_75t_L g1887 ( .A1(n_1720), .A2(n_1888), .B(n_1891), .Y(n_1887) );
INVx3_ASAP7_75t_L g1720 ( .A(n_1721), .Y(n_1720) );
OR2x2_ASAP7_75t_L g1754 ( .A(n_1721), .B(n_1755), .Y(n_1754) );
AND2x2_ASAP7_75t_L g1886 ( .A(n_1721), .B(n_1728), .Y(n_1886) );
OR2x2_ASAP7_75t_L g1721 ( .A(n_1722), .B(n_1725), .Y(n_1721) );
AND2x2_ASAP7_75t_L g1737 ( .A(n_1728), .B(n_1738), .Y(n_1737) );
OR2x2_ASAP7_75t_L g1755 ( .A(n_1728), .B(n_1738), .Y(n_1755) );
INVx2_ASAP7_75t_L g1761 ( .A(n_1728), .Y(n_1761) );
AND2x2_ASAP7_75t_L g1765 ( .A(n_1728), .B(n_1749), .Y(n_1765) );
OR2x2_ASAP7_75t_L g1776 ( .A(n_1728), .B(n_1749), .Y(n_1776) );
AOI22xp5_ASAP7_75t_L g1829 ( .A1(n_1728), .A2(n_1797), .B1(n_1830), .B2(n_1834), .Y(n_1829) );
OAI221xp5_ASAP7_75t_L g1856 ( .A1(n_1728), .A2(n_1855), .B1(n_1857), .B2(n_1865), .C(n_1867), .Y(n_1856) );
AND2x4_ASAP7_75t_L g1728 ( .A(n_1729), .B(n_1730), .Y(n_1728) );
OAI21xp5_ASAP7_75t_SL g1731 ( .A1(n_1732), .A2(n_1736), .B(n_1742), .Y(n_1731) );
NAND2xp5_ASAP7_75t_L g1794 ( .A(n_1733), .B(n_1795), .Y(n_1794) );
A2O1A1Ixp33_ASAP7_75t_SL g1826 ( .A1(n_1733), .A2(n_1827), .B(n_1829), .C(n_1837), .Y(n_1826) );
AOI211xp5_ASAP7_75t_L g1857 ( .A1(n_1733), .A2(n_1858), .B(n_1860), .C(n_1864), .Y(n_1857) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1734), .Y(n_1753) );
NAND2xp5_ASAP7_75t_L g1767 ( .A(n_1734), .B(n_1768), .Y(n_1767) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1737), .Y(n_1736) );
AOI322xp5_ASAP7_75t_L g1807 ( .A1(n_1737), .A2(n_1760), .A3(n_1808), .B1(n_1810), .B2(n_1813), .C1(n_1816), .C2(n_1821), .Y(n_1807) );
INVx2_ASAP7_75t_SL g1749 ( .A(n_1738), .Y(n_1749) );
HB1xp67_ASAP7_75t_L g1759 ( .A(n_1738), .Y(n_1759) );
AOI22xp5_ASAP7_75t_L g1742 ( .A1(n_1743), .A2(n_1747), .B1(n_1748), .B2(n_1750), .Y(n_1742) );
INVxp67_ASAP7_75t_L g1898 ( .A(n_1743), .Y(n_1898) );
AND2x2_ASAP7_75t_L g1743 ( .A(n_1744), .B(n_1745), .Y(n_1743) );
INVx1_ASAP7_75t_L g1809 ( .A(n_1745), .Y(n_1809) );
NOR2xp33_ASAP7_75t_L g1892 ( .A(n_1745), .B(n_1893), .Y(n_1892) );
INVx1_ASAP7_75t_L g1876 ( .A(n_1748), .Y(n_1876) );
INVx2_ASAP7_75t_SL g1787 ( .A(n_1749), .Y(n_1787) );
NOR2xp33_ASAP7_75t_L g1752 ( .A(n_1753), .B(n_1754), .Y(n_1752) );
AND2x2_ASAP7_75t_L g1808 ( .A(n_1753), .B(n_1809), .Y(n_1808) );
INVx1_ASAP7_75t_L g1821 ( .A(n_1754), .Y(n_1821) );
INVx1_ASAP7_75t_L g1839 ( .A(n_1755), .Y(n_1839) );
OAI21xp33_ASAP7_75t_SL g1850 ( .A1(n_1755), .A2(n_1851), .B(n_1853), .Y(n_1850) );
AOI21xp5_ASAP7_75t_L g1756 ( .A1(n_1757), .A2(n_1762), .B(n_1764), .Y(n_1756) );
INVx1_ASAP7_75t_L g1757 ( .A(n_1758), .Y(n_1757) );
NAND2xp5_ASAP7_75t_L g1758 ( .A(n_1759), .B(n_1760), .Y(n_1758) );
INVx1_ASAP7_75t_L g1790 ( .A(n_1759), .Y(n_1790) );
NAND2xp5_ASAP7_75t_L g1805 ( .A(n_1759), .B(n_1806), .Y(n_1805) );
NAND2xp5_ASAP7_75t_L g1834 ( .A(n_1759), .B(n_1835), .Y(n_1834) );
INVx1_ASAP7_75t_L g1855 ( .A(n_1759), .Y(n_1855) );
INVx1_ASAP7_75t_L g1862 ( .A(n_1759), .Y(n_1862) );
AOI211xp5_ASAP7_75t_SL g1877 ( .A1(n_1760), .A2(n_1878), .B(n_1879), .C(n_1880), .Y(n_1877) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1763), .Y(n_1762) );
A2O1A1Ixp33_ASAP7_75t_L g1873 ( .A1(n_1763), .A2(n_1874), .B(n_1876), .C(n_1877), .Y(n_1873) );
AND2x2_ASAP7_75t_L g1764 ( .A(n_1765), .B(n_1766), .Y(n_1764) );
NAND2xp5_ASAP7_75t_L g1777 ( .A(n_1765), .B(n_1778), .Y(n_1777) );
AOI21xp5_ASAP7_75t_L g1837 ( .A1(n_1765), .A2(n_1838), .B(n_1839), .Y(n_1837) );
INVx1_ASAP7_75t_L g1843 ( .A(n_1765), .Y(n_1843) );
INVx1_ASAP7_75t_L g1766 ( .A(n_1767), .Y(n_1766) );
NOR2xp33_ASAP7_75t_L g1799 ( .A(n_1767), .B(n_1800), .Y(n_1799) );
NAND2xp5_ASAP7_75t_L g1792 ( .A(n_1768), .B(n_1770), .Y(n_1792) );
NAND2xp5_ASAP7_75t_L g1769 ( .A(n_1770), .B(n_1772), .Y(n_1769) );
NAND2xp5_ASAP7_75t_L g1779 ( .A(n_1770), .B(n_1780), .Y(n_1779) );
INVx1_ASAP7_75t_L g1770 ( .A(n_1771), .Y(n_1770) );
OAI211xp5_ASAP7_75t_L g1822 ( .A1(n_1772), .A2(n_1795), .B(n_1823), .C(n_1824), .Y(n_1822) );
INVx1_ASAP7_75t_L g1772 ( .A(n_1773), .Y(n_1772) );
OR2x2_ASAP7_75t_L g1773 ( .A(n_1774), .B(n_1776), .Y(n_1773) );
NAND2xp5_ASAP7_75t_L g1817 ( .A(n_1774), .B(n_1818), .Y(n_1817) );
AND2x2_ASAP7_75t_L g1835 ( .A(n_1774), .B(n_1836), .Y(n_1835) );
NOR2x1_ASAP7_75t_L g1868 ( .A(n_1774), .B(n_1825), .Y(n_1868) );
INVx2_ASAP7_75t_L g1774 ( .A(n_1775), .Y(n_1774) );
NAND2xp5_ASAP7_75t_L g1785 ( .A(n_1775), .B(n_1786), .Y(n_1785) );
AND2x2_ASAP7_75t_L g1878 ( .A(n_1775), .B(n_1782), .Y(n_1878) );
INVx2_ASAP7_75t_L g1797 ( .A(n_1776), .Y(n_1797) );
AND2x2_ASAP7_75t_L g1854 ( .A(n_1778), .B(n_1855), .Y(n_1854) );
INVx1_ASAP7_75t_L g1778 ( .A(n_1779), .Y(n_1778) );
NOR2xp33_ASAP7_75t_L g1890 ( .A(n_1779), .B(n_1855), .Y(n_1890) );
INVx1_ASAP7_75t_L g1815 ( .A(n_1780), .Y(n_1815) );
NAND2xp5_ASAP7_75t_L g1781 ( .A(n_1782), .B(n_1784), .Y(n_1781) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1783), .Y(n_1782) );
INVx1_ASAP7_75t_L g1784 ( .A(n_1785), .Y(n_1784) );
INVx1_ASAP7_75t_L g1786 ( .A(n_1787), .Y(n_1786) );
INVx1_ASAP7_75t_L g1801 ( .A(n_1787), .Y(n_1801) );
OAI21xp33_ASAP7_75t_L g1888 ( .A1(n_1787), .A2(n_1814), .B(n_1889), .Y(n_1888) );
OAI221xp5_ASAP7_75t_L g1788 ( .A1(n_1789), .A2(n_1793), .B1(n_1794), .B2(n_1796), .C(n_1798), .Y(n_1788) );
NAND2xp5_ASAP7_75t_L g1789 ( .A(n_1790), .B(n_1791), .Y(n_1789) );
INVx1_ASAP7_75t_L g1791 ( .A(n_1792), .Y(n_1791) );
INVx1_ASAP7_75t_SL g1804 ( .A(n_1795), .Y(n_1804) );
NOR3xp33_ASAP7_75t_L g1880 ( .A(n_1795), .B(n_1809), .C(n_1859), .Y(n_1880) );
INVxp67_ASAP7_75t_L g1798 ( .A(n_1799), .Y(n_1798) );
NOR2xp33_ASAP7_75t_L g1831 ( .A(n_1801), .B(n_1832), .Y(n_1831) );
OAI211xp5_ASAP7_75t_SL g1802 ( .A1(n_1803), .A2(n_1805), .B(n_1807), .C(n_1822), .Y(n_1802) );
OAI311xp33_ASAP7_75t_L g1840 ( .A1(n_1803), .A2(n_1841), .A3(n_1842), .B1(n_1850), .C1(n_1856), .Y(n_1840) );
INVx1_ASAP7_75t_L g1845 ( .A(n_1806), .Y(n_1845) );
OR2x2_ASAP7_75t_L g1814 ( .A(n_1809), .B(n_1815), .Y(n_1814) );
INVx1_ASAP7_75t_L g1810 ( .A(n_1811), .Y(n_1810) );
INVx1_ASAP7_75t_L g1813 ( .A(n_1814), .Y(n_1813) );
NAND2xp33_ASAP7_75t_L g1816 ( .A(n_1817), .B(n_1819), .Y(n_1816) );
INVx1_ASAP7_75t_L g1819 ( .A(n_1820), .Y(n_1819) );
INVx1_ASAP7_75t_L g1824 ( .A(n_1825), .Y(n_1824) );
INVx1_ASAP7_75t_L g1827 ( .A(n_1828), .Y(n_1827) );
INVx1_ASAP7_75t_L g1830 ( .A(n_1831), .Y(n_1830) );
INVx1_ASAP7_75t_L g1864 ( .A(n_1832), .Y(n_1864) );
INVx1_ASAP7_75t_L g1841 ( .A(n_1834), .Y(n_1841) );
INVxp67_ASAP7_75t_L g1884 ( .A(n_1835), .Y(n_1884) );
OAI21xp33_ASAP7_75t_L g1842 ( .A1(n_1843), .A2(n_1844), .B(n_1848), .Y(n_1842) );
AND2x2_ASAP7_75t_L g1844 ( .A(n_1845), .B(n_1846), .Y(n_1844) );
INVx1_ASAP7_75t_L g1846 ( .A(n_1847), .Y(n_1846) );
INVx1_ASAP7_75t_L g1851 ( .A(n_1852), .Y(n_1851) );
A2O1A1Ixp33_ASAP7_75t_L g1883 ( .A1(n_1853), .A2(n_1884), .B(n_1885), .C(n_1887), .Y(n_1883) );
INVx1_ASAP7_75t_L g1853 ( .A(n_1854), .Y(n_1853) );
INVx1_ASAP7_75t_L g1858 ( .A(n_1859), .Y(n_1858) );
INVx1_ASAP7_75t_L g1860 ( .A(n_1861), .Y(n_1860) );
NAND2xp5_ASAP7_75t_L g1861 ( .A(n_1862), .B(n_1863), .Y(n_1861) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1866), .Y(n_1871) );
NAND2xp5_ASAP7_75t_L g1869 ( .A(n_1870), .B(n_1871), .Y(n_1869) );
AOI21xp5_ASAP7_75t_L g1872 ( .A1(n_1873), .A2(n_1881), .B(n_1883), .Y(n_1872) );
CKINVDCx14_ASAP7_75t_R g1881 ( .A(n_1882), .Y(n_1881) );
INVx1_ASAP7_75t_L g1885 ( .A(n_1886), .Y(n_1885) );
INVxp33_ASAP7_75t_L g1889 ( .A(n_1890), .Y(n_1889) );
INVx1_ASAP7_75t_L g1895 ( .A(n_1896), .Y(n_1895) );
HB1xp67_ASAP7_75t_L g1899 ( .A(n_1900), .Y(n_1899) );
INVx1_ASAP7_75t_L g1900 ( .A(n_1901), .Y(n_1900) );
HB1xp67_ASAP7_75t_L g1959 ( .A(n_1903), .Y(n_1959) );
NAND3xp33_ASAP7_75t_L g1903 ( .A(n_1904), .B(n_1929), .C(n_1931), .Y(n_1903) );
INVx1_ASAP7_75t_L g1921 ( .A(n_1922), .Y(n_1921) );
INVx1_ASAP7_75t_L g1926 ( .A(n_1927), .Y(n_1926) );
NOR2xp33_ASAP7_75t_SL g1931 ( .A(n_1932), .B(n_1944), .Y(n_1931) );
INVx1_ASAP7_75t_L g1942 ( .A(n_1943), .Y(n_1942) );
NAND2xp5_ASAP7_75t_L g1944 ( .A(n_1945), .B(n_1946), .Y(n_1944) );
CKINVDCx14_ASAP7_75t_R g1947 ( .A(n_1948), .Y(n_1947) );
BUFx2_ASAP7_75t_L g1948 ( .A(n_1949), .Y(n_1948) );
INVx1_ASAP7_75t_L g1949 ( .A(n_1950), .Y(n_1949) );
INVx1_ASAP7_75t_L g1950 ( .A(n_1951), .Y(n_1950) );
HB1xp67_ASAP7_75t_SL g1953 ( .A(n_1954), .Y(n_1953) );
A2O1A1Ixp33_ASAP7_75t_L g1961 ( .A1(n_1955), .A2(n_1962), .B(n_1964), .C(n_1965), .Y(n_1961) );
INVxp33_ASAP7_75t_SL g1956 ( .A(n_1957), .Y(n_1956) );
INVx1_ASAP7_75t_L g1958 ( .A(n_1959), .Y(n_1958) );
HB1xp67_ASAP7_75t_L g1960 ( .A(n_1961), .Y(n_1960) );
INVx1_ASAP7_75t_L g1962 ( .A(n_1963), .Y(n_1962) );
endmodule