module fake_jpeg_31002_n_187 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_187);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_49),
.Y(n_57)
);

BUFx6f_ASAP7_75t_SL g58 ( 
.A(n_19),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_33),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_9),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_7),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g85 ( 
.A(n_75),
.B(n_51),
.Y(n_85)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_1),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_72),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_90),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_82),
.A2(n_51),
.B1(n_73),
.B2(n_72),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_96),
.B1(n_76),
.B2(n_67),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_55),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_66),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_74),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_83),
.C(n_80),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_73),
.B1(n_72),
.B2(n_66),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_100),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_88),
.B(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_99),
.B(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_89),
.B(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_55),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_106),
.Y(n_127)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_81),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_63),
.Y(n_132)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_113),
.Y(n_116)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_70),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_95),
.C(n_85),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_117),
.C(n_132),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_106),
.A2(n_108),
.B1(n_112),
.B2(n_92),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_123),
.B1(n_6),
.B2(n_8),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_90),
.B(n_82),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_SL g155 ( 
.A1(n_118),
.A2(n_31),
.B(n_44),
.C(n_43),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_54),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_122),
.B(n_131),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_92),
.B1(n_60),
.B2(n_65),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_130),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_5),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_104),
.B(n_61),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_56),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_105),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_25),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_59),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_136),
.B(n_10),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_146),
.Y(n_160)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_147),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_148),
.C(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_143),
.B(n_146),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_57),
.B(n_52),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_144),
.B(n_149),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_156),
.B1(n_142),
.B2(n_14),
.Y(n_166)
);

NOR2x1p5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_28),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_29),
.C(n_46),
.Y(n_148)
);

AO22x1_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_126),
.B1(n_128),
.B2(n_116),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

BUFx24_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_151),
.B(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_11),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_155),
.B(n_35),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_161),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_160),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_133),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_23),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_163),
.Y(n_173)
);

OAI321xp33_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_155),
.A3(n_137),
.B1(n_12),
.B2(n_14),
.C(n_17),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_164),
.A2(n_155),
.B(n_154),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_170),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_164),
.A2(n_15),
.A3(n_16),
.B1(n_18),
.B2(n_21),
.C1(n_36),
.C2(n_37),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_168),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_176),
.A2(n_173),
.B1(n_172),
.B2(n_165),
.Y(n_179)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

OAI21x1_ASAP7_75t_L g180 ( 
.A1(n_178),
.A2(n_179),
.B(n_170),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_175),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_165),
.C(n_169),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_167),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_157),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_162),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_157),
.C(n_39),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_186),
.B(n_47),
.Y(n_187)
);


endmodule