module fake_jpeg_31448_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_57),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_1),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_1),
.B(n_2),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_51),
.B1(n_55),
.B2(n_58),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_29),
.B(n_30),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_51),
.Y(n_90)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_53),
.Y(n_92)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_81),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_61),
.B(n_46),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_79),
.A2(n_55),
.B1(n_47),
.B2(n_53),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_58),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_12),
.B(n_42),
.Y(n_109)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_91),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_56),
.C(n_45),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_77),
.C(n_5),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_52),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_4),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_44),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_2),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_11),
.Y(n_108)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_89),
.A2(n_77),
.B1(n_71),
.B2(n_6),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_102),
.B(n_107),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_108),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_12),
.B1(n_94),
.B2(n_18),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_106),
.B1(n_111),
.B2(n_94),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_92),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_109),
.B(n_110),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_85),
.B(n_26),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_41),
.B1(n_13),
.B2(n_15),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_83),
.Y(n_115)
);

BUFx24_ASAP7_75t_SL g116 ( 
.A(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_119),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_117),
.B(n_118),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_106),
.A2(n_17),
.B1(n_20),
.B2(n_23),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_121),
.B(n_105),
.Y(n_125)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_110),
.B(n_107),
.C(n_102),
.D(n_111),
.Y(n_124)
);

A2O1A1O1Ixp25_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_118),
.B(n_100),
.C(n_117),
.D(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_114),
.C(n_112),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_128),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_126),
.C(n_129),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_121),
.Y(n_132)
);

OAI221xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_122),
.B1(n_27),
.B2(n_32),
.C(n_35),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_25),
.B1(n_36),
.B2(n_37),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_38),
.Y(n_135)
);


endmodule