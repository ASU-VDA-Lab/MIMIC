module fake_jpeg_8060_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_31),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_29),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_26),
.B(n_24),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_54),
.Y(n_70)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_34),
.A2(n_19),
.B1(n_30),
.B2(n_29),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_62),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_34),
.A2(n_19),
.B1(n_28),
.B2(n_31),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_63),
.B(n_24),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_18),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_15),
.B1(n_21),
.B2(n_20),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_78),
.B1(n_52),
.B2(n_56),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_39),
.B1(n_38),
.B2(n_21),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_81),
.C(n_72),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_56),
.B1(n_46),
.B2(n_17),
.Y(n_99)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_76),
.Y(n_84)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_74),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_25),
.B1(n_33),
.B2(n_36),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_75),
.A2(n_46),
.B1(n_53),
.B2(n_49),
.Y(n_103)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_47),
.B1(n_52),
.B2(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_83),
.B(n_89),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_100),
.B1(n_103),
.B2(n_76),
.Y(n_107)
);

OR2x2_ASAP7_75t_SL g86 ( 
.A(n_82),
.B(n_17),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_88),
.B(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_61),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_1),
.C(n_2),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_0),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_45),
.B(n_73),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_95),
.B(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_42),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_53),
.B1(n_49),
.B2(n_71),
.Y(n_113)
);

OAI22x1_ASAP7_75t_SL g100 ( 
.A1(n_64),
.A2(n_40),
.B1(n_41),
.B2(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_69),
.B(n_9),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_66),
.B(n_36),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_73),
.Y(n_112)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_105),
.B(n_123),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_80),
.C(n_46),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_122),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_99),
.B1(n_91),
.B2(n_87),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_100),
.B1(n_96),
.B2(n_85),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_113),
.B1(n_84),
.B2(n_87),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_97),
.B(n_95),
.Y(n_139)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_114),
.B(n_116),
.Y(n_138)
);

AO22x1_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_44),
.B1(n_50),
.B2(n_71),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_125),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_53),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_44),
.B1(n_71),
.B2(n_50),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_50),
.B1(n_55),
.B2(n_74),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_0),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_124),
.B(n_25),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_41),
.C(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_86),
.A2(n_18),
.B(n_17),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_93),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_126),
.B(n_141),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_143),
.B1(n_113),
.B2(n_123),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_131),
.B(n_139),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_108),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_133),
.Y(n_163)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_108),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_94),
.Y(n_136)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_18),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_25),
.B(n_2),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_142),
.A2(n_145),
.B(n_125),
.Y(n_161)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_144),
.B(n_115),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_1),
.B(n_2),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_147),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_135),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_150),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_107),
.B1(n_132),
.B2(n_119),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_153),
.A2(n_157),
.B(n_159),
.Y(n_166)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_156),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_109),
.B(n_105),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_129),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_161),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_106),
.B(n_117),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_162),
.A2(n_144),
.B(n_121),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_164),
.A2(n_178),
.B1(n_162),
.B2(n_149),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_154),
.B(n_126),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_177),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_153),
.A2(n_110),
.B1(n_133),
.B2(n_134),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_170),
.A2(n_171),
.B(n_151),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_121),
.A3(n_137),
.B1(n_142),
.B2(n_136),
.C1(n_145),
.C2(n_124),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_157),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_137),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_175),
.C(n_161),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_122),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_147),
.A2(n_121),
.B1(n_115),
.B2(n_116),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_186),
.B(n_45),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_174),
.B(n_158),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_180),
.B(n_167),
.Y(n_195)
);

MAJx2_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_159),
.C(n_160),
.Y(n_181)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_3),
.C(n_5),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_164),
.B(n_168),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_171),
.A2(n_155),
.B1(n_151),
.B2(n_149),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_185),
.A2(n_190),
.B1(n_3),
.B2(n_5),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_188),
.C(n_189),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_163),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_163),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_176),
.A2(n_55),
.B1(n_45),
.B2(n_4),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_196),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_195),
.Y(n_201)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_179),
.A2(n_166),
.B(n_170),
.C(n_178),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_194),
.B(n_200),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_183),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_187),
.B(n_11),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_198),
.A2(n_190),
.B1(n_181),
.B2(n_189),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_182),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_8),
.C(n_10),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_200),
.Y(n_210)
);

NOR2xp67_ASAP7_75t_R g205 ( 
.A(n_199),
.B(n_182),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_10),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_207),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_201),
.A2(n_193),
.B(n_194),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_212),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_211),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_193),
.Y(n_211)
);

XOR2x2_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_207),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_213),
.A2(n_206),
.B(n_13),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

AOI21x1_ASAP7_75t_L g217 ( 
.A1(n_209),
.A2(n_11),
.B(n_13),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_11),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_218),
.A2(n_14),
.B(n_215),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_210),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_14),
.C(n_219),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_222),
.C(n_220),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_14),
.Y(n_224)
);


endmodule