module fake_jpeg_24889_n_270 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx11_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

CKINVDCx9p33_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_42),
.B(n_26),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_45),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_23),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_21),
.Y(n_54)
);

OR2x2_ASAP7_75t_SL g101 ( 
.A(n_54),
.B(n_64),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_33),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_62),
.Y(n_97)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_23),
.B1(n_32),
.B2(n_19),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_59),
.B1(n_18),
.B2(n_34),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_23),
.B1(n_32),
.B2(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_27),
.Y(n_62)
);

HAxp5_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_18),
.CON(n_64),
.SN(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_24),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_65),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_70),
.Y(n_104)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_68),
.B(n_78),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_16),
.B1(n_19),
.B2(n_27),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_85),
.B1(n_91),
.B2(n_35),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_36),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_30),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_74),
.Y(n_110)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_76),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_42),
.A2(n_28),
.B1(n_16),
.B2(n_26),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_77),
.A2(n_18),
.B1(n_17),
.B2(n_2),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_35),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_15),
.Y(n_95)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_71),
.B1(n_51),
.B2(n_89),
.Y(n_92)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_43),
.A2(n_20),
.B1(n_29),
.B2(n_22),
.Y(n_85)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_25),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_90),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_43),
.A2(n_20),
.B1(n_29),
.B2(n_22),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_93),
.A2(n_71),
.B1(n_51),
.B2(n_86),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_95),
.B(n_13),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_96),
.A2(n_114),
.B1(n_118),
.B2(n_57),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_54),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_116),
.Y(n_124)
);

OA22x2_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_62),
.B1(n_59),
.B2(n_77),
.Y(n_105)
);

AND2x4_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_81),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_34),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_109),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_50),
.B(n_34),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_63),
.B(n_17),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_87),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_56),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_80),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_122),
.A2(n_1),
.B1(n_5),
.B2(n_7),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_121),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_127),
.B(n_134),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_128),
.A2(n_131),
.B1(n_135),
.B2(n_154),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_83),
.B(n_82),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_86),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_132),
.B(n_139),
.Y(n_166)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_74),
.B(n_73),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_143),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_98),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_141),
.Y(n_172)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_138),
.B(n_140),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_73),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_104),
.B(n_60),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_114),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_63),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g174 ( 
.A(n_144),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_113),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_148),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_120),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_149),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_100),
.B(n_57),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_152),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_100),
.B(n_108),
.Y(n_153)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_168),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_101),
.B1(n_97),
.B2(n_96),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_163),
.B1(n_165),
.B2(n_167),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_128),
.A2(n_101),
.B1(n_97),
.B2(n_94),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_159),
.A2(n_157),
.B1(n_165),
.B2(n_163),
.Y(n_207)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_109),
.B(n_97),
.C(n_99),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_94),
.B1(n_120),
.B2(n_102),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_102),
.B1(n_107),
.B2(n_111),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_130),
.A2(n_122),
.B1(n_87),
.B2(n_66),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_126),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_111),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_179),
.Y(n_204)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_108),
.B1(n_116),
.B2(n_95),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_137),
.B1(n_148),
.B2(n_149),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_63),
.Y(n_183)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_150),
.B(n_156),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_186),
.A2(n_203),
.B(n_189),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_184),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_196),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_138),
.C(n_152),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_175),
.C(n_161),
.Y(n_211)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_194),
.Y(n_221)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_178),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_182),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_198),
.A2(n_174),
.B1(n_129),
.B2(n_125),
.Y(n_224)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_145),
.C(n_146),
.Y(n_199)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_183),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_171),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_154),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_177),
.B(n_141),
.Y(n_206)
);

BUFx24_ASAP7_75t_SL g219 ( 
.A(n_206),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_170),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_164),
.B(n_147),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_208),
.A2(n_166),
.B(n_179),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_209),
.B(n_207),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_185),
.A2(n_176),
.B1(n_173),
.B2(n_167),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_220),
.C(n_223),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_225),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_185),
.A2(n_167),
.B1(n_181),
.B2(n_162),
.Y(n_214)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_164),
.C(n_158),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_226),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_158),
.C(n_167),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_225),
.B1(n_190),
.B2(n_193),
.Y(n_237)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

AOI321xp33_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_202),
.A3(n_199),
.B1(n_201),
.B2(n_188),
.C(n_205),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_212),
.B(n_217),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_191),
.C(n_202),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_230),
.C(n_233),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_188),
.C(n_186),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_238),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_195),
.C(n_194),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_221),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_234),
.Y(n_247)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_237),
.B(n_239),
.Y(n_245)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_210),
.Y(n_242)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_214),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_231),
.Y(n_254)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_229),
.B(n_203),
.CI(n_219),
.CON(n_248),
.SN(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_197),
.C(n_187),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_241),
.C(n_227),
.Y(n_252)
);

OAI21x1_ASAP7_75t_SL g250 ( 
.A1(n_240),
.A2(n_226),
.B(n_204),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_250),
.A2(n_232),
.B1(n_235),
.B2(n_228),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_233),
.B(n_14),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_14),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_256),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_245),
.Y(n_256)
);

NOR2x1_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_244),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_R g263 ( 
.A(n_259),
.B(n_261),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_246),
.Y(n_260)
);

OAI21x1_ASAP7_75t_L g261 ( 
.A1(n_253),
.A2(n_243),
.B(n_242),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_174),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_252),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_263),
.A2(n_262),
.B(n_260),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_266),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_264),
.A2(n_248),
.B1(n_174),
.B2(n_129),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_267),
.A2(n_144),
.B(n_9),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_7),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_7),
.Y(n_270)
);


endmodule