module fake_jpeg_23769_n_101 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_25),
.A2(n_17),
.B1(n_24),
.B2(n_19),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_2),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_15),
.B(n_19),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_34),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_3),
.Y(n_32)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_12),
.Y(n_46)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_24),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_14),
.B1(n_34),
.B2(n_22),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_30),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_47),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_15),
.C(n_12),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_13),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_60),
.B1(n_6),
.B2(n_7),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_36),
.B1(n_41),
.B2(n_43),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_67)
);

BUFx24_ASAP7_75t_SL g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_56),
.B(n_46),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_45),
.Y(n_73)
);

OA21x2_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_34),
.B(n_21),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_14),
.B1(n_21),
.B2(n_22),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_22),
.B1(n_5),
.B2(n_4),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_73),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_39),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_69),
.C(n_74),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_35),
.B1(n_39),
.B2(n_42),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_51),
.B1(n_60),
.B2(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_45),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_8),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_72),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_83),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_50),
.C(n_54),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_50),
.C(n_67),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_88),
.C(n_89),
.Y(n_90)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_86),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_74),
.B(n_68),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_67),
.C(n_63),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_73),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_84),
.B1(n_81),
.B2(n_83),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_92),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_89),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_60),
.C(n_59),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_82),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_96),
.C(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_92),
.Y(n_98)
);

AOI321xp33_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_98),
.A3(n_91),
.B1(n_95),
.B2(n_59),
.C(n_10),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_80),
.Y(n_101)
);


endmodule