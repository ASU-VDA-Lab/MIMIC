module fake_netlist_6_1996_n_125 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_2, n_5, n_19, n_29, n_25, n_125);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;
input n_29;
input n_25;

output n_125;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_68;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_99;
wire n_85;
wire n_78;
wire n_84;
wire n_100;
wire n_121;
wire n_47;
wire n_62;
wire n_75;
wire n_109;
wire n_122;
wire n_45;
wire n_34;
wire n_70;
wire n_120;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_94;
wire n_108;
wire n_97;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_35;
wire n_115;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVxp67_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_16),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

INVxp67_ASAP7_75t_SL g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_2),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVxp67_ASAP7_75t_SL g50 ( 
.A(n_17),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_0),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_30),
.B(n_0),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_53),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_51),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_59),
.B(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_45),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_45),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_65),
.B(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_51),
.C(n_38),
.Y(n_84)
);

AO21x2_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_73),
.B(n_76),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_62),
.B1(n_55),
.B2(n_60),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_37),
.B(n_40),
.Y(n_87)
);

AO21x2_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_54),
.B(n_33),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_55),
.B1(n_62),
.B2(n_6),
.Y(n_89)
);

AND2x4_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_62),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_R g91 ( 
.A(n_81),
.B(n_2),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_62),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_55),
.Y(n_95)
);

AND2x4_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_24),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_55),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

AND2x4_ASAP7_75t_SL g99 ( 
.A(n_96),
.B(n_93),
.Y(n_99)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_93),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_82),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_82),
.Y(n_102)
);

AO221x2_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_87),
.B1(n_91),
.B2(n_80),
.C(n_84),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_98),
.A2(n_91),
.B1(n_96),
.B2(n_80),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_99),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_88),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_101),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

AOI211xp5_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_109),
.B(n_90),
.C(n_88),
.Y(n_113)
);

NOR3xp33_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_92),
.C(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_111),
.Y(n_116)
);

NAND2xp33_ASAP7_75t_SL g117 ( 
.A(n_113),
.B(n_88),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_5),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_114),
.B1(n_89),
.B2(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_85),
.B1(n_90),
.B2(n_95),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_85),
.B1(n_86),
.B2(n_100),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_85),
.B1(n_6),
.B2(n_5),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_R g124 ( 
.A1(n_123),
.A2(n_85),
.B1(n_22),
.B2(n_25),
.Y(n_124)
);

AOI221xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_121),
.B1(n_122),
.B2(n_27),
.C(n_8),
.Y(n_125)
);


endmodule