module fake_jpeg_16895_n_183 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_183);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_SL g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_6),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_32),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_34),
.Y(n_38)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_32),
.A2(n_22),
.B1(n_19),
.B2(n_24),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_46),
.B(n_18),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_13),
.B(n_35),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_28),
.B(n_29),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_0),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_22),
.B1(n_24),
.B2(n_12),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_58),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_38),
.B1(n_44),
.B2(n_41),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_48),
.B1(n_65),
.B2(n_53),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_22),
.B1(n_16),
.B2(n_12),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_59),
.B(n_70),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

AO22x1_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_61),
.B1(n_37),
.B2(n_31),
.Y(n_78)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_16),
.B1(n_18),
.B2(n_12),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_63),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_46),
.A2(n_16),
.B1(n_24),
.B2(n_18),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_35),
.C(n_30),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_27),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_33),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_31),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_39),
.B(n_23),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

OAI32xp33_ASAP7_75t_L g72 ( 
.A1(n_42),
.A2(n_15),
.A3(n_25),
.B1(n_14),
.B2(n_21),
.Y(n_72)
);

OAI32xp33_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_52),
.A3(n_15),
.B1(n_68),
.B2(n_14),
.Y(n_90)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_37),
.B1(n_31),
.B2(n_40),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_78),
.B1(n_80),
.B2(n_56),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_1),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_1),
.B(n_57),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_29),
.B1(n_27),
.B2(n_15),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_30),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_90),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_93),
.C(n_64),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_21),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_21),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_94),
.A2(n_72),
.B1(n_54),
.B2(n_73),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_17),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_54),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_109),
.B1(n_113),
.B2(n_114),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_71),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_102),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_93),
.C(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_101),
.B(n_112),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_17),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_105),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_17),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_106),
.A2(n_108),
.B(n_117),
.Y(n_128)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_55),
.B1(n_58),
.B2(n_57),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_110),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_57),
.B1(n_62),
.B2(n_30),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_80),
.B1(n_79),
.B2(n_88),
.Y(n_124)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_62),
.B1(n_17),
.B2(n_4),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_83),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_6),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_81),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_75),
.Y(n_134)
);

AND2x4_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_7),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_131),
.C(n_121),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_88),
.B(n_82),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_121),
.A2(n_124),
.B(n_104),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_133),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_78),
.B1(n_95),
.B2(n_90),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_117),
.B1(n_79),
.B2(n_115),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_76),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_76),
.Y(n_132)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g133 ( 
.A(n_99),
.B(n_91),
.CI(n_75),
.CON(n_133),
.SN(n_133)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_134),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_111),
.B(n_117),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_136),
.A2(n_141),
.B1(n_146),
.B2(n_124),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_143),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_99),
.B(n_117),
.C(n_95),
.D(n_101),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_138),
.B(n_145),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_113),
.C(n_112),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_128),
.A2(n_104),
.B(n_110),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_144),
.A2(n_123),
.B1(n_134),
.B2(n_129),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_114),
.B(n_8),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_150),
.A2(n_152),
.B1(n_136),
.B2(n_141),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_129),
.B1(n_140),
.B2(n_142),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_153),
.A2(n_155),
.B1(n_120),
.B2(n_122),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_137),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_164),
.C(n_8),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_143),
.C(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_163),
.C(n_127),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_138),
.B(n_127),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_145),
.C(n_133),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_130),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_163),
.A2(n_148),
.B(n_152),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_168),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_160),
.B(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

OAI221xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_171),
.B1(n_164),
.B2(n_161),
.C(n_158),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_159),
.B(n_7),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

OAI221xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_9),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_179),
.C(n_10),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_170),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_177),
.A2(n_172),
.B(n_176),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_181),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_178),
.B(n_11),
.Y(n_183)
);


endmodule