module fake_jpeg_24106_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_49),
.Y(n_70)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_28),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_21),
.B(n_0),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_24),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_31),
.B1(n_34),
.B2(n_18),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_62),
.B(n_63),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_31),
.B1(n_36),
.B2(n_18),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_56),
.A2(n_68),
.B1(n_74),
.B2(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_71),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_31),
.B1(n_34),
.B2(n_18),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_31),
.B1(n_34),
.B2(n_23),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_72),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_66),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_36),
.B1(n_27),
.B2(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_27),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_21),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_81),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_42),
.A2(n_36),
.B1(n_25),
.B2(n_24),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_35),
.Y(n_77)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_39),
.A2(n_24),
.B1(n_17),
.B2(n_19),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_78),
.A2(n_19),
.B1(n_17),
.B2(n_29),
.Y(n_121)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_26),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_84),
.Y(n_115)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_26),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_17),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_50),
.A2(n_29),
.B1(n_21),
.B2(n_22),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_88),
.B(n_100),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_57),
.B(n_50),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_91),
.B(n_99),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_60),
.B(n_35),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_65),
.B(n_48),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_41),
.C(n_47),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_79),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_103),
.A2(n_111),
.B1(n_114),
.B2(n_116),
.Y(n_158)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_60),
.B(n_32),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_32),
.B1(n_26),
.B2(n_22),
.Y(n_127)
);

OR2x2_ASAP7_75t_SL g109 ( 
.A(n_65),
.B(n_16),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_33),
.B(n_8),
.C(n_9),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_117),
.Y(n_131)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_70),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_70),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_47),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

NAND2x1_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_48),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_120),
.A2(n_121),
.B(n_38),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_85),
.B(n_19),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_86),
.B(n_29),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_64),
.B1(n_67),
.B2(n_72),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_124),
.A2(n_128),
.B1(n_151),
.B2(n_153),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_126),
.B(n_127),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_64),
.B1(n_67),
.B2(n_55),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_22),
.B1(n_76),
.B2(n_55),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_144),
.B1(n_92),
.B2(n_122),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_120),
.A2(n_82),
.B(n_2),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_136),
.B(n_140),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_133),
.C(n_134),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_71),
.C(n_83),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_47),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_41),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_96),
.C(n_119),
.Y(n_177)
);

NAND2x1_ASAP7_75t_SL g136 ( 
.A(n_87),
.B(n_76),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_101),
.A2(n_80),
.B1(n_61),
.B2(n_59),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_142),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_87),
.B(n_61),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_145),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_93),
.A2(n_84),
.B1(n_33),
.B2(n_66),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_89),
.B(n_33),
.Y(n_145)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_95),
.A2(n_66),
.B1(n_37),
.B2(n_38),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_152),
.B(n_156),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_95),
.A2(n_117),
.B1(n_111),
.B2(n_89),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_102),
.A2(n_37),
.B1(n_38),
.B2(n_3),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_155),
.A2(n_106),
.B1(n_38),
.B2(n_37),
.Y(n_194)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_105),
.B1(n_92),
.B2(n_97),
.Y(n_181)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_162),
.B(n_168),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_138),
.A2(n_104),
.B1(n_118),
.B2(n_116),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_163),
.A2(n_166),
.B1(n_171),
.B2(n_172),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_102),
.B(n_110),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_175),
.B(n_179),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_149),
.A2(n_114),
.B1(n_105),
.B2(n_103),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_153),
.B(n_135),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_173),
.Y(n_210)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_186),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_128),
.B1(n_132),
.B2(n_133),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_131),
.A2(n_136),
.B1(n_134),
.B2(n_143),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_173),
.A2(n_176),
.B1(n_181),
.B2(n_147),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_131),
.A2(n_91),
.B(n_109),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_124),
.B1(n_145),
.B2(n_130),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_182),
.C(n_112),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_141),
.B(n_96),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_178),
.B(n_188),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_126),
.A2(n_107),
.B(n_99),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_90),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_192),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_90),
.C(n_108),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_1),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_183),
.A2(n_2),
.B(n_3),
.Y(n_215)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_125),
.B(n_94),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_146),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_190),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_148),
.B(n_108),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_191),
.Y(n_214)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_159),
.B1(n_142),
.B2(n_112),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_205),
.B1(n_217),
.B2(n_218),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_38),
.B1(n_94),
.B2(n_98),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_198),
.B(n_211),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_37),
.Y(n_201)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_204),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_161),
.A2(n_98),
.B1(n_37),
.B2(n_3),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_1),
.C(n_2),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_208),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_1),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_160),
.A2(n_9),
.B(n_15),
.C(n_14),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_209),
.B(n_179),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_215),
.Y(n_239)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_171),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_212),
.B(n_216),
.Y(n_245)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_169),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_172),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_219),
.B(n_223),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_160),
.A2(n_5),
.B(n_6),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_183),
.B(n_165),
.Y(n_235)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_170),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_224),
.A2(n_170),
.B1(n_185),
.B2(n_183),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_203),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_225),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_213),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_226),
.B(n_233),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_229),
.Y(n_255)
);

BUFx4f_ASAP7_75t_SL g230 ( 
.A(n_223),
.Y(n_230)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_247),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_203),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_215),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_176),
.B(n_164),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_248),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_161),
.B1(n_162),
.B2(n_177),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_238),
.A2(n_244),
.B1(n_205),
.B2(n_208),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_221),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_175),
.Y(n_241)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_212),
.A2(n_216),
.B1(n_195),
.B2(n_218),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_200),
.Y(n_247)
);

NAND2xp33_ASAP7_75t_SL g248 ( 
.A(n_199),
.B(n_167),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_247),
.B1(n_242),
.B2(n_241),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_249),
.A2(n_256),
.B1(n_263),
.B2(n_229),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_202),
.C(n_201),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_252),
.C(n_254),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_211),
.C(n_199),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_234),
.B1(n_232),
.B2(n_227),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_210),
.C(n_206),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_245),
.A2(n_217),
.B1(n_224),
.B2(n_219),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_235),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_196),
.C(n_192),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_228),
.C(n_226),
.Y(n_282)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_230),
.Y(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_268),
.Y(n_269)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_250),
.A2(n_225),
.B(n_233),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_286),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_227),
.B1(n_236),
.B2(n_244),
.Y(n_273)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_283),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_281),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_236),
.B1(n_230),
.B2(n_238),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_276),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_214),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_280),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_193),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_248),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_284),
.C(n_285),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_174),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_228),
.C(n_230),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_186),
.C(n_204),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_214),
.C(n_198),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_269),
.A2(n_274),
.B1(n_268),
.B2(n_265),
.Y(n_288)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

INVx13_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_257),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_249),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_299),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_266),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_284),
.C(n_282),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_302),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_243),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_285),
.C(n_286),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_305),
.Y(n_316)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_288),
.B(n_276),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_306),
.A2(n_287),
.B1(n_294),
.B2(n_209),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_259),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_309),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_243),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_295),
.B1(n_187),
.B2(n_221),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_259),
.C(n_263),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_293),
.B1(n_291),
.B2(n_296),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_311),
.B1(n_315),
.B2(n_317),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_258),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_298),
.B1(n_299),
.B2(n_281),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_305),
.A2(n_292),
.B1(n_266),
.B2(n_275),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_319),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_313),
.A2(n_304),
.B(n_187),
.Y(n_319)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_314),
.A2(n_174),
.B(n_9),
.Y(n_320)
);

AO21x1_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_10),
.B(n_11),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_6),
.C(n_10),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_13),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_324),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_325),
.A2(n_321),
.B(n_316),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_314),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_322),
.C(n_323),
.Y(n_329)
);

AOI21x1_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_326),
.B(n_310),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_317),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_16),
.Y(n_332)
);


endmodule