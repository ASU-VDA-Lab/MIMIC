module fake_jpeg_17293_n_114 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_26),
.B(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_28),
.B(n_30),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_25),
.B(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_29),
.B(n_32),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_1),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_3),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_4),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_10),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_19),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_33),
.A2(n_22),
.B1(n_14),
.B2(n_12),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_36),
.B1(n_7),
.B2(n_8),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_50),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_31),
.A2(n_17),
.B1(n_14),
.B2(n_22),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_53),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_26),
.B(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_4),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_57),
.Y(n_79)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_45),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_64),
.B1(n_67),
.B2(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_61),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_36),
.C(n_7),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_65),
.C(n_69),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_6),
.B(n_8),
.Y(n_65)
);

AO21x1_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_40),
.B(n_54),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_69),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_41),
.B(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_78),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_49),
.B(n_55),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_55),
.B(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_82),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_58),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_56),
.C(n_66),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_90),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_72),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_62),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_77),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_60),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_79),
.B1(n_87),
.B2(n_83),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_89),
.C(n_86),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_92),
.C(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_103),
.A2(n_90),
.B1(n_98),
.B2(n_77),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_105),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_94),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

OAI321xp33_ASAP7_75t_L g107 ( 
.A1(n_101),
.A2(n_91),
.A3(n_92),
.B1(n_79),
.B2(n_59),
.C(n_60),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_99),
.B(n_102),
.C(n_70),
.D(n_75),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_76),
.C(n_75),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_111),
.A2(n_109),
.B(n_112),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);


endmodule