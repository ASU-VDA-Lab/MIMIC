module real_jpeg_12525_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_401, n_6, n_402, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_401;
input n_6;
input n_402;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_0),
.Y(n_108)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_3),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_3),
.B(n_95),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_3),
.B(n_32),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_3),
.B(n_29),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_3),
.B(n_53),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_3),
.B(n_40),
.Y(n_293)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_5),
.B(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_5),
.B(n_53),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_5),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_5),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_5),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_5),
.B(n_40),
.Y(n_327)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_6),
.Y(n_97)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_7),
.B(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_7),
.B(n_108),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_7),
.B(n_95),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_7),
.B(n_26),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_7),
.B(n_29),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_8),
.B(n_29),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_8),
.B(n_53),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_8),
.B(n_26),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_8),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_8),
.B(n_40),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_12),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_12),
.B(n_45),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_12),
.B(n_95),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_12),
.B(n_32),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_12),
.B(n_26),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_13),
.B(n_26),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_13),
.B(n_29),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_13),
.B(n_95),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_13),
.B(n_32),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_13),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_13),
.B(n_53),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_13),
.B(n_40),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_13),
.B(n_45),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_14),
.B(n_32),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_14),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_14),
.B(n_108),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_14),
.B(n_29),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_14),
.B(n_40),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_14),
.B(n_45),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_15),
.B(n_53),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_15),
.B(n_40),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_15),
.B(n_26),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_15),
.B(n_108),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_15),
.B(n_95),
.Y(n_208)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_119),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_118),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_79),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_21),
.B(n_79),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_64),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_48),
.C(n_55),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_23),
.B(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_37),
.C(n_41),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.C(n_31),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_25),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_25),
.B(n_57),
.C(n_62),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_25),
.A2(n_31),
.B1(n_63),
.B2(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_25),
.A2(n_63),
.B1(n_109),
.B2(n_110),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_25),
.B(n_109),
.C(n_252),
.Y(n_272)
);

INVx5_ASAP7_75t_SL g148 ( 
.A(n_26),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_28),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_28),
.A2(n_83),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_28),
.B(n_290),
.C(n_293),
.Y(n_338)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_30),
.B(n_38),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_31),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_31),
.B(n_93),
.C(n_98),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_31),
.A2(n_86),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_31),
.B(n_200),
.C(n_202),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_31),
.A2(n_86),
.B1(n_93),
.B2(n_94),
.Y(n_372)
);

CKINVDCx14_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_33),
.B(n_51),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_33),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_33),
.B(n_43),
.Y(n_269)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_38),
.B(n_136),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_44),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_44),
.B(n_179),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_44),
.B(n_137),
.Y(n_329)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_48),
.A2(n_55),
.B1(n_56),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.C(n_52),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_49),
.B(n_52),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_50),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_50),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_53),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_57),
.A2(n_58),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_107),
.C(n_109),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_62),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_61),
.A2(n_62),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_62),
.B(n_98),
.C(n_264),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_78),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_73),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_89),
.C(n_90),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_67),
.A2(n_71),
.B1(n_365),
.B2(n_366),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_68),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_69),
.A2(n_70),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_70),
.B(n_303),
.C(n_305),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_113),
.C(n_114),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_80),
.B(n_394),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_99),
.C(n_103),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_81),
.B(n_388),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_87),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_88),
.C(n_92),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_89),
.B(n_90),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_91),
.B(n_134),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_105),
.C(n_111),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_93),
.A2(n_94),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_93),
.A2(n_94),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_93),
.A2(n_94),
.B1(n_111),
.B2(n_360),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_94),
.B(n_160),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_94),
.B(n_343),
.C(n_345),
.Y(n_361)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_96),
.B(n_179),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_98),
.A2(n_261),
.B1(n_262),
.B2(n_265),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_98),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_98),
.A2(n_265),
.B1(n_371),
.B2(n_372),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_99),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_101),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_105),
.A2(n_106),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_107),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_107),
.B(n_139),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_107),
.A2(n_141),
.B1(n_207),
.B2(n_208),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_107),
.A2(n_109),
.B1(n_110),
.B2(n_141),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_107),
.B(n_208),
.C(n_306),
.Y(n_343)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_111),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_113),
.Y(n_395)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI321xp33_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_382),
.A3(n_391),
.B1(n_396),
.B2(n_397),
.C(n_401),
.Y(n_119)
);

AOI321xp33_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_314),
.A3(n_348),
.B1(n_376),
.B2(n_381),
.C(n_402),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_255),
.C(n_309),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_226),
.B(n_254),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_194),
.B(n_225),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_163),
.B(n_193),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_142),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_126),
.B(n_142),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.C(n_138),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_145),
.B1(n_146),
.B2(n_154),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_127),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_127),
.B(n_190),
.Y(n_189)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_129),
.CI(n_130),
.CON(n_127),
.SN(n_127)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_131),
.A2(n_132),
.B1(n_138),
.B2(n_191),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_133),
.B(n_135),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_136),
.B(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_137),
.B(n_148),
.Y(n_200)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_138),
.Y(n_191)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_155),
.B2(n_162),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_154),
.C(n_162),
.Y(n_195)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_147),
.B(n_150),
.C(n_153),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_156),
.B(n_158),
.C(n_159),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_160),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_160),
.A2(n_161),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_160),
.B(n_277),
.C(n_280),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_187),
.B(n_192),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_176),
.B(n_186),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_171),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_166),
.B(n_171),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_174),
.C(n_175),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_181),
.B(n_185),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_178),
.B(n_180),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_188),
.B(n_189),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_195),
.B(n_196),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_211),
.B2(n_212),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_213),
.C(n_224),
.Y(n_227)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_204),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_205),
.C(n_206),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_209),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_223),
.B2(n_224),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_222),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_219),
.C(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_218),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_227),
.B(n_228),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_244),
.B2(n_253),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_243),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_231),
.B(n_243),
.C(n_253),
.Y(n_310)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_239),
.B2(n_240),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_234),
.B(n_241),
.C(n_242),
.Y(n_273)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g398 ( 
.A(n_235),
.Y(n_398)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_237),
.CI(n_238),
.CON(n_235),
.SN(n_235)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_236),
.B(n_237),
.C(n_238),
.Y(n_282)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_244),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g399 ( 
.A(n_244),
.Y(n_399)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_246),
.CI(n_250),
.CON(n_244),
.SN(n_244)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_245),
.B(n_246),
.C(n_250),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B(n_249),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_248),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_249),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_281)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI21xp33_ASAP7_75t_L g377 ( 
.A1(n_256),
.A2(n_378),
.B(n_379),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_286),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_257),
.B(n_286),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_274),
.C(n_285),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_258),
.B(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_273),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_266),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_260),
.B(n_266),
.C(n_273),
.Y(n_308)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_263),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_272),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_270),
.C(n_272),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_274),
.A2(n_275),
.B1(n_285),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_282),
.C(n_284),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_279),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_282),
.Y(n_283)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_308),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_297),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_297),
.C(n_308),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_294),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_295),
.C(n_296),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_298),
.B(n_300),
.C(n_301),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_305),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_303),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_310),
.B(n_311),
.Y(n_378)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_315),
.A2(n_377),
.B(n_380),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_316),
.B(n_317),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_347),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_320),
.C(n_347),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_339),
.B2(n_340),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_321),
.B(n_341),
.C(n_342),
.Y(n_375)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_324),
.B1(n_331),
.B2(n_332),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_323),
.B(n_333),
.C(n_338),
.Y(n_354)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_325),
.B(n_327),
.C(n_329),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_329),
.B2(n_330),
.Y(n_326)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_327),
.Y(n_330)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_337),
.B2(n_338),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_345),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_350),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_375),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_362),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_362),
.C(n_375),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_353),
.B(n_357),
.C(n_361),
.Y(n_390)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_361),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_364),
.B1(n_367),
.B2(n_368),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_363),
.B(n_369),
.C(n_374),
.Y(n_386)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_369),
.A2(n_370),
.B1(n_373),
.B2(n_374),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_374),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_383),
.B(n_384),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_390),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_386),
.B(n_387),
.C(n_390),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_392),
.B(n_393),
.Y(n_397)
);


endmodule