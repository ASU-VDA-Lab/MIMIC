module fake_aes_1022_n_47 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_47);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_47;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_46;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_7), .Y(n_10) );
CKINVDCx20_ASAP7_75t_R g11 ( .A(n_8), .Y(n_11) );
INVx3_ASAP7_75t_L g12 ( .A(n_3), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g13 ( .A(n_1), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_2), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_2), .Y(n_18) );
BUFx3_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_12), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_12), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_11), .Y(n_22) );
BUFx3_ASAP7_75t_L g23 ( .A(n_16), .Y(n_23) );
NOR2xp33_ASAP7_75t_L g24 ( .A(n_12), .B(n_15), .Y(n_24) );
INVx3_ASAP7_75t_L g25 ( .A(n_14), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_24), .B(n_10), .Y(n_26) );
AOI222xp33_ASAP7_75t_L g27 ( .A1(n_22), .A2(n_18), .B1(n_13), .B2(n_17), .C1(n_14), .C2(n_15), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
AND2x4_ASAP7_75t_L g29 ( .A(n_25), .B(n_15), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_25), .Y(n_30) );
OAI211xp5_ASAP7_75t_SL g31 ( .A1(n_27), .A2(n_17), .B(n_14), .C(n_20), .Y(n_31) );
OAI22xp5_ASAP7_75t_L g32 ( .A1(n_26), .A2(n_11), .B1(n_30), .B2(n_29), .Y(n_32) );
INVx8_ASAP7_75t_L g33 ( .A(n_29), .Y(n_33) );
NAND2x1p5_ASAP7_75t_L g34 ( .A(n_33), .B(n_29), .Y(n_34) );
NAND2xp5_ASAP7_75t_L g35 ( .A(n_32), .B(n_28), .Y(n_35) );
NAND3xp33_ASAP7_75t_L g36 ( .A(n_31), .B(n_28), .C(n_24), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_36), .Y(n_37) );
NAND3xp33_ASAP7_75t_SL g38 ( .A(n_34), .B(n_20), .C(n_21), .Y(n_38) );
NOR2xp33_ASAP7_75t_L g39 ( .A(n_35), .B(n_21), .Y(n_39) );
NAND4xp75_ASAP7_75t_L g40 ( .A(n_37), .B(n_0), .C(n_1), .D(n_3), .Y(n_40) );
AOI221xp5_ASAP7_75t_SL g41 ( .A1(n_39), .A2(n_25), .B1(n_19), .B2(n_23), .C(n_4), .Y(n_41) );
NOR2x1_ASAP7_75t_L g42 ( .A(n_38), .B(n_19), .Y(n_42) );
NOR4xp25_ASAP7_75t_L g43 ( .A(n_40), .B(n_19), .C(n_23), .D(n_5), .Y(n_43) );
INVx1_ASAP7_75t_L g44 ( .A(n_42), .Y(n_44) );
INVxp67_ASAP7_75t_L g45 ( .A(n_44), .Y(n_45) );
NAND3xp33_ASAP7_75t_SL g46 ( .A(n_43), .B(n_41), .C(n_23), .Y(n_46) );
AOI22xp5_ASAP7_75t_SL g47 ( .A1(n_45), .A2(n_9), .B1(n_44), .B2(n_46), .Y(n_47) );
endmodule