module real_jpeg_20830_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_255;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_202;
wire n_179;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_1),
.A2(n_40),
.B1(n_41),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_1),
.A2(n_5),
.B1(n_44),
.B2(n_46),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_46),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_2),
.A2(n_3),
.B1(n_20),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_28),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_2),
.A2(n_28),
.B1(n_40),
.B2(n_41),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_2),
.A2(n_5),
.B1(n_28),
.B2(n_44),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_SL g146 ( 
.A1(n_2),
.A2(n_24),
.B(n_31),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_2),
.B(n_21),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_L g174 ( 
.A1(n_2),
.A2(n_5),
.B(n_10),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_2),
.B(n_95),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_SL g197 ( 
.A1(n_2),
.A2(n_41),
.B(n_49),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_8),
.B1(n_19),
.B2(n_20),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_3),
.A2(n_25),
.B(n_28),
.C(n_146),
.Y(n_145)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_5),
.A2(n_10),
.B1(n_42),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_5),
.B(n_73),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_5),
.A2(n_7),
.B1(n_44),
.B2(n_53),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_5),
.A2(n_8),
.B1(n_19),
.B2(n_44),
.Y(n_148)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_53),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_8),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_8),
.A2(n_19),
.B1(n_40),
.B2(n_41),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_9),
.A2(n_20),
.B(n_22),
.C(n_30),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_101),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_99),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_84),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_15),
.B(n_84),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_61),
.C(n_67),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_16),
.B(n_61),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_60),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_17),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_17),
.A2(n_60),
.B1(n_86),
.B2(n_97),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_17),
.B(n_116),
.C(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_17),
.A2(n_60),
.B1(n_151),
.B2(n_154),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_17),
.A2(n_60),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_17),
.B(n_231),
.C(n_233),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_21),
.B(n_26),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_18),
.A2(n_21),
.B1(n_82),
.B2(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_22),
.B(n_29),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_23),
.A2(n_48),
.B(n_49),
.C(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_23),
.B(n_49),
.Y(n_58)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_24),
.A2(n_28),
.B(n_50),
.C(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_27),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_28),
.A2(n_41),
.B(n_42),
.C(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_28),
.B(n_74),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_28),
.B(n_43),
.Y(n_180)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_47),
.B2(n_59),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_34),
.A2(n_35),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_34),
.B(n_59),
.C(n_60),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_45),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_37),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_43),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_43),
.B1(n_45),
.B2(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_38),
.A2(n_43),
.B1(n_80),
.B2(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_43),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_41),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_43),
.A2(n_63),
.B(n_78),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_43),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_44),
.B(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B(n_54),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_56),
.B1(n_57),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_52),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_55),
.A2(n_66),
.B(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_56),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_61),
.A2(n_62),
.B(n_64),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_64),
.A2(n_87),
.B1(n_88),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_64),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_64),
.B(n_158),
.C(n_160),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_64),
.A2(n_142),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_67),
.A2(n_68),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_76),
.B(n_81),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_69),
.A2(n_81),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_69),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_69),
.A2(n_77),
.B1(n_106),
.B2(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_75),
.Y(n_69)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_71),
.B(n_134),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_72),
.A2(n_73),
.B1(n_135),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_74),
.A2(n_113),
.B(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_77),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_79),
.A2(n_129),
.B(n_130),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_81),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_98),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_87),
.A2(n_88),
.B1(n_116),
.B2(n_153),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_111),
.C(n_116),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_88),
.B(n_142),
.C(n_143),
.Y(n_236)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_94),
.B(n_95),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_120),
.B(n_257),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_117),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_103),
.B(n_117),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.C(n_109),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_104),
.B(n_108),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_109),
.A2(n_110),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_111),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_112),
.A2(n_114),
.B1(n_190),
.B2(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_112),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_114),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_114),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_114),
.B(n_147),
.C(n_188),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_114),
.A2(n_190),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_114),
.B(n_206),
.C(n_213),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_138),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_116),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_116),
.A2(n_127),
.B1(n_128),
.B2(n_153),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_116),
.B(n_128),
.C(n_195),
.Y(n_204)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_251),
.B(n_256),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_239),
.B(n_250),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_163),
.B(n_221),
.C(n_238),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_149),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_124),
.B(n_149),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_140),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_137),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_126),
.B(n_137),
.C(n_140),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_131),
.B2(n_132),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_128),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_127),
.B(n_132),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_128),
.B(n_173),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_148),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_138),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_180),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_147),
.A2(n_156),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_155),
.C(n_157),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_150),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_155),
.B(n_157),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_170),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_220),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_215),
.B(n_219),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_203),
.B(n_214),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_192),
.B(n_202),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_183),
.B(n_191),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_175),
.B(n_182),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_171),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_179),
.B(n_181),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_185),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_194),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_201),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_196),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_198),
.B(n_200),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_204),
.B(n_205),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_208),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_212),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_217),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_222),
.B(n_223),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_236),
.B2(n_237),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_229),
.B2(n_230),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_230),
.C(n_237),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_236),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_240),
.B(n_241),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_249),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_247),
.C(n_249),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_253),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);


endmodule