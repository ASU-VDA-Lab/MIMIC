module fake_jpeg_4336_n_265 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_265);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_28),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_33),
.B1(n_22),
.B2(n_24),
.Y(n_40)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_12),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_25),
.Y(n_43)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVxp67_ASAP7_75t_SL g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_45),
.B(n_20),
.Y(n_60)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_34),
.B(n_33),
.C(n_27),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_17),
.C(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_47),
.Y(n_65)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_57),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_22),
.B1(n_30),
.B2(n_24),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_60),
.B(n_29),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_29),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_33),
.B1(n_22),
.B2(n_20),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_24),
.B1(n_33),
.B2(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_27),
.Y(n_73)
);

AOI32xp33_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_57),
.A3(n_60),
.B1(n_61),
.B2(n_53),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_49),
.B(n_50),
.C(n_54),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_79),
.Y(n_95)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_17),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_76),
.B(n_77),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_34),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_68),
.B(n_70),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_71),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

BUFx2_ASAP7_75t_SL g74 ( 
.A(n_58),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_59),
.B1(n_52),
.B2(n_38),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_57),
.B(n_56),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_26),
.B(n_21),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_90),
.B1(n_97),
.B2(n_72),
.Y(n_105)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_86),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_53),
.B1(n_54),
.B2(n_60),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_77),
.B1(n_66),
.B2(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_47),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_88),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_91),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_65),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_71),
.B1(n_83),
.B2(n_48),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_50),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_110)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_63),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_96),
.B(n_66),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_59),
.B1(n_38),
.B2(n_52),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_98),
.A2(n_82),
.B1(n_93),
.B2(n_41),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_101),
.C(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_67),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_103),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_72),
.C(n_62),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_109),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_66),
.A3(n_64),
.B1(n_76),
.B2(n_67),
.Y(n_103)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_66),
.A3(n_64),
.B1(n_76),
.B2(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_95),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_93),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_83),
.B1(n_92),
.B2(n_41),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_75),
.B1(n_64),
.B2(n_79),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_97),
.B1(n_82),
.B2(n_93),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_80),
.B(n_91),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_75),
.C(n_68),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_116),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_26),
.C(n_39),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_97),
.C(n_89),
.Y(n_132)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_115),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_117),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_119),
.Y(n_152)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_95),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_132),
.C(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_58),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_88),
.B(n_80),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_133),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_125),
.B1(n_105),
.B2(n_111),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_131),
.Y(n_144)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_85),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_37),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_99),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_107),
.A2(n_47),
.B(n_35),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_136),
.A2(n_113),
.B1(n_37),
.B2(n_35),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_138),
.A2(n_139),
.B1(n_147),
.B2(n_153),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_116),
.B1(n_112),
.B2(n_102),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_119),
.B(n_110),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_148),
.Y(n_178)
);

NOR2x1_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_109),
.Y(n_141)
);

XOR2x1_ASAP7_75t_SL g171 ( 
.A(n_141),
.B(n_35),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_130),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_121),
.B1(n_132),
.B2(n_124),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_104),
.B1(n_103),
.B2(n_92),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_47),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_48),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_13),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_48),
.B1(n_19),
.B2(n_39),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_19),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_158),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_169),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_120),
.C(n_130),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_145),
.C(n_36),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_166),
.B(n_171),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_158),
.A2(n_134),
.B1(n_124),
.B2(n_131),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_123),
.B1(n_135),
.B2(n_39),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_168),
.A2(n_173),
.B1(n_146),
.B2(n_171),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_123),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_174),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_147),
.A2(n_39),
.B1(n_31),
.B2(n_18),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_175),
.B(n_177),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_17),
.B1(n_58),
.B2(n_13),
.Y(n_176)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_180),
.B(n_155),
.Y(n_185)
);

AO221x1_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_142),
.B1(n_157),
.B2(n_151),
.C(n_36),
.Y(n_182)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_142),
.Y(n_183)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_184),
.A2(n_188),
.B1(n_196),
.B2(n_167),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_185),
.Y(n_206)
);

XNOR2x1_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_155),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_198),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g187 ( 
.A(n_165),
.B(n_149),
.CI(n_144),
.CON(n_187),
.SN(n_187)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_187),
.B(n_190),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_163),
.A2(n_18),
.B1(n_14),
.B2(n_144),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_195),
.C(n_160),
.Y(n_202)
);

BUFx12_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_36),
.C(n_31),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_31),
.B1(n_1),
.B2(n_2),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_16),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_0),
.B(n_1),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_199),
.A2(n_178),
.B1(n_192),
.B2(n_191),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_162),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_203),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_184),
.B1(n_196),
.B2(n_187),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_207),
.C(n_210),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_173),
.Y(n_203)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_36),
.C(n_27),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_36),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_36),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_212),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_27),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_194),
.B(n_0),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_199),
.B(n_190),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_16),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_207),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_181),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_217),
.A2(n_225),
.B(n_226),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_6),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_27),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_206),
.A2(n_190),
.B(n_189),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_222),
.A2(n_210),
.B(n_208),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_213),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_227),
.B(n_4),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_0),
.Y(n_225)
);

XOR2x2_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_3),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_3),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_3),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_229),
.B(n_208),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_230),
.A2(n_235),
.B(n_239),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_231),
.B(n_238),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_200),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_237),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_27),
.C(n_4),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_234),
.A2(n_222),
.B(n_228),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_3),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_236),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_240),
.B(n_6),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_242),
.B(n_243),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_223),
.B(n_224),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_233),
.A2(n_16),
.B(n_7),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_246),
.B(n_7),
.Y(n_255)
);

OAI31xp33_ASAP7_75t_SL g247 ( 
.A1(n_235),
.A2(n_7),
.A3(n_8),
.B(n_9),
.Y(n_247)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_247),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_248),
.A2(n_234),
.B(n_232),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_251),
.B(n_254),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_249),
.C(n_244),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_247),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_255),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_248),
.B(n_16),
.Y(n_254)
);

A2O1A1O1Ixp25_ASAP7_75t_L g257 ( 
.A1(n_256),
.A2(n_8),
.B(n_9),
.C(n_10),
.D(n_11),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_257),
.A2(n_260),
.B(n_10),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_253),
.A2(n_8),
.B(n_10),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_262),
.B(n_258),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_259),
.B(n_10),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_264),
.A2(n_11),
.B(n_23),
.Y(n_265)
);


endmodule