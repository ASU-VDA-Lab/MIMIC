module fake_jpeg_28726_n_158 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_5),
.B(n_9),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_12),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_71),
.Y(n_82)
);

CKINVDCx9p33_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_73),
.A2(n_68),
.B1(n_59),
.B2(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_1),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_2),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_30),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_76),
.B(n_63),
.Y(n_80)
);

CKINVDCx9p33_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_92),
.B1(n_70),
.B2(n_53),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_74),
.B(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_84),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_76),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_72),
.A2(n_57),
.B1(n_65),
.B2(n_50),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_70),
.B1(n_73),
.B2(n_56),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_59),
.B1(n_57),
.B2(n_52),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_78),
.B1(n_32),
.B2(n_34),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_71),
.B(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_55),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_67),
.B1(n_64),
.B2(n_62),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_103),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_51),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_8),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_96),
.A2(n_109),
.B1(n_20),
.B2(n_24),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_100),
.Y(n_127)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_33),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_101),
.B(n_49),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_50),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_102),
.B(n_78),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_3),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_6),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_108),
.Y(n_115)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_109),
.A2(n_5),
.B(n_6),
.Y(n_111)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_SL g143 ( 
.A1(n_111),
.A2(n_122),
.B(n_125),
.C(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_116),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_7),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_7),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_118),
.B(n_19),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_119),
.B(n_125),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_8),
.C(n_9),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_46),
.B(n_47),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_10),
.B(n_12),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_123),
.B(n_129),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_124),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_17),
.C(n_18),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_48),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_135),
.B1(n_141),
.B2(n_143),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_112),
.B1(n_131),
.B2(n_141),
.Y(n_147)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_138),
.B(n_139),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_140),
.B(n_122),
.CI(n_119),
.CON(n_145),
.SN(n_145)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_127),
.B(n_124),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_147),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_115),
.C(n_117),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_149),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_112),
.B1(n_132),
.B2(n_142),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_143),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_152),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_152),
.C(n_150),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_144),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_147),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_148),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_146),
.Y(n_158)
);


endmodule