module fake_ariane_1828_n_2326 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_32, n_410, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_267, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_439, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_429, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_413, n_392, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_383, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_409, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_430, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_428, n_159, n_358, n_105, n_30, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_425, n_431, n_118, n_121, n_411, n_353, n_22, n_241, n_29, n_357, n_412, n_191, n_382, n_80, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_351, n_39, n_393, n_359, n_155, n_127, n_2326);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_410;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_267;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_439;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_429;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_413;
input n_392;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_409;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_430;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_425;
input n_431;
input n_118;
input n_121;
input n_411;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_2326;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_1298;
wire n_737;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_995;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_2233;
wire n_495;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2098;
wire n_661;
wire n_1751;
wire n_533;
wire n_1917;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_612;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_1442;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_1884;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_1253;
wire n_762;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_2185;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2087;
wire n_931;
wire n_669;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_489;
wire n_2294;
wire n_2274;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_471;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_2262;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_1817;
wire n_2168;
wire n_552;
wire n_2312;
wire n_670;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_1609;
wire n_1053;
wire n_600;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_2075;
wire n_1726;
wire n_1945;
wire n_1015;
wire n_545;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_501;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_1402;
wire n_957;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_1373;
wire n_1081;
wire n_742;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_1191;
wire n_618;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2320;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_453;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_519;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_1127;
wire n_556;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_1720;
wire n_663;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_1003;
wire n_701;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_671;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_97),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_157),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_415),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_397),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_342),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_312),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_174),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_225),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_367),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_71),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_62),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_395),
.Y(n_453)
);

BUFx10_ASAP7_75t_L g454 ( 
.A(n_303),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_422),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_192),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_407),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_403),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_213),
.Y(n_459)
);

BUFx10_ASAP7_75t_L g460 ( 
.A(n_235),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_239),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_159),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_5),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_382),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_23),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_288),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_170),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_396),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_438),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_333),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_251),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_18),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_143),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_345),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_91),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_69),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_278),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_149),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_410),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_5),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_439),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_412),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_371),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_361),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_247),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_59),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_105),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_274),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_223),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_10),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_329),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_290),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_58),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_197),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_386),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_378),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_282),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_108),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_291),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_180),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_229),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_131),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_38),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_173),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_313),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_293),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_286),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_344),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_409),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_160),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_88),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_168),
.Y(n_512)
);

BUFx5_ASAP7_75t_L g513 ( 
.A(n_405),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_258),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_26),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_374),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_335),
.Y(n_517)
);

CKINVDCx14_ASAP7_75t_R g518 ( 
.A(n_339),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_72),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_354),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_7),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_321),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_36),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_385),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_317),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_201),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_211),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_4),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_142),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_15),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_242),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_431),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_419),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_434),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_328),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_280),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_158),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_275),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_404),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_347),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_147),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_167),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_323),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_366),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_352),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_242),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_217),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_376),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_350),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_306),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_390),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_377),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_424),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_184),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_426),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_127),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_215),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_417),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_381),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_54),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_244),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_228),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_357),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_178),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_104),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_362),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_269),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_359),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_84),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_189),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_209),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_360),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_89),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_120),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_257),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_432),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_315),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_285),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_441),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_235),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_428),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_261),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_45),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_351),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_317),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_436),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_383),
.Y(n_587)
);

CKINVDCx14_ASAP7_75t_R g588 ( 
.A(n_258),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_338),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_332),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_372),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_433),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_41),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_183),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_302),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_233),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_398),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_312),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_231),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_256),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_212),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_257),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_184),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_216),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_341),
.Y(n_605)
);

BUFx10_ASAP7_75t_L g606 ( 
.A(n_278),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_402),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_370),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_437),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_368),
.Y(n_610)
);

BUFx10_ASAP7_75t_L g611 ( 
.A(n_82),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_77),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_399),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_107),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_364),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_114),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_336),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_429),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_337),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_394),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_24),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_270),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_435),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_267),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_294),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_401),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_126),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_236),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_388),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_16),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_413),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_146),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_406),
.Y(n_633)
);

BUFx10_ASAP7_75t_L g634 ( 
.A(n_348),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_12),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_400),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_241),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_254),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_309),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_272),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_86),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_430),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_349),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_289),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_214),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_285),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_262),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_110),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_63),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_46),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_379),
.Y(n_651)
);

BUFx2_ASAP7_75t_SL g652 ( 
.A(n_340),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_273),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_123),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_25),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_189),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_271),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_380),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_177),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_363),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_414),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_343),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_175),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_114),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_19),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_268),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_440),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_373),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_226),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_220),
.Y(n_670)
);

BUFx10_ASAP7_75t_L g671 ( 
.A(n_387),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_355),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_284),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_297),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_1),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_298),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_175),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_14),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_389),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_311),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_3),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_263),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_176),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_68),
.Y(n_684)
);

BUFx10_ASAP7_75t_L g685 ( 
.A(n_334),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_294),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_77),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_427),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_100),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_95),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_98),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_420),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_191),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_122),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_276),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_331),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_160),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_71),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_313),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_243),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_220),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_279),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_299),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_300),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_216),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_174),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_284),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_198),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_283),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_137),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_153),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_73),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_91),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_68),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_207),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_28),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_144),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_230),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_353),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_48),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_322),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_112),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_375),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_81),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_365),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_356),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_277),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_200),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_176),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_187),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_6),
.Y(n_731)
);

INVx1_ASAP7_75t_SL g732 ( 
.A(n_297),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_130),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_423),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_277),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_306),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_244),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_147),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_0),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_411),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_20),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_109),
.Y(n_742)
);

BUFx5_ASAP7_75t_L g743 ( 
.A(n_181),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_255),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_115),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_158),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_218),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_93),
.Y(n_748)
);

BUFx10_ASAP7_75t_L g749 ( 
.A(n_99),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_369),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_318),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_54),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_253),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_274),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_302),
.Y(n_755)
);

INVx1_ASAP7_75t_SL g756 ( 
.A(n_292),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_14),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_240),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_288),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_137),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_391),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_177),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_320),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_283),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_384),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_222),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_208),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_190),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_210),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_126),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_346),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_212),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_109),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_291),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_231),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_162),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_179),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_281),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_124),
.Y(n_779)
);

INVxp67_ASAP7_75t_SL g780 ( 
.A(n_425),
.Y(n_780)
);

CKINVDCx16_ASAP7_75t_R g781 ( 
.A(n_416),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_311),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_392),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_204),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_141),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_57),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_358),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_408),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_321),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_141),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_173),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_421),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_84),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_61),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_418),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_32),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_210),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_49),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_300),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_315),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_296),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_393),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_653),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_743),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_743),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_653),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_673),
.Y(n_807)
);

INVxp33_ASAP7_75t_SL g808 ( 
.A(n_632),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_588),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_673),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_789),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_775),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_743),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_781),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_743),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_797),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_743),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_743),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_743),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_789),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_524),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_743),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_461),
.Y(n_823)
);

INVxp33_ASAP7_75t_SL g824 ( 
.A(n_586),
.Y(n_824)
);

INVxp67_ASAP7_75t_SL g825 ( 
.A(n_461),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_461),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_461),
.Y(n_827)
);

INVxp67_ASAP7_75t_SL g828 ( 
.A(n_461),
.Y(n_828)
);

INVxp67_ASAP7_75t_SL g829 ( 
.A(n_473),
.Y(n_829)
);

INVxp67_ASAP7_75t_SL g830 ( 
.A(n_473),
.Y(n_830)
);

CKINVDCx16_ASAP7_75t_R g831 ( 
.A(n_454),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_443),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_634),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_563),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_463),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_466),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_475),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_477),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_480),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_634),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_473),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_492),
.Y(n_842)
);

INVxp33_ASAP7_75t_SL g843 ( 
.A(n_642),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_497),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_512),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_448),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_514),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_515),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_634),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_636),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_473),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_526),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_528),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_537),
.Y(n_854)
);

INVxp67_ASAP7_75t_SL g855 ( 
.A(n_473),
.Y(n_855)
);

INVxp33_ASAP7_75t_SL g856 ( 
.A(n_448),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_550),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_538),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_547),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_451),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_671),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_447),
.Y(n_862)
);

INVxp67_ASAP7_75t_SL g863 ( 
.A(n_511),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_564),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_455),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_567),
.Y(n_866)
);

INVxp33_ASAP7_75t_L g867 ( 
.A(n_577),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_602),
.Y(n_868)
);

INVxp33_ASAP7_75t_SL g869 ( 
.A(n_451),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_511),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_511),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_671),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_511),
.Y(n_873)
);

INVxp33_ASAP7_75t_L g874 ( 
.A(n_616),
.Y(n_874)
);

OA21x2_ASAP7_75t_L g875 ( 
.A1(n_805),
.A2(n_445),
.B(n_444),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_865),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_865),
.B(n_825),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_841),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_828),
.B(n_550),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_805),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_841),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_851),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_813),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_813),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_829),
.B(n_569),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_824),
.B(n_518),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_862),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_SL g888 ( 
.A1(n_834),
.A2(n_798),
.B1(n_449),
.B2(n_459),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_851),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_823),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_823),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_820),
.B(n_454),
.Y(n_892)
);

OA21x2_ASAP7_75t_L g893 ( 
.A1(n_815),
.A2(n_464),
.B(n_450),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_826),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_826),
.Y(n_895)
);

OAI21x1_ASAP7_75t_L g896 ( 
.A1(n_804),
.A2(n_491),
.B(n_474),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_815),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_830),
.B(n_516),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_827),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_817),
.Y(n_900)
);

BUFx12f_ASAP7_75t_L g901 ( 
.A(n_809),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_804),
.A2(n_534),
.B(n_532),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_827),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_817),
.Y(n_904)
);

BUFx2_ASAP7_75t_L g905 ( 
.A(n_809),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_870),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_820),
.B(n_454),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_855),
.B(n_535),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_818),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_870),
.Y(n_910)
);

INVx5_ASAP7_75t_L g911 ( 
.A(n_818),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_871),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_871),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_873),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_863),
.B(n_558),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_819),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_819),
.A2(n_822),
.B(n_873),
.Y(n_917)
);

OAI21x1_ASAP7_75t_L g918 ( 
.A1(n_822),
.A2(n_587),
.B(n_581),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_833),
.B(n_589),
.Y(n_919)
);

INVxp33_ASAP7_75t_SL g920 ( 
.A(n_814),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_850),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_832),
.Y(n_922)
);

NAND2xp33_ASAP7_75t_L g923 ( 
.A(n_821),
.B(n_511),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_803),
.B(n_569),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_835),
.Y(n_925)
);

BUFx12f_ASAP7_75t_L g926 ( 
.A(n_814),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_824),
.A2(n_603),
.B1(n_703),
.B2(n_580),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_833),
.B(n_590),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_836),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_837),
.Y(n_930)
);

OA21x2_ASAP7_75t_L g931 ( 
.A1(n_838),
.A2(n_605),
.B(n_591),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_839),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_867),
.B(n_460),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_842),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_844),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_840),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_884),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_921),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_887),
.Y(n_939)
);

CKINVDCx16_ASAP7_75t_R g940 ( 
.A(n_901),
.Y(n_940)
);

NOR2x1p5_ASAP7_75t_L g941 ( 
.A(n_901),
.B(n_840),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_926),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_884),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_925),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_926),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_880),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_925),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_920),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_920),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_922),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_905),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_922),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_905),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_R g954 ( 
.A(n_936),
.B(n_849),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_936),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_886),
.B(n_872),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_888),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_927),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_895),
.Y(n_959)
);

AOI21x1_ASAP7_75t_L g960 ( 
.A1(n_880),
.A2(n_617),
.B(n_607),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_929),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_929),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_930),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_883),
.Y(n_964)
);

CKINVDCx20_ASAP7_75t_R g965 ( 
.A(n_933),
.Y(n_965)
);

BUFx10_ASAP7_75t_L g966 ( 
.A(n_879),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_919),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_933),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_895),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_928),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_876),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_892),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_892),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_883),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_876),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_907),
.A2(n_843),
.B1(n_821),
.B2(n_856),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_907),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_930),
.B(n_831),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_877),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_897),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_935),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_932),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_897),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_935),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_935),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_935),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_935),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_932),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_895),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_900),
.Y(n_990)
);

BUFx8_ASAP7_75t_L g991 ( 
.A(n_879),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_879),
.B(n_849),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_879),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_967),
.B(n_923),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_946),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_978),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_964),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_946),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_970),
.B(n_993),
.Y(n_999)
);

BUFx4f_ASAP7_75t_L g1000 ( 
.A(n_950),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_966),
.Y(n_1001)
);

OAI22x1_ASAP7_75t_L g1002 ( 
.A1(n_958),
.A2(n_861),
.B1(n_816),
.B2(n_812),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_991),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_938),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_991),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_964),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_974),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_972),
.B(n_856),
.Y(n_1008)
);

NAND2xp33_ASAP7_75t_L g1009 ( 
.A(n_955),
.B(n_900),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_937),
.Y(n_1010)
);

AND2x6_ASAP7_75t_L g1011 ( 
.A(n_974),
.B(n_885),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_980),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_966),
.Y(n_1013)
);

AND2x6_ASAP7_75t_L g1014 ( 
.A(n_980),
.B(n_885),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_966),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_939),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_952),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_981),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_961),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_983),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_962),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_973),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_983),
.Y(n_1023)
);

AND2x4_ASAP7_75t_SL g1024 ( 
.A(n_965),
.B(n_662),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_951),
.B(n_846),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_963),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_992),
.B(n_924),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_988),
.B(n_885),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_956),
.B(n_869),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_990),
.Y(n_1030)
);

AND2x6_ASAP7_75t_L g1031 ( 
.A(n_990),
.B(n_885),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_944),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_939),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_982),
.B(n_934),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_947),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_937),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_953),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_937),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_943),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_959),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_971),
.B(n_861),
.Y(n_1041)
);

NOR2x1p5_ASAP7_75t_L g1042 ( 
.A(n_948),
.B(n_949),
.Y(n_1042)
);

BUFx10_ASAP7_75t_L g1043 ( 
.A(n_942),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_943),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_959),
.Y(n_1045)
);

NAND2x1p5_ASAP7_75t_L g1046 ( 
.A(n_943),
.B(n_934),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_959),
.Y(n_1047)
);

BUFx10_ASAP7_75t_L g1048 ( 
.A(n_942),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_969),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_977),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_954),
.B(n_904),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_975),
.B(n_898),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_969),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_969),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_981),
.B(n_991),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_965),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_989),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_989),
.Y(n_1058)
);

INVx4_ASAP7_75t_L g1059 ( 
.A(n_984),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_979),
.B(n_869),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_989),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_987),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_960),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_985),
.B(n_908),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_986),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_979),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_945),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_940),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_976),
.B(n_915),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_968),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_968),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_997),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1028),
.B(n_843),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1060),
.B(n_977),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_997),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1006),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1006),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_1069),
.A2(n_918),
.B(n_902),
.C(n_896),
.Y(n_1078)
);

OAI221xp5_ASAP7_75t_L g1079 ( 
.A1(n_1069),
.A2(n_860),
.B1(n_857),
.B2(n_957),
.C(n_506),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1007),
.Y(n_1080)
);

INVx8_ASAP7_75t_L g1081 ( 
.A(n_1067),
.Y(n_1081)
);

NOR2x1p5_ASAP7_75t_L g1082 ( 
.A(n_1068),
.B(n_941),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1017),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_1033),
.Y(n_1084)
);

INVxp67_ASAP7_75t_L g1085 ( 
.A(n_1050),
.Y(n_1085)
);

AO22x2_ASAP7_75t_L g1086 ( 
.A1(n_1066),
.A2(n_1056),
.B1(n_1071),
.B2(n_1055),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1060),
.B(n_874),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_1049),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_1016),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_1003),
.B(n_924),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1007),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1012),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_1004),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1019),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1021),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1026),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1012),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_1018),
.B(n_1000),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_1003),
.B(n_924),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_1049),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1005),
.B(n_924),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1034),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1052),
.B(n_808),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_1025),
.B(n_808),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1020),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_1049),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_1070),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1020),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1023),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_1070),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1000),
.A2(n_452),
.B1(n_504),
.B2(n_499),
.Y(n_1111)
);

INVxp67_ASAP7_75t_L g1112 ( 
.A(n_999),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_1013),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1023),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1030),
.Y(n_1115)
);

NAND2x1p5_ASAP7_75t_L g1116 ( 
.A(n_1005),
.B(n_881),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_1008),
.Y(n_1117)
);

AO22x2_ASAP7_75t_L g1118 ( 
.A1(n_1055),
.A2(n_624),
.B1(n_650),
.B2(n_594),
.Y(n_1118)
);

NAND2xp33_ASAP7_75t_L g1119 ( 
.A(n_1046),
.B(n_904),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1027),
.B(n_845),
.Y(n_1120)
);

OAI221xp5_ASAP7_75t_L g1121 ( 
.A1(n_996),
.A2(n_1008),
.B1(n_1022),
.B2(n_1029),
.C(n_1041),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1030),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_1037),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_1024),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_1067),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1032),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1013),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1034),
.B(n_909),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1032),
.Y(n_1129)
);

CKINVDCx8_ASAP7_75t_R g1130 ( 
.A(n_1067),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1035),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1024),
.B(n_806),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_1013),
.Y(n_1133)
);

AOI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_994),
.A2(n_723),
.B1(n_734),
.B2(n_672),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1034),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1064),
.B(n_909),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1035),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1029),
.A2(n_918),
.B(n_902),
.C(n_896),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1027),
.B(n_1001),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_995),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1040),
.Y(n_1141)
);

NAND2x1p5_ASAP7_75t_L g1142 ( 
.A(n_1068),
.B(n_881),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1040),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_998),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1062),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1001),
.B(n_847),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1036),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1022),
.B(n_507),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1038),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1009),
.B(n_529),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1045),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1039),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1044),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_1065),
.B(n_1013),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1053),
.Y(n_1155)
);

OR2x2_ASAP7_75t_SL g1156 ( 
.A(n_1067),
.B(n_614),
.Y(n_1156)
);

OR2x6_ASAP7_75t_L g1157 ( 
.A(n_1042),
.B(n_848),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1009),
.B(n_599),
.Y(n_1158)
);

OAI221xp5_ASAP7_75t_L g1159 ( 
.A1(n_1051),
.A2(n_505),
.B1(n_732),
.B2(n_756),
.C(n_686),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1011),
.B(n_916),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1053),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1047),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1010),
.Y(n_1163)
);

INVx4_ASAP7_75t_L g1164 ( 
.A(n_1015),
.Y(n_1164)
);

OR2x2_ASAP7_75t_SL g1165 ( 
.A(n_1043),
.B(n_639),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1010),
.Y(n_1166)
);

INVxp67_ASAP7_75t_L g1167 ( 
.A(n_1051),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1049),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1046),
.A2(n_665),
.B1(n_730),
.B2(n_659),
.Y(n_1169)
);

AND2x6_ASAP7_75t_L g1170 ( 
.A(n_1015),
.B(n_458),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1065),
.B(n_735),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1088),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1139),
.B(n_1015),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_1081),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1117),
.A2(n_689),
.B(n_736),
.C(n_646),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1112),
.B(n_1059),
.Y(n_1176)
);

BUFx4f_ASAP7_75t_L g1177 ( 
.A(n_1081),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1150),
.B(n_1018),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1088),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1104),
.B(n_1059),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1078),
.A2(n_1063),
.B(n_1054),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1158),
.B(n_1043),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1087),
.B(n_1102),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1082),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1119),
.A2(n_1058),
.B(n_1057),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1135),
.B(n_1011),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1103),
.B(n_1011),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1136),
.A2(n_1058),
.B(n_1057),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1076),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1073),
.B(n_1011),
.Y(n_1190)
);

OAI21xp33_ASAP7_75t_L g1191 ( 
.A1(n_1148),
.A2(n_465),
.B(n_456),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1076),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1083),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1094),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1080),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1080),
.A2(n_917),
.B(n_1061),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1121),
.A2(n_1061),
.B(n_780),
.C(n_646),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1097),
.A2(n_917),
.B(n_893),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1134),
.B(n_1048),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1120),
.B(n_1014),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_SL g1201 ( 
.A(n_1130),
.B(n_1048),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1128),
.A2(n_916),
.B(n_893),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1120),
.B(n_1014),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1079),
.A2(n_1167),
.B(n_1159),
.C(n_1171),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1160),
.A2(n_689),
.B(n_736),
.C(n_457),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1139),
.B(n_1014),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1138),
.A2(n_1031),
.B(n_1014),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1095),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1096),
.B(n_1014),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1146),
.B(n_1031),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1155),
.A2(n_1161),
.B(n_1162),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1097),
.Y(n_1212)
);

AO32x2_ASAP7_75t_L g1213 ( 
.A1(n_1086),
.A2(n_457),
.A3(n_931),
.B1(n_893),
.B2(n_875),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1146),
.B(n_1154),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1074),
.A2(n_778),
.B(n_628),
.C(n_635),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1098),
.A2(n_640),
.B(n_645),
.C(n_621),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1111),
.A2(n_1002),
.B1(n_1031),
.B2(n_754),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1093),
.B(n_1090),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1163),
.A2(n_893),
.B(n_875),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1163),
.A2(n_875),
.B(n_911),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1154),
.B(n_1031),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1166),
.A2(n_911),
.B(n_931),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1166),
.A2(n_911),
.B(n_931),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1132),
.B(n_807),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1126),
.A2(n_668),
.B(n_679),
.C(n_667),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1169),
.B(n_755),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1085),
.B(n_777),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1126),
.A2(n_725),
.B(n_726),
.C(n_719),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1084),
.B(n_1031),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1105),
.Y(n_1230)
);

AOI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1105),
.A2(n_891),
.B(n_890),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1141),
.A2(n_911),
.B(n_931),
.Y(n_1232)
);

AOI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1108),
.A2(n_891),
.B(n_890),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1143),
.A2(n_911),
.B(n_481),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_L g1235 ( 
.A(n_1123),
.B(n_498),
.C(n_442),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1145),
.B(n_810),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1108),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1147),
.A2(n_465),
.B1(n_467),
.B2(n_456),
.Y(n_1238)
);

NOR2x1_ASAP7_75t_L g1239 ( 
.A(n_1157),
.B(n_811),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1137),
.B(n_467),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1129),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1151),
.A2(n_765),
.B(n_458),
.Y(n_1242)
);

NAND3xp33_ASAP7_75t_L g1243 ( 
.A(n_1107),
.B(n_501),
.C(n_500),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1109),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_1110),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1100),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1149),
.A2(n_771),
.B(n_765),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1090),
.B(n_471),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1131),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1099),
.B(n_471),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1099),
.B(n_472),
.Y(n_1251)
);

O2A1O1Ixp33_ASAP7_75t_SL g1252 ( 
.A1(n_1152),
.A2(n_648),
.B(n_649),
.C(n_647),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1153),
.A2(n_771),
.B(n_540),
.Y(n_1253)
);

NAND3xp33_ASAP7_75t_L g1254 ( 
.A(n_1140),
.B(n_503),
.C(n_502),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1100),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1101),
.B(n_472),
.Y(n_1256)
);

BUFx12f_ASAP7_75t_L g1257 ( 
.A(n_1157),
.Y(n_1257)
);

NOR2xp67_ASAP7_75t_L g1258 ( 
.A(n_1133),
.B(n_881),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1101),
.B(n_1086),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1144),
.A2(n_750),
.B(n_740),
.Y(n_1260)
);

INVx4_ASAP7_75t_L g1261 ( 
.A(n_1133),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1124),
.B(n_460),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1109),
.A2(n_549),
.B(n_484),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1100),
.A2(n_633),
.B(n_566),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1106),
.A2(n_802),
.B(n_508),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1224),
.B(n_1089),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1180),
.B(n_1173),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_1245),
.Y(n_1268)
);

NAND2xp33_ASAP7_75t_SL g1269 ( 
.A(n_1176),
.B(n_1164),
.Y(n_1269)
);

AOI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1231),
.A2(n_1075),
.B(n_1072),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1204),
.A2(n_1125),
.B1(n_1142),
.B2(n_1127),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1193),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1199),
.B(n_1165),
.Y(n_1273)
);

NAND2x1p5_ASAP7_75t_L g1274 ( 
.A(n_1177),
.B(n_1174),
.Y(n_1274)
);

INVx4_ASAP7_75t_L g1275 ( 
.A(n_1177),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1183),
.B(n_1118),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1227),
.B(n_1156),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1189),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1226),
.B(n_1116),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1174),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1187),
.A2(n_1113),
.B1(n_1127),
.B2(n_1164),
.Y(n_1281)
);

OR2x6_ASAP7_75t_L g1282 ( 
.A(n_1257),
.B(n_1118),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1214),
.B(n_1115),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1182),
.B(n_1113),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1173),
.B(n_1106),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1197),
.A2(n_1190),
.B1(n_1191),
.B2(n_1217),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1194),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1239),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1192),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1229),
.B(n_1077),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1208),
.B(n_1091),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1184),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1241),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1218),
.B(n_1092),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1249),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1188),
.A2(n_1170),
.B(n_1122),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1201),
.B(n_1114),
.Y(n_1297)
);

CKINVDCx8_ASAP7_75t_R g1298 ( 
.A(n_1172),
.Y(n_1298)
);

BUFx8_ASAP7_75t_L g1299 ( 
.A(n_1262),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1207),
.A2(n_1168),
.B(n_1106),
.Y(n_1300)
);

CKINVDCx16_ASAP7_75t_R g1301 ( 
.A(n_1248),
.Y(n_1301)
);

OR2x6_ASAP7_75t_L g1302 ( 
.A(n_1206),
.B(n_1168),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1195),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1250),
.B(n_852),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_SL g1305 ( 
.A1(n_1175),
.A2(n_666),
.B(n_669),
.C(n_655),
.Y(n_1305)
);

INVxp67_ASAP7_75t_L g1306 ( 
.A(n_1251),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1215),
.A2(n_675),
.B(n_676),
.C(n_674),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1172),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1212),
.Y(n_1309)
);

OR2x6_ASAP7_75t_L g1310 ( 
.A(n_1259),
.B(n_1168),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1260),
.A2(n_592),
.B(n_623),
.C(n_455),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1178),
.B(n_1170),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1181),
.A2(n_1170),
.B(n_494),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_SL g1314 ( 
.A1(n_1216),
.A2(n_680),
.B(n_681),
.C(n_677),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1172),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1210),
.B(n_1200),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_SL g1317 ( 
.A(n_1256),
.B(n_485),
.C(n_476),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1179),
.Y(n_1318)
);

NAND3xp33_ASAP7_75t_L g1319 ( 
.A(n_1205),
.B(n_485),
.C(n_476),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1240),
.A2(n_767),
.B1(n_774),
.B2(n_489),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1203),
.Y(n_1321)
);

AOI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1233),
.A2(n_899),
.B(n_894),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1185),
.A2(n_1170),
.B(n_494),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1230),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1237),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1209),
.A2(n_776),
.B1(n_489),
.B2(n_486),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1254),
.A2(n_769),
.B1(n_782),
.B2(n_493),
.Y(n_1327)
);

AOI33xp33_ASAP7_75t_L g1328 ( 
.A1(n_1252),
.A2(n_700),
.A3(n_693),
.B1(n_702),
.B2(n_695),
.B3(n_687),
.Y(n_1328)
);

BUFx4f_ASAP7_75t_L g1329 ( 
.A(n_1179),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1261),
.B(n_1221),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1244),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1179),
.B(n_470),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1202),
.A2(n_543),
.B(n_462),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1236),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1238),
.A2(n_709),
.B(n_710),
.C(n_704),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1235),
.B(n_487),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1246),
.B(n_470),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1211),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1246),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1213),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1243),
.B(n_488),
.Y(n_1341)
);

O2A1O1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1225),
.A2(n_713),
.B(n_715),
.C(n_712),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1196),
.A2(n_899),
.B(n_894),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1263),
.B(n_490),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1220),
.A2(n_578),
.B(n_554),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1247),
.Y(n_1346)
);

NAND2x1p5_ASAP7_75t_L g1347 ( 
.A(n_1261),
.B(n_853),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1213),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1186),
.A2(n_782),
.B1(n_799),
.B2(n_769),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1228),
.A2(n_784),
.B1(n_770),
.B2(n_493),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1255),
.B(n_479),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1253),
.A2(n_478),
.B1(n_536),
.B2(n_460),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1213),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1264),
.B(n_1255),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1222),
.A2(n_578),
.B(n_554),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_1265),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1258),
.B(n_490),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1242),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1198),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1219),
.B(n_625),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1232),
.B(n_760),
.Y(n_1361)
);

OAI21xp33_ASAP7_75t_L g1362 ( 
.A1(n_1223),
.A2(n_764),
.B(n_762),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1338),
.B(n_1234),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1268),
.Y(n_1364)
);

INVx1_ASAP7_75t_SL g1365 ( 
.A(n_1315),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1298),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1339),
.Y(n_1367)
);

INVx5_ASAP7_75t_L g1368 ( 
.A(n_1302),
.Y(n_1368)
);

INVx5_ASAP7_75t_SL g1369 ( 
.A(n_1280),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1272),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1308),
.Y(n_1371)
);

INVx3_ASAP7_75t_SL g1372 ( 
.A(n_1275),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1329),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1274),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1267),
.B(n_762),
.Y(n_1375)
);

BUFx12f_ASAP7_75t_L g1376 ( 
.A(n_1299),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1273),
.A2(n_767),
.B1(n_768),
.B2(n_764),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1287),
.Y(n_1378)
);

INVx6_ASAP7_75t_SL g1379 ( 
.A(n_1310),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1292),
.Y(n_1380)
);

INVx5_ASAP7_75t_L g1381 ( 
.A(n_1302),
.Y(n_1381)
);

BUFx12f_ASAP7_75t_L g1382 ( 
.A(n_1299),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1280),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1278),
.Y(n_1384)
);

BUFx12f_ASAP7_75t_L g1385 ( 
.A(n_1308),
.Y(n_1385)
);

NAND2x1p5_ASAP7_75t_L g1386 ( 
.A(n_1330),
.B(n_914),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1266),
.Y(n_1387)
);

OR2x6_ASAP7_75t_L g1388 ( 
.A(n_1310),
.B(n_903),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1301),
.B(n_478),
.Y(n_1389)
);

INVx5_ASAP7_75t_L g1390 ( 
.A(n_1302),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1330),
.B(n_903),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1288),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1289),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1318),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1293),
.Y(n_1395)
);

NAND2x1_ASAP7_75t_L g1396 ( 
.A(n_1300),
.B(n_895),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1295),
.Y(n_1397)
);

INVx2_ASAP7_75t_SL g1398 ( 
.A(n_1347),
.Y(n_1398)
);

INVx1_ASAP7_75t_SL g1399 ( 
.A(n_1321),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1303),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1334),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1359),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1309),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1325),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1282),
.A2(n_478),
.B1(n_606),
.B2(n_536),
.Y(n_1405)
);

BUFx12f_ASAP7_75t_L g1406 ( 
.A(n_1304),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1324),
.Y(n_1407)
);

NAND2x1p5_ASAP7_75t_L g1408 ( 
.A(n_1285),
.B(n_878),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1331),
.B(n_721),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1297),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1284),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1291),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1306),
.B(n_536),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1354),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_1277),
.Y(n_1415)
);

BUFx4_ASAP7_75t_SL g1416 ( 
.A(n_1319),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1294),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1283),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1290),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1279),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1316),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1340),
.B(n_724),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1270),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1312),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1332),
.Y(n_1425)
);

INVx3_ASAP7_75t_SL g1426 ( 
.A(n_1337),
.Y(n_1426)
);

BUFx2_ASAP7_75t_SL g1427 ( 
.A(n_1351),
.Y(n_1427)
);

INVx5_ASAP7_75t_L g1428 ( 
.A(n_1282),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1341),
.B(n_606),
.Y(n_1429)
);

CKINVDCx6p67_ASAP7_75t_R g1430 ( 
.A(n_1276),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1333),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1286),
.A2(n_611),
.B1(n_749),
.B2(n_606),
.Y(n_1432)
);

BUFx4_ASAP7_75t_SL g1433 ( 
.A(n_1346),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1336),
.A2(n_770),
.B1(n_772),
.B2(n_768),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1360),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1269),
.Y(n_1436)
);

INVx2_ASAP7_75t_R g1437 ( 
.A(n_1358),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1281),
.Y(n_1438)
);

AO21x2_ASAP7_75t_L g1439 ( 
.A1(n_1423),
.A2(n_1296),
.B(n_1313),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1396),
.A2(n_1322),
.B(n_1343),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1435),
.A2(n_1305),
.B(n_1307),
.C(n_1314),
.Y(n_1441)
);

INVx4_ASAP7_75t_L g1442 ( 
.A(n_1385),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1363),
.A2(n_1323),
.B(n_1355),
.Y(n_1443)
);

OAI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1387),
.A2(n_1344),
.B1(n_1271),
.B2(n_1361),
.Y(n_1444)
);

AOI221xp5_ASAP7_75t_L g1445 ( 
.A1(n_1432),
.A2(n_1335),
.B1(n_1350),
.B2(n_776),
.C(n_784),
.Y(n_1445)
);

AO21x2_ASAP7_75t_L g1446 ( 
.A1(n_1422),
.A2(n_1345),
.B(n_1348),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1432),
.A2(n_1362),
.B1(n_1311),
.B2(n_1342),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1384),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1407),
.B(n_1353),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1363),
.A2(n_1362),
.B(n_1356),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1370),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_L g1452 ( 
.A(n_1429),
.B(n_1357),
.C(n_1352),
.Y(n_1452)
);

BUFx12f_ASAP7_75t_L g1453 ( 
.A(n_1376),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1382),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_SL g1455 ( 
.A1(n_1427),
.A2(n_779),
.B1(n_785),
.B2(n_773),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1434),
.A2(n_1328),
.B(n_1326),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1367),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1406),
.A2(n_1317),
.B1(n_1349),
.B2(n_685),
.Y(n_1458)
);

OA21x2_ASAP7_75t_L g1459 ( 
.A1(n_1431),
.A2(n_858),
.B(n_854),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1378),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1393),
.Y(n_1461)
);

A2O1A1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1375),
.A2(n_1320),
.B(n_654),
.C(n_670),
.Y(n_1462)
);

AOI211xp5_ASAP7_75t_L g1463 ( 
.A1(n_1377),
.A2(n_1327),
.B(n_747),
.C(n_748),
.Y(n_1463)
);

AO31x2_ASAP7_75t_L g1464 ( 
.A1(n_1400),
.A2(n_864),
.A3(n_866),
.B(n_859),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1407),
.B(n_878),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1395),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1411),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1419),
.B(n_1399),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1436),
.A2(n_654),
.B(n_637),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1402),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1438),
.A2(n_759),
.B(n_728),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1408),
.A2(n_868),
.B(n_766),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_1380),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1405),
.A2(n_779),
.B1(n_785),
.B2(n_773),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1411),
.B(n_763),
.Y(n_1475)
);

AND2x6_ASAP7_75t_L g1476 ( 
.A(n_1421),
.B(n_446),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1438),
.A2(n_790),
.B(n_786),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1386),
.A2(n_796),
.B(n_794),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1430),
.A2(n_685),
.B1(n_671),
.B2(n_611),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1404),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1386),
.A2(n_801),
.B(n_800),
.Y(n_1481)
);

CKINVDCx6p67_ASAP7_75t_R g1482 ( 
.A(n_1372),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_SL g1483 ( 
.A(n_1420),
.B(n_685),
.Y(n_1483)
);

BUFx10_ASAP7_75t_L g1484 ( 
.A(n_1373),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1397),
.A2(n_670),
.B(n_637),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1403),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1419),
.B(n_678),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1399),
.B(n_678),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1402),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1401),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1410),
.B(n_1414),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1412),
.A2(n_729),
.B(n_699),
.Y(n_1492)
);

NOR2xp67_ASAP7_75t_L g1493 ( 
.A(n_1428),
.B(n_878),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1440),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1486),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1451),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1489),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1460),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1466),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1445),
.A2(n_1405),
.B1(n_1415),
.B2(n_1375),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1489),
.B(n_1437),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1448),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1461),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1439),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1470),
.B(n_1437),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1480),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1470),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1468),
.B(n_1410),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1446),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1446),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1464),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1447),
.A2(n_1428),
.B1(n_1424),
.B2(n_1401),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1467),
.B(n_1414),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1468),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1464),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1457),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1464),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1449),
.Y(n_1518)
);

BUFx2_ASAP7_75t_SL g1519 ( 
.A(n_1476),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1449),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1439),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1491),
.B(n_1364),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1491),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1447),
.A2(n_1428),
.B1(n_1424),
.B2(n_1389),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1490),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1459),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1459),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1471),
.A2(n_1426),
.B1(n_1428),
.B2(n_1433),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1485),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1443),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1452),
.A2(n_1418),
.B1(n_1417),
.B2(n_1413),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1492),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1450),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1450),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1487),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1444),
.B(n_1418),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_1482),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1475),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1473),
.B(n_1365),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1488),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1487),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1516),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1502),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1497),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_R g1545 ( 
.A(n_1537),
.B(n_1454),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1522),
.B(n_1364),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_R g1547 ( 
.A(n_1537),
.B(n_1453),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1513),
.B(n_1392),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1513),
.B(n_1442),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1516),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1516),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1539),
.B(n_1442),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1495),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1500),
.A2(n_1477),
.B1(n_1471),
.B2(n_1445),
.Y(n_1554)
);

NOR2x1_ASAP7_75t_SL g1555 ( 
.A(n_1528),
.B(n_1519),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1539),
.B(n_1365),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1522),
.B(n_1469),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1502),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1495),
.Y(n_1559)
);

NAND2xp33_ASAP7_75t_R g1560 ( 
.A(n_1523),
.B(n_1366),
.Y(n_1560)
);

CKINVDCx16_ASAP7_75t_R g1561 ( 
.A(n_1537),
.Y(n_1561)
);

CKINVDCx16_ASAP7_75t_R g1562 ( 
.A(n_1538),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1507),
.B(n_1383),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1495),
.Y(n_1564)
);

INVxp67_ASAP7_75t_L g1565 ( 
.A(n_1507),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1520),
.B(n_1465),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1496),
.Y(n_1567)
);

CKINVDCx16_ASAP7_75t_R g1568 ( 
.A(n_1540),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1496),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1523),
.B(n_1514),
.Y(n_1570)
);

AO31x2_ASAP7_75t_L g1571 ( 
.A1(n_1509),
.A2(n_1462),
.A3(n_1469),
.B(n_1474),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1498),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1520),
.B(n_1518),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1519),
.B(n_1388),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1508),
.B(n_1372),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_1541),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1500),
.A2(n_1444),
.B1(n_1477),
.B2(n_1456),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1514),
.B(n_1421),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1498),
.Y(n_1579)
);

NAND3xp33_ASAP7_75t_SL g1580 ( 
.A(n_1528),
.B(n_1483),
.C(n_1463),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1499),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1533),
.B(n_1421),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1533),
.A2(n_1441),
.B(n_1433),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1499),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1518),
.B(n_1465),
.Y(n_1585)
);

INVxp67_ASAP7_75t_L g1586 ( 
.A(n_1534),
.Y(n_1586)
);

INVx4_ASAP7_75t_L g1587 ( 
.A(n_1505),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1525),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1535),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1503),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1501),
.Y(n_1591)
);

NOR2xp67_ASAP7_75t_L g1592 ( 
.A(n_1586),
.B(n_1534),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1586),
.Y(n_1593)
);

INVx4_ASAP7_75t_L g1594 ( 
.A(n_1561),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1553),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1587),
.B(n_1505),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1559),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1587),
.B(n_1501),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1564),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1582),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1570),
.B(n_1544),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1591),
.B(n_1494),
.Y(n_1602)
);

INVxp67_ASAP7_75t_SL g1603 ( 
.A(n_1544),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1570),
.B(n_1525),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1562),
.B(n_1494),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1551),
.B(n_1494),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1556),
.B(n_1494),
.Y(n_1607)
);

INVxp67_ASAP7_75t_SL g1608 ( 
.A(n_1565),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1582),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1590),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1567),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1565),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1580),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1563),
.B(n_1530),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1568),
.B(n_1536),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1569),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1543),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1572),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1579),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1558),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1589),
.B(n_1535),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1555),
.B(n_1536),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1581),
.B(n_1511),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1601),
.B(n_1557),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1622),
.B(n_1549),
.Y(n_1625)
);

OAI22xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1615),
.A2(n_1577),
.B1(n_1483),
.B2(n_1588),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1623),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1594),
.Y(n_1628)
);

AO21x2_ASAP7_75t_L g1629 ( 
.A1(n_1592),
.A2(n_1577),
.B(n_1580),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1610),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1593),
.A2(n_1583),
.B(n_1554),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1594),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1610),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1611),
.Y(n_1634)
);

OA21x2_ASAP7_75t_L g1635 ( 
.A1(n_1592),
.A2(n_1609),
.B(n_1600),
.Y(n_1635)
);

AOI211xp5_ASAP7_75t_L g1636 ( 
.A1(n_1613),
.A2(n_1583),
.B(n_1622),
.C(n_1474),
.Y(n_1636)
);

OAI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1608),
.A2(n_1554),
.B(n_1576),
.Y(n_1637)
);

OAI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1613),
.A2(n_1560),
.B1(n_1615),
.B2(n_1594),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1622),
.B(n_1548),
.Y(n_1639)
);

INVxp67_ASAP7_75t_L g1640 ( 
.A(n_1613),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1604),
.B(n_1584),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1623),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1622),
.B(n_1605),
.Y(n_1643)
);

OAI21xp33_ASAP7_75t_SL g1644 ( 
.A1(n_1603),
.A2(n_1542),
.B(n_1552),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1600),
.B(n_1609),
.Y(n_1645)
);

INVx4_ASAP7_75t_L g1646 ( 
.A(n_1613),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1610),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1611),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1616),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1616),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1618),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1613),
.A2(n_1578),
.B(n_1574),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1639),
.B(n_1605),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1649),
.Y(n_1654)
);

OAI211xp5_ASAP7_75t_L g1655 ( 
.A1(n_1631),
.A2(n_1637),
.B(n_1636),
.C(n_1646),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1639),
.B(n_1596),
.Y(n_1656)
);

NAND3xp33_ASAP7_75t_L g1657 ( 
.A(n_1646),
.B(n_1612),
.C(n_1609),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1629),
.A2(n_1621),
.B(n_1600),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1643),
.B(n_1596),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1643),
.B(n_1606),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1625),
.B(n_1606),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1625),
.B(n_1607),
.Y(n_1662)
);

OA332x1_ASAP7_75t_L g1663 ( 
.A1(n_1632),
.A2(n_1545),
.A3(n_1547),
.B1(n_1619),
.B2(n_1618),
.B3(n_1598),
.C1(n_1550),
.C2(n_1607),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1629),
.A2(n_1626),
.B1(n_1646),
.B2(n_1640),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1634),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1649),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1650),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1628),
.B(n_1598),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1628),
.B(n_1602),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1650),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1635),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1624),
.A2(n_1575),
.B1(n_1548),
.B2(n_1524),
.Y(n_1672)
);

NOR2x1_ASAP7_75t_L g1673 ( 
.A(n_1638),
.B(n_1619),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1644),
.B(n_1602),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1648),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1651),
.B(n_1595),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1635),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1651),
.Y(n_1678)
);

INVx4_ASAP7_75t_L g1679 ( 
.A(n_1635),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1641),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1627),
.B(n_1595),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1630),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1627),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1680),
.B(n_1642),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1679),
.B(n_1642),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1658),
.B(n_1645),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1654),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1659),
.B(n_1614),
.Y(n_1688)
);

AND2x4_ASAP7_75t_SL g1689 ( 
.A(n_1668),
.B(n_1566),
.Y(n_1689)
);

OR2x6_ASAP7_75t_L g1690 ( 
.A(n_1679),
.B(n_1652),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1654),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1665),
.B(n_1675),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1655),
.B(n_1597),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1653),
.B(n_1597),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1653),
.B(n_1599),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1656),
.B(n_1599),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1679),
.A2(n_1515),
.B1(n_1517),
.B2(n_1511),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1656),
.B(n_1630),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1683),
.B(n_1546),
.Y(n_1699)
);

BUFx3_ASAP7_75t_L g1700 ( 
.A(n_1671),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1671),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1668),
.B(n_1633),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1673),
.B(n_1633),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1674),
.B(n_1647),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1666),
.Y(n_1705)
);

AOI221x1_ASAP7_75t_L g1706 ( 
.A1(n_1657),
.A2(n_1456),
.B1(n_1409),
.B2(n_1647),
.C(n_1366),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1674),
.B(n_1573),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1666),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1677),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1677),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1669),
.B(n_1573),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1700),
.B(n_1660),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1689),
.B(n_1669),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1689),
.B(n_1660),
.Y(n_1714)
);

INVxp67_ASAP7_75t_SL g1715 ( 
.A(n_1700),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1687),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1687),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1711),
.B(n_1661),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1691),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1691),
.Y(n_1720)
);

INVx2_ASAP7_75t_SL g1721 ( 
.A(n_1700),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1699),
.B(n_1681),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1703),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1702),
.B(n_1662),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1698),
.B(n_1707),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1692),
.B(n_1676),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1693),
.B(n_1684),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1686),
.B(n_1672),
.Y(n_1728)
);

INVxp67_ASAP7_75t_L g1729 ( 
.A(n_1709),
.Y(n_1729)
);

OAI21x1_ASAP7_75t_L g1730 ( 
.A1(n_1701),
.A2(n_1664),
.B(n_1682),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1705),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1703),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1707),
.B(n_1662),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1704),
.B(n_1667),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1703),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1685),
.B(n_1670),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1708),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1709),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1710),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1704),
.B(n_1670),
.Y(n_1740)
);

XOR2x2_ASAP7_75t_L g1741 ( 
.A(n_1703),
.B(n_1455),
.Y(n_1741)
);

NAND3xp33_ASAP7_75t_L g1742 ( 
.A(n_1706),
.B(n_1701),
.C(n_1685),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1701),
.B(n_1678),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1694),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1685),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1715),
.B(n_1678),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1728),
.B(n_1727),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1725),
.B(n_1695),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1722),
.B(n_1695),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1712),
.B(n_1688),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1712),
.B(n_1724),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1715),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1734),
.B(n_1696),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1734),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1740),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1740),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1713),
.Y(n_1757)
);

INVx3_ASAP7_75t_L g1758 ( 
.A(n_1736),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1716),
.Y(n_1759)
);

INVxp67_ASAP7_75t_L g1760 ( 
.A(n_1721),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1717),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1744),
.B(n_1685),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1719),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1721),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1714),
.B(n_1690),
.Y(n_1765)
);

OAI21xp33_ASAP7_75t_L g1766 ( 
.A1(n_1728),
.A2(n_1690),
.B(n_1697),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1718),
.B(n_1690),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1720),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1741),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1741),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1726),
.B(n_1663),
.Y(n_1771)
);

INVx2_ASAP7_75t_SL g1772 ( 
.A(n_1745),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1745),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1731),
.Y(n_1774)
);

INVx4_ASAP7_75t_L g1775 ( 
.A(n_1736),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1733),
.B(n_1663),
.Y(n_1776)
);

NAND4xp25_ASAP7_75t_SL g1777 ( 
.A(n_1742),
.B(n_1458),
.C(n_1479),
.D(n_1531),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1737),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1729),
.B(n_791),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1738),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1723),
.B(n_791),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1736),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1739),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1723),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1729),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1743),
.B(n_793),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1732),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1735),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1730),
.A2(n_1425),
.B1(n_1578),
.B2(n_1517),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_SL g1790 ( 
.A(n_1741),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1712),
.Y(n_1791)
);

AND2x2_ASAP7_75t_SL g1792 ( 
.A(n_1728),
.B(n_1373),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_1712),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1712),
.Y(n_1794)
);

BUFx2_ASAP7_75t_L g1795 ( 
.A(n_1751),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1752),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1752),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1773),
.Y(n_1798)
);

AOI221xp5_ASAP7_75t_SL g1799 ( 
.A1(n_1760),
.A2(n_582),
.B1(n_561),
.B2(n_749),
.C(n_611),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1748),
.B(n_510),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1753),
.B(n_0),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1765),
.B(n_561),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1758),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1750),
.B(n_1566),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1753),
.B(n_1),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1773),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1749),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1784),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1787),
.Y(n_1809)
);

NAND4xp25_ASAP7_75t_L g1810 ( 
.A(n_1760),
.B(n_1764),
.C(n_1794),
.D(n_1791),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1788),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1790),
.Y(n_1812)
);

AOI222xp33_ASAP7_75t_L g1813 ( 
.A1(n_1770),
.A2(n_749),
.B1(n_1512),
.B2(n_1509),
.C1(n_522),
.C2(n_519),
.Y(n_1813)
);

INVxp67_ASAP7_75t_L g1814 ( 
.A(n_1769),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1746),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1746),
.Y(n_1816)
);

AND2x2_ASAP7_75t_SL g1817 ( 
.A(n_1769),
.B(n_1373),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1793),
.B(n_521),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1754),
.Y(n_1819)
);

NAND3xp33_ASAP7_75t_L g1820 ( 
.A(n_1785),
.B(n_525),
.C(n_523),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1767),
.B(n_1585),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1755),
.B(n_527),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1782),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1792),
.Y(n_1824)
);

OR2x6_ASAP7_75t_L g1825 ( 
.A(n_1770),
.B(n_1398),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1756),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1776),
.B(n_530),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1772),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1775),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1765),
.B(n_531),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1757),
.B(n_2),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1781),
.B(n_1775),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1771),
.B(n_541),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1762),
.B(n_2),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1766),
.B(n_542),
.Y(n_1835)
);

BUFx3_ASAP7_75t_L g1836 ( 
.A(n_1780),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1786),
.B(n_546),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1779),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1783),
.B(n_556),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1777),
.B(n_557),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1759),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1761),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1763),
.B(n_1768),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1774),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1778),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1789),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1747),
.B(n_560),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1751),
.B(n_562),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1753),
.B(n_3),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1752),
.Y(n_1850)
);

INVx1_ASAP7_75t_SL g1851 ( 
.A(n_1790),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1752),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1777),
.A2(n_1504),
.B1(n_1521),
.B2(n_1574),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1753),
.B(n_4),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1747),
.B(n_565),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_SL g1856 ( 
.A(n_1747),
.B(n_1383),
.Y(n_1856)
);

OAI21xp33_ASAP7_75t_L g1857 ( 
.A1(n_1851),
.A2(n_571),
.B(n_570),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1804),
.B(n_573),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1812),
.B(n_1848),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1823),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1827),
.B(n_574),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1833),
.B(n_575),
.Y(n_1862)
);

OAI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1840),
.A2(n_585),
.B(n_583),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1807),
.B(n_593),
.Y(n_1864)
);

OAI31xp33_ASAP7_75t_L g1865 ( 
.A1(n_1811),
.A2(n_1571),
.A3(n_1416),
.B(n_1374),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1798),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1806),
.Y(n_1867)
);

AOI222xp33_ASAP7_75t_L g1868 ( 
.A1(n_1808),
.A2(n_595),
.B1(n_596),
.B2(n_601),
.C1(n_600),
.C2(n_598),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1824),
.A2(n_1617),
.B1(n_1620),
.B2(n_1504),
.Y(n_1869)
);

INVxp67_ASAP7_75t_L g1870 ( 
.A(n_1856),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1801),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1805),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1849),
.Y(n_1873)
);

NOR2x1_ASAP7_75t_L g1874 ( 
.A(n_1820),
.B(n_561),
.Y(n_1874)
);

NAND4xp25_ASAP7_75t_L g1875 ( 
.A(n_1810),
.B(n_1394),
.C(n_1416),
.D(n_1371),
.Y(n_1875)
);

OAI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1828),
.A2(n_1369),
.B1(n_612),
.B2(n_622),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1846),
.A2(n_1853),
.B1(n_1825),
.B2(n_1838),
.Y(n_1877)
);

AOI222xp33_ASAP7_75t_L g1878 ( 
.A1(n_1809),
.A2(n_604),
.B1(n_627),
.B2(n_641),
.C1(n_638),
.C2(n_630),
.Y(n_1878)
);

INVx4_ASAP7_75t_L g1879 ( 
.A(n_1830),
.Y(n_1879)
);

OAI21xp33_ASAP7_75t_L g1880 ( 
.A1(n_1832),
.A2(n_656),
.B(n_644),
.Y(n_1880)
);

AOI211xp5_ASAP7_75t_L g1881 ( 
.A1(n_1803),
.A2(n_663),
.B(n_664),
.C(n_657),
.Y(n_1881)
);

INVx2_ASAP7_75t_SL g1882 ( 
.A(n_1834),
.Y(n_1882)
);

INVxp67_ASAP7_75t_L g1883 ( 
.A(n_1856),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1847),
.B(n_561),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1854),
.B(n_8),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_SL g1886 ( 
.A(n_1855),
.B(n_582),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1836),
.B(n_682),
.Y(n_1887)
);

OAI21xp33_ASAP7_75t_L g1888 ( 
.A1(n_1829),
.A2(n_684),
.B(n_683),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1831),
.B(n_690),
.Y(n_1889)
);

OAI221xp5_ASAP7_75t_L g1890 ( 
.A1(n_1799),
.A2(n_694),
.B1(n_698),
.B2(n_697),
.C(n_691),
.Y(n_1890)
);

OAI33xp33_ASAP7_75t_L g1891 ( 
.A1(n_1796),
.A2(n_707),
.A3(n_705),
.B1(n_708),
.B2(n_706),
.B3(n_701),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1821),
.B(n_711),
.Y(n_1892)
);

AOI21xp33_ASAP7_75t_L g1893 ( 
.A1(n_1799),
.A2(n_716),
.B(n_714),
.Y(n_1893)
);

AOI21xp33_ASAP7_75t_SL g1894 ( 
.A1(n_1820),
.A2(n_9),
.B(n_11),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1797),
.Y(n_1895)
);

AOI21xp33_ASAP7_75t_L g1896 ( 
.A1(n_1817),
.A2(n_718),
.B(n_717),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1800),
.B(n_720),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1825),
.Y(n_1898)
);

OAI31xp33_ASAP7_75t_L g1899 ( 
.A1(n_1835),
.A2(n_1571),
.A3(n_1526),
.B(n_1527),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1850),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1852),
.Y(n_1901)
);

OAI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1815),
.A2(n_727),
.B(n_722),
.Y(n_1902)
);

INVxp67_ASAP7_75t_L g1903 ( 
.A(n_1837),
.Y(n_1903)
);

INVx1_ASAP7_75t_SL g1904 ( 
.A(n_1818),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1819),
.B(n_731),
.Y(n_1905)
);

OAI221xp5_ASAP7_75t_L g1906 ( 
.A1(n_1816),
.A2(n_737),
.B1(n_739),
.B2(n_738),
.C(n_733),
.Y(n_1906)
);

OR2x6_ASAP7_75t_L g1907 ( 
.A(n_1802),
.B(n_1373),
.Y(n_1907)
);

OAI22xp33_ASAP7_75t_L g1908 ( 
.A1(n_1843),
.A2(n_1504),
.B1(n_1421),
.B2(n_1521),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1826),
.B(n_741),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1822),
.B(n_12),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1841),
.B(n_1571),
.Y(n_1911)
);

OAI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1842),
.A2(n_742),
.B1(n_745),
.B2(n_744),
.Y(n_1912)
);

OAI21xp33_ASAP7_75t_L g1913 ( 
.A1(n_1844),
.A2(n_751),
.B(n_746),
.Y(n_1913)
);

AOI322xp5_ASAP7_75t_L g1914 ( 
.A1(n_1845),
.A2(n_1526),
.A3(n_1527),
.B1(n_1510),
.B2(n_753),
.C1(n_752),
.C2(n_757),
.Y(n_1914)
);

NAND3xp33_ASAP7_75t_L g1915 ( 
.A(n_1813),
.B(n_582),
.C(n_758),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1839),
.Y(n_1916)
);

OAI21xp33_ASAP7_75t_L g1917 ( 
.A1(n_1851),
.A2(n_582),
.B(n_1530),
.Y(n_1917)
);

OAI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1814),
.A2(n_1481),
.B(n_1478),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1795),
.B(n_13),
.Y(n_1919)
);

NOR3xp33_ASAP7_75t_L g1920 ( 
.A(n_1851),
.B(n_468),
.C(n_453),
.Y(n_1920)
);

A2O1A1Ixp33_ASAP7_75t_L g1921 ( 
.A1(n_1851),
.A2(n_582),
.B(n_592),
.C(n_652),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1851),
.B(n_13),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1823),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1851),
.B(n_17),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1795),
.B(n_18),
.Y(n_1925)
);

OAI32xp33_ASAP7_75t_L g1926 ( 
.A1(n_1814),
.A2(n_22),
.A3(n_19),
.B1(n_21),
.B2(n_23),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1851),
.B(n_26),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1851),
.A2(n_1476),
.B1(n_1510),
.B2(n_1391),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1795),
.B(n_27),
.Y(n_1929)
);

INVxp67_ASAP7_75t_L g1930 ( 
.A(n_1795),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1795),
.B(n_27),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1851),
.B(n_28),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1795),
.B(n_29),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1851),
.B(n_29),
.Y(n_1934)
);

INVx4_ASAP7_75t_L g1935 ( 
.A(n_1830),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1851),
.B(n_30),
.Y(n_1936)
);

NOR2x1_ASAP7_75t_L g1937 ( 
.A(n_1820),
.B(n_31),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1851),
.A2(n_468),
.B(n_453),
.Y(n_1938)
);

OAI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1814),
.A2(n_1476),
.B(n_1472),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1823),
.Y(n_1940)
);

NAND3x2_ASAP7_75t_L g1941 ( 
.A(n_1795),
.B(n_32),
.C(n_33),
.Y(n_1941)
);

OAI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1814),
.A2(n_482),
.B(n_469),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1823),
.Y(n_1943)
);

INVx2_ASAP7_75t_SL g1944 ( 
.A(n_1795),
.Y(n_1944)
);

OAI322xp33_ASAP7_75t_L g1945 ( 
.A1(n_1814),
.A2(n_1529),
.A3(n_651),
.B1(n_761),
.B2(n_495),
.C1(n_783),
.C2(n_496),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1851),
.B(n_34),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1823),
.Y(n_1947)
);

AOI211xp5_ASAP7_75t_L g1948 ( 
.A1(n_1851),
.A2(n_495),
.B(n_496),
.C(n_483),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1795),
.Y(n_1949)
);

OAI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1814),
.A2(n_761),
.B(n_651),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1795),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1795),
.B(n_35),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1823),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1949),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1944),
.B(n_37),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1931),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1952),
.B(n_39),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1879),
.Y(n_1958)
);

INVx1_ASAP7_75t_SL g1959 ( 
.A(n_1919),
.Y(n_1959)
);

NAND2x1_ASAP7_75t_L g1960 ( 
.A(n_1951),
.B(n_1388),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1879),
.Y(n_1961)
);

NOR2x1_ASAP7_75t_L g1962 ( 
.A(n_1922),
.B(n_39),
.Y(n_1962)
);

NAND2x1p5_ASAP7_75t_L g1963 ( 
.A(n_1935),
.B(n_1493),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1925),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1929),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1935),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1933),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1930),
.B(n_40),
.Y(n_1968)
);

NOR2xp67_ASAP7_75t_L g1969 ( 
.A(n_1860),
.B(n_41),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1923),
.B(n_42),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1882),
.B(n_42),
.Y(n_1971)
);

INVxp67_ASAP7_75t_L g1972 ( 
.A(n_1937),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1885),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1892),
.B(n_43),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1924),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1927),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1932),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1858),
.B(n_44),
.Y(n_1978)
);

CKINVDCx16_ASAP7_75t_R g1979 ( 
.A(n_1859),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1871),
.B(n_45),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1934),
.Y(n_1981)
);

NOR2x1_ASAP7_75t_L g1982 ( 
.A(n_1936),
.B(n_47),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1946),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1872),
.B(n_47),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1940),
.B(n_49),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1943),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1873),
.B(n_1894),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1864),
.B(n_50),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1891),
.B(n_50),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1947),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1868),
.B(n_51),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1953),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1878),
.B(n_52),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1905),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1909),
.Y(n_1995)
);

NOR2x1_ASAP7_75t_L g1996 ( 
.A(n_1887),
.B(n_53),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1897),
.B(n_55),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1910),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1889),
.Y(n_1999)
);

INVx1_ASAP7_75t_SL g2000 ( 
.A(n_1862),
.Y(n_2000)
);

OR2x2_ASAP7_75t_L g2001 ( 
.A(n_1866),
.B(n_55),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1920),
.B(n_56),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1867),
.B(n_57),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1895),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1900),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1901),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1907),
.Y(n_2007)
);

INVxp67_ASAP7_75t_L g2008 ( 
.A(n_1874),
.Y(n_2008)
);

INVxp67_ASAP7_75t_SL g2009 ( 
.A(n_1941),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1902),
.B(n_1948),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1904),
.B(n_58),
.Y(n_2011)
);

INVxp67_ASAP7_75t_L g2012 ( 
.A(n_1861),
.Y(n_2012)
);

OR2x2_ASAP7_75t_L g2013 ( 
.A(n_1916),
.B(n_1942),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_1950),
.B(n_59),
.Y(n_2014)
);

INVx1_ASAP7_75t_SL g2015 ( 
.A(n_1896),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1881),
.B(n_60),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1857),
.B(n_60),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1912),
.B(n_61),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1898),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1926),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1903),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1938),
.B(n_63),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1945),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1906),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1913),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1890),
.Y(n_2026)
);

OAI21x1_ASAP7_75t_SL g2027 ( 
.A1(n_1876),
.A2(n_64),
.B(n_65),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1915),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1870),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1883),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1921),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1880),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_L g2033 ( 
.A(n_1875),
.B(n_64),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1863),
.B(n_1484),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_L g2035 ( 
.A(n_1979),
.B(n_1888),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1969),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1969),
.Y(n_2037)
);

NAND3xp33_ASAP7_75t_L g2038 ( 
.A(n_1972),
.B(n_1914),
.C(n_1917),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1961),
.B(n_1877),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1959),
.B(n_1893),
.Y(n_2040)
);

NOR2x1_ASAP7_75t_L g2041 ( 
.A(n_1966),
.B(n_1884),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1962),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1982),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1956),
.B(n_1886),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1964),
.B(n_1918),
.Y(n_2045)
);

INVx1_ASAP7_75t_SL g2046 ( 
.A(n_1955),
.Y(n_2046)
);

NOR2xp33_ASAP7_75t_L g2047 ( 
.A(n_1965),
.B(n_1928),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1982),
.Y(n_2048)
);

INVxp67_ASAP7_75t_SL g2049 ( 
.A(n_1957),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1967),
.B(n_1939),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2003),
.Y(n_2051)
);

OAI211xp5_ASAP7_75t_SL g2052 ( 
.A1(n_2029),
.A2(n_1899),
.B(n_1869),
.C(n_1865),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2001),
.Y(n_2053)
);

OAI21xp5_ASAP7_75t_L g2054 ( 
.A1(n_2009),
.A2(n_1911),
.B(n_1908),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1954),
.B(n_66),
.Y(n_2055)
);

CKINVDCx16_ASAP7_75t_R g2056 ( 
.A(n_2010),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1973),
.B(n_67),
.Y(n_2057)
);

OR2x2_ASAP7_75t_L g2058 ( 
.A(n_2030),
.B(n_67),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1970),
.B(n_69),
.Y(n_2059)
);

NOR3xp33_ASAP7_75t_L g2060 ( 
.A(n_2012),
.B(n_788),
.C(n_787),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2011),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1968),
.B(n_70),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_2027),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1985),
.B(n_72),
.Y(n_2064)
);

AOI21xp33_ASAP7_75t_L g2065 ( 
.A1(n_1998),
.A2(n_1987),
.B(n_2000),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1986),
.B(n_73),
.Y(n_2066)
);

AOI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_1971),
.A2(n_1993),
.B(n_1991),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1994),
.B(n_74),
.Y(n_2068)
);

HB1xp67_ASAP7_75t_L g2069 ( 
.A(n_2020),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1996),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1990),
.B(n_75),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1997),
.Y(n_2072)
);

OR2x2_ASAP7_75t_L g2073 ( 
.A(n_1992),
.B(n_75),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1988),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1974),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2018),
.Y(n_2076)
);

NAND2x1_ASAP7_75t_L g2077 ( 
.A(n_2004),
.B(n_76),
.Y(n_2077)
);

AND3x1_ASAP7_75t_L g2078 ( 
.A(n_2033),
.B(n_76),
.C(n_78),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1978),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1995),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2015),
.B(n_78),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_2005),
.B(n_79),
.Y(n_2082)
);

OA21x2_ASAP7_75t_L g2083 ( 
.A1(n_2006),
.A2(n_792),
.B(n_788),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1975),
.B(n_79),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1980),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1984),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1976),
.B(n_80),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1963),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2022),
.Y(n_2089)
);

AOI21xp33_ASAP7_75t_L g2090 ( 
.A1(n_2031),
.A2(n_795),
.B(n_509),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2013),
.Y(n_2091)
);

AOI22xp33_ASAP7_75t_L g2092 ( 
.A1(n_1977),
.A2(n_1506),
.B1(n_1379),
.B2(n_1532),
.Y(n_2092)
);

NOR2xp33_ASAP7_75t_L g2093 ( 
.A(n_1981),
.B(n_82),
.Y(n_2093)
);

NAND3xp33_ASAP7_75t_L g2094 ( 
.A(n_1983),
.B(n_551),
.C(n_446),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1989),
.B(n_83),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2002),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_2016),
.B(n_85),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_L g2098 ( 
.A(n_2021),
.B(n_85),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_2032),
.B(n_86),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2017),
.B(n_1999),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_2023),
.B(n_87),
.Y(n_2101)
);

NOR2xp33_ASAP7_75t_L g2102 ( 
.A(n_2014),
.B(n_87),
.Y(n_2102)
);

AOI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_2026),
.A2(n_1506),
.B1(n_1532),
.B2(n_1368),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2019),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2025),
.B(n_89),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2024),
.B(n_90),
.Y(n_2106)
);

NOR2xp33_ASAP7_75t_L g2107 ( 
.A(n_2034),
.B(n_90),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2028),
.Y(n_2108)
);

NAND3xp33_ASAP7_75t_L g2109 ( 
.A(n_2007),
.B(n_551),
.C(n_446),
.Y(n_2109)
);

OR2x6_ASAP7_75t_L g2110 ( 
.A(n_2008),
.B(n_446),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1960),
.B(n_92),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1979),
.B(n_94),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_1979),
.B(n_94),
.Y(n_2113)
);

NOR3x1_ASAP7_75t_L g2114 ( 
.A(n_2009),
.B(n_95),
.C(n_96),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1979),
.B(n_96),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1979),
.Y(n_2116)
);

NAND4xp25_ASAP7_75t_L g2117 ( 
.A(n_2029),
.B(n_101),
.C(n_97),
.D(n_99),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1979),
.B(n_101),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1979),
.Y(n_2119)
);

NAND2x1_ASAP7_75t_L g2120 ( 
.A(n_1958),
.B(n_102),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1979),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1979),
.B(n_103),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1979),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1979),
.B(n_103),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1979),
.B(n_104),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1979),
.B(n_105),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1979),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1979),
.Y(n_2128)
);

OR2x2_ASAP7_75t_L g2129 ( 
.A(n_1979),
.B(n_106),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1979),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1979),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1979),
.Y(n_2132)
);

NOR2xp33_ASAP7_75t_L g2133 ( 
.A(n_2056),
.B(n_110),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2112),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2113),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2118),
.Y(n_2136)
);

NOR2x1_ASAP7_75t_L g2137 ( 
.A(n_2116),
.B(n_111),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2056),
.B(n_112),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2129),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2119),
.Y(n_2140)
);

NAND4xp25_ASAP7_75t_L g2141 ( 
.A(n_2121),
.B(n_2123),
.C(n_2128),
.D(n_2127),
.Y(n_2141)
);

OAI221xp5_ASAP7_75t_L g2142 ( 
.A1(n_2046),
.A2(n_533),
.B1(n_539),
.B2(n_520),
.C(n_517),
.Y(n_2142)
);

NOR2xp33_ASAP7_75t_L g2143 ( 
.A(n_2131),
.B(n_113),
.Y(n_2143)
);

INVxp67_ASAP7_75t_SL g2144 ( 
.A(n_2130),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_2114),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_SL g2146 ( 
.A(n_2132),
.B(n_2091),
.Y(n_2146)
);

INVx3_ASAP7_75t_L g2147 ( 
.A(n_2077),
.Y(n_2147)
);

AOI211xp5_ASAP7_75t_L g2148 ( 
.A1(n_2065),
.A2(n_118),
.B(n_116),
.C(n_117),
.Y(n_2148)
);

O2A1O1Ixp33_ASAP7_75t_L g2149 ( 
.A1(n_2069),
.A2(n_119),
.B(n_117),
.C(n_118),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_SL g2150 ( 
.A(n_2115),
.B(n_513),
.Y(n_2150)
);

NAND3xp33_ASAP7_75t_L g2151 ( 
.A(n_2104),
.B(n_551),
.C(n_446),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2035),
.B(n_121),
.Y(n_2152)
);

INVx1_ASAP7_75t_SL g2153 ( 
.A(n_2122),
.Y(n_2153)
);

AOI21xp5_ASAP7_75t_L g2154 ( 
.A1(n_2124),
.A2(n_122),
.B(n_123),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2062),
.B(n_2120),
.Y(n_2155)
);

NAND3xp33_ASAP7_75t_L g2156 ( 
.A(n_2125),
.B(n_572),
.C(n_551),
.Y(n_2156)
);

NAND3xp33_ASAP7_75t_L g2157 ( 
.A(n_2126),
.B(n_572),
.C(n_551),
.Y(n_2157)
);

NAND4xp25_ASAP7_75t_SL g2158 ( 
.A(n_2080),
.B(n_128),
.C(n_125),
.D(n_127),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2042),
.Y(n_2159)
);

XOR2x2_ASAP7_75t_L g2160 ( 
.A(n_2078),
.B(n_128),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2043),
.Y(n_2161)
);

O2A1O1Ixp33_ASAP7_75t_L g2162 ( 
.A1(n_2048),
.A2(n_2070),
.B(n_2095),
.C(n_2101),
.Y(n_2162)
);

NAND3xp33_ASAP7_75t_L g2163 ( 
.A(n_2093),
.B(n_608),
.C(n_572),
.Y(n_2163)
);

A2O1A1Ixp33_ASAP7_75t_L g2164 ( 
.A1(n_2098),
.A2(n_545),
.B(n_548),
.C(n_544),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2082),
.B(n_129),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_2117),
.B(n_130),
.Y(n_2166)
);

AND2x4_ASAP7_75t_L g2167 ( 
.A(n_2055),
.B(n_132),
.Y(n_2167)
);

NOR3xp33_ASAP7_75t_L g2168 ( 
.A(n_2040),
.B(n_553),
.C(n_552),
.Y(n_2168)
);

AOI211xp5_ASAP7_75t_L g2169 ( 
.A1(n_2039),
.A2(n_135),
.B(n_133),
.C(n_134),
.Y(n_2169)
);

NOR2xp33_ASAP7_75t_L g2170 ( 
.A(n_2051),
.B(n_136),
.Y(n_2170)
);

AOI211x1_ASAP7_75t_SL g2171 ( 
.A1(n_2054),
.A2(n_140),
.B(n_138),
.C(n_139),
.Y(n_2171)
);

NOR3xp33_ASAP7_75t_L g2172 ( 
.A(n_2036),
.B(n_559),
.C(n_555),
.Y(n_2172)
);

NOR2x1_ASAP7_75t_L g2173 ( 
.A(n_2073),
.B(n_138),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2066),
.B(n_139),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2059),
.Y(n_2175)
);

NAND4xp25_ASAP7_75t_L g2176 ( 
.A(n_2108),
.B(n_143),
.C(n_140),
.D(n_142),
.Y(n_2176)
);

OAI211xp5_ASAP7_75t_SL g2177 ( 
.A1(n_2045),
.A2(n_146),
.B(n_144),
.C(n_145),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2071),
.B(n_145),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2049),
.B(n_148),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2064),
.Y(n_2180)
);

NOR3xp33_ASAP7_75t_L g2181 ( 
.A(n_2037),
.B(n_576),
.C(n_568),
.Y(n_2181)
);

NOR3xp33_ASAP7_75t_L g2182 ( 
.A(n_2081),
.B(n_584),
.C(n_579),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2099),
.Y(n_2183)
);

NOR2xp33_ASAP7_75t_L g2184 ( 
.A(n_2053),
.B(n_2058),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_2068),
.B(n_150),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2089),
.B(n_151),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2102),
.B(n_2072),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2107),
.B(n_151),
.Y(n_2188)
);

A2O1A1Ixp33_ASAP7_75t_SL g2189 ( 
.A1(n_2159),
.A2(n_2060),
.B(n_2088),
.C(n_2086),
.Y(n_2189)
);

AOI221x1_ASAP7_75t_L g2190 ( 
.A1(n_2141),
.A2(n_2057),
.B1(n_2087),
.B2(n_2084),
.C(n_2085),
.Y(n_2190)
);

AOI221xp5_ASAP7_75t_L g2191 ( 
.A1(n_2162),
.A2(n_2052),
.B1(n_2074),
.B2(n_2079),
.C(n_2075),
.Y(n_2191)
);

NAND4xp25_ASAP7_75t_L g2192 ( 
.A(n_2171),
.B(n_2041),
.C(n_2038),
.D(n_2047),
.Y(n_2192)
);

AOI221xp5_ASAP7_75t_L g2193 ( 
.A1(n_2133),
.A2(n_2067),
.B1(n_2061),
.B2(n_2063),
.C(n_2050),
.Y(n_2193)
);

O2A1O1Ixp33_ASAP7_75t_L g2194 ( 
.A1(n_2138),
.A2(n_2100),
.B(n_2083),
.C(n_2096),
.Y(n_2194)
);

OAI211xp5_ASAP7_75t_SL g2195 ( 
.A1(n_2146),
.A2(n_2041),
.B(n_2044),
.C(n_2076),
.Y(n_2195)
);

AOI211xp5_ASAP7_75t_SL g2196 ( 
.A1(n_2144),
.A2(n_2105),
.B(n_2097),
.C(n_2090),
.Y(n_2196)
);

INVx1_ASAP7_75t_SL g2197 ( 
.A(n_2174),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_R g2198 ( 
.A(n_2140),
.B(n_2106),
.Y(n_2198)
);

NAND4xp25_ASAP7_75t_L g2199 ( 
.A(n_2147),
.B(n_2094),
.C(n_2109),
.D(n_2111),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2160),
.Y(n_2200)
);

AOI221xp5_ASAP7_75t_L g2201 ( 
.A1(n_2139),
.A2(n_2092),
.B1(n_2103),
.B2(n_2110),
.C(n_608),
.Y(n_2201)
);

OAI311xp33_ASAP7_75t_L g2202 ( 
.A1(n_2155),
.A2(n_2110),
.A3(n_154),
.B1(n_152),
.C1(n_153),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2167),
.B(n_2137),
.Y(n_2203)
);

AOI221x1_ASAP7_75t_L g2204 ( 
.A1(n_2161),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.C(n_157),
.Y(n_2204)
);

AOI221xp5_ASAP7_75t_L g2205 ( 
.A1(n_2134),
.A2(n_608),
.B1(n_609),
.B2(n_610),
.C(n_597),
.Y(n_2205)
);

AOI21xp5_ASAP7_75t_SL g2206 ( 
.A1(n_2149),
.A2(n_161),
.B(n_163),
.Y(n_2206)
);

OAI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_2143),
.A2(n_1381),
.B1(n_1390),
.B2(n_1368),
.Y(n_2207)
);

NAND3xp33_ASAP7_75t_SL g2208 ( 
.A(n_2153),
.B(n_615),
.C(n_613),
.Y(n_2208)
);

AOI21xp5_ASAP7_75t_L g2209 ( 
.A1(n_2158),
.A2(n_163),
.B(n_164),
.Y(n_2209)
);

AOI221xp5_ASAP7_75t_L g2210 ( 
.A1(n_2135),
.A2(n_620),
.B1(n_626),
.B2(n_619),
.C(n_618),
.Y(n_2210)
);

NOR2xp33_ASAP7_75t_L g2211 ( 
.A(n_2177),
.B(n_165),
.Y(n_2211)
);

NAND4xp75_ASAP7_75t_L g2212 ( 
.A(n_2173),
.B(n_169),
.C(n_166),
.D(n_168),
.Y(n_2212)
);

OAI21xp33_ASAP7_75t_L g2213 ( 
.A1(n_2145),
.A2(n_631),
.B(n_629),
.Y(n_2213)
);

OAI22xp5_ASAP7_75t_L g2214 ( 
.A1(n_2148),
.A2(n_1381),
.B1(n_1390),
.B2(n_1368),
.Y(n_2214)
);

AOI221xp5_ASAP7_75t_L g2215 ( 
.A1(n_2136),
.A2(n_2184),
.B1(n_2182),
.B2(n_2168),
.C(n_2180),
.Y(n_2215)
);

AOI22xp33_ASAP7_75t_L g2216 ( 
.A1(n_2183),
.A2(n_895),
.B1(n_910),
.B2(n_906),
.Y(n_2216)
);

OAI321xp33_ASAP7_75t_L g2217 ( 
.A1(n_2187),
.A2(n_171),
.A3(n_172),
.B1(n_179),
.B2(n_180),
.C(n_181),
.Y(n_2217)
);

AOI221xp5_ASAP7_75t_L g2218 ( 
.A1(n_2175),
.A2(n_660),
.B1(n_661),
.B2(n_658),
.C(n_643),
.Y(n_2218)
);

OAI21xp33_ASAP7_75t_SL g2219 ( 
.A1(n_2170),
.A2(n_2152),
.B(n_2186),
.Y(n_2219)
);

AOI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_2164),
.A2(n_182),
.B(n_185),
.Y(n_2220)
);

AOI22xp33_ASAP7_75t_L g2221 ( 
.A1(n_2150),
.A2(n_906),
.B1(n_912),
.B2(n_910),
.Y(n_2221)
);

OAI22xp33_ASAP7_75t_SL g2222 ( 
.A1(n_2179),
.A2(n_692),
.B1(n_696),
.B2(n_688),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_2198),
.Y(n_2223)
);

AOI21xp33_ASAP7_75t_L g2224 ( 
.A1(n_2194),
.A2(n_2157),
.B(n_2156),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_L g2225 ( 
.A(n_2203),
.B(n_2176),
.Y(n_2225)
);

AOI221xp5_ASAP7_75t_L g2226 ( 
.A1(n_2222),
.A2(n_2181),
.B1(n_2172),
.B2(n_2154),
.C(n_2163),
.Y(n_2226)
);

NOR4xp25_ASAP7_75t_L g2227 ( 
.A(n_2195),
.B(n_2178),
.C(n_2165),
.D(n_2185),
.Y(n_2227)
);

OAI321xp33_ASAP7_75t_L g2228 ( 
.A1(n_2192),
.A2(n_2151),
.A3(n_2169),
.B1(n_2166),
.B2(n_2188),
.C(n_2142),
.Y(n_2228)
);

AO22x2_ASAP7_75t_L g2229 ( 
.A1(n_2212),
.A2(n_190),
.B1(n_186),
.B2(n_188),
.Y(n_2229)
);

AOI211xp5_ASAP7_75t_L g2230 ( 
.A1(n_2208),
.A2(n_195),
.B(n_193),
.C(n_194),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2196),
.B(n_194),
.Y(n_2231)
);

A2O1A1Ixp33_ASAP7_75t_L g2232 ( 
.A1(n_2200),
.A2(n_197),
.B(n_195),
.C(n_196),
.Y(n_2232)
);

AOI211xp5_ASAP7_75t_L g2233 ( 
.A1(n_2189),
.A2(n_2193),
.B(n_2213),
.C(n_2191),
.Y(n_2233)
);

AOI21xp5_ASAP7_75t_L g2234 ( 
.A1(n_2209),
.A2(n_196),
.B(n_198),
.Y(n_2234)
);

CKINVDCx5p33_ASAP7_75t_R g2235 ( 
.A(n_2197),
.Y(n_2235)
);

NAND4xp25_ASAP7_75t_L g2236 ( 
.A(n_2190),
.B(n_201),
.C(n_199),
.D(n_200),
.Y(n_2236)
);

OAI211xp5_ASAP7_75t_SL g2237 ( 
.A1(n_2215),
.A2(n_203),
.B(n_199),
.C(n_202),
.Y(n_2237)
);

AOI322xp5_ASAP7_75t_L g2238 ( 
.A1(n_2219),
.A2(n_202),
.A3(n_203),
.B1(n_204),
.B2(n_205),
.C1(n_206),
.C2(n_208),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2229),
.B(n_2211),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2229),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2235),
.Y(n_2241)
);

NAND4xp75_ASAP7_75t_L g2242 ( 
.A(n_2231),
.B(n_2204),
.C(n_2220),
.D(n_2205),
.Y(n_2242)
);

AOI221xp5_ASAP7_75t_L g2243 ( 
.A1(n_2227),
.A2(n_2206),
.B1(n_2201),
.B2(n_2199),
.C(n_2202),
.Y(n_2243)
);

AOI221xp5_ASAP7_75t_L g2244 ( 
.A1(n_2225),
.A2(n_2221),
.B1(n_2216),
.B2(n_2218),
.C(n_2210),
.Y(n_2244)
);

NOR2xp33_ASAP7_75t_L g2245 ( 
.A(n_2236),
.B(n_2217),
.Y(n_2245)
);

AOI31xp33_ASAP7_75t_L g2246 ( 
.A1(n_2223),
.A2(n_2214),
.A3(n_2207),
.B(n_223),
.Y(n_2246)
);

AOI21xp5_ASAP7_75t_L g2247 ( 
.A1(n_2233),
.A2(n_219),
.B(n_221),
.Y(n_2247)
);

OAI211xp5_ASAP7_75t_SL g2248 ( 
.A1(n_2226),
.A2(n_228),
.B(n_224),
.C(n_227),
.Y(n_2248)
);

AOI22xp33_ASAP7_75t_L g2249 ( 
.A1(n_2234),
.A2(n_906),
.B1(n_912),
.B2(n_910),
.Y(n_2249)
);

NOR2x1_ASAP7_75t_L g2250 ( 
.A(n_2241),
.B(n_2232),
.Y(n_2250)
);

HB1xp67_ASAP7_75t_L g2251 ( 
.A(n_2240),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2239),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2243),
.B(n_2230),
.Y(n_2253)
);

AOI211xp5_ASAP7_75t_L g2254 ( 
.A1(n_2245),
.A2(n_2228),
.B(n_2224),
.C(n_2237),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2242),
.B(n_2238),
.Y(n_2255)
);

AND2x4_ASAP7_75t_L g2256 ( 
.A(n_2247),
.B(n_227),
.Y(n_2256)
);

NOR3xp33_ASAP7_75t_L g2257 ( 
.A(n_2248),
.B(n_229),
.C(n_230),
.Y(n_2257)
);

A2O1A1Ixp33_ASAP7_75t_L g2258 ( 
.A1(n_2244),
.A2(n_234),
.B(n_232),
.C(n_233),
.Y(n_2258)
);

AOI21xp5_ASAP7_75t_L g2259 ( 
.A1(n_2255),
.A2(n_2246),
.B(n_2249),
.Y(n_2259)
);

CKINVDCx5p33_ASAP7_75t_R g2260 ( 
.A(n_2252),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2250),
.B(n_232),
.Y(n_2261)
);

CKINVDCx5p33_ASAP7_75t_R g2262 ( 
.A(n_2253),
.Y(n_2262)
);

CKINVDCx5p33_ASAP7_75t_R g2263 ( 
.A(n_2256),
.Y(n_2263)
);

HB1xp67_ASAP7_75t_L g2264 ( 
.A(n_2257),
.Y(n_2264)
);

BUFx2_ASAP7_75t_L g2265 ( 
.A(n_2258),
.Y(n_2265)
);

BUFx6f_ASAP7_75t_L g2266 ( 
.A(n_2254),
.Y(n_2266)
);

NAND3xp33_ASAP7_75t_L g2267 ( 
.A(n_2251),
.B(n_913),
.C(n_912),
.Y(n_2267)
);

INVxp67_ASAP7_75t_L g2268 ( 
.A(n_2261),
.Y(n_2268)
);

OAI22xp5_ASAP7_75t_L g2269 ( 
.A1(n_2260),
.A2(n_913),
.B1(n_912),
.B2(n_882),
.Y(n_2269)
);

NOR3xp33_ASAP7_75t_SL g2270 ( 
.A(n_2262),
.B(n_237),
.C(n_238),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2263),
.Y(n_2271)
);

OAI22x1_ASAP7_75t_L g2272 ( 
.A1(n_2265),
.A2(n_245),
.B1(n_240),
.B2(n_241),
.Y(n_2272)
);

INVx3_ASAP7_75t_L g2273 ( 
.A(n_2266),
.Y(n_2273)
);

AO22x2_ASAP7_75t_L g2274 ( 
.A1(n_2259),
.A2(n_249),
.B1(n_246),
.B2(n_248),
.Y(n_2274)
);

XNOR2x1_ASAP7_75t_L g2275 ( 
.A(n_2266),
.B(n_248),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2266),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2264),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2267),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2274),
.Y(n_2279)
);

OAI21xp5_ASAP7_75t_L g2280 ( 
.A1(n_2268),
.A2(n_250),
.B(n_252),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2274),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2273),
.Y(n_2282)
);

AOI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_2271),
.A2(n_513),
.B1(n_889),
.B2(n_878),
.Y(n_2283)
);

HB1xp67_ASAP7_75t_L g2284 ( 
.A(n_2276),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2270),
.B(n_2277),
.Y(n_2285)
);

NOR2x1p5_ASAP7_75t_L g2286 ( 
.A(n_2278),
.B(n_259),
.Y(n_2286)
);

INVx1_ASAP7_75t_SL g2287 ( 
.A(n_2275),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2284),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2279),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2281),
.Y(n_2290)
);

INVx3_ASAP7_75t_L g2291 ( 
.A(n_2282),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2286),
.Y(n_2292)
);

HB1xp67_ASAP7_75t_L g2293 ( 
.A(n_2285),
.Y(n_2293)
);

INVx3_ASAP7_75t_L g2294 ( 
.A(n_2287),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2280),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2283),
.Y(n_2296)
);

NAND3xp33_ASAP7_75t_L g2297 ( 
.A(n_2289),
.B(n_2269),
.C(n_2272),
.Y(n_2297)
);

NOR2x1_ASAP7_75t_L g2298 ( 
.A(n_2291),
.B(n_2294),
.Y(n_2298)
);

OAI21xp5_ASAP7_75t_L g2299 ( 
.A1(n_2290),
.A2(n_2293),
.B(n_2294),
.Y(n_2299)
);

CKINVDCx20_ASAP7_75t_R g2300 ( 
.A(n_2292),
.Y(n_2300)
);

HB1xp67_ASAP7_75t_L g2301 ( 
.A(n_2295),
.Y(n_2301)
);

OAI22xp5_ASAP7_75t_SL g2302 ( 
.A1(n_2296),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_2302)
);

OAI22xp5_ASAP7_75t_SL g2303 ( 
.A1(n_2288),
.A2(n_265),
.B1(n_266),
.B2(n_268),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2298),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2301),
.Y(n_2305)
);

OR2x6_ASAP7_75t_L g2306 ( 
.A(n_2299),
.B(n_2297),
.Y(n_2306)
);

OAI21xp5_ASAP7_75t_L g2307 ( 
.A1(n_2300),
.A2(n_270),
.B(n_271),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2305),
.B(n_2303),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2304),
.Y(n_2309)
);

OAI22xp5_ASAP7_75t_L g2310 ( 
.A1(n_2306),
.A2(n_2302),
.B1(n_286),
.B2(n_287),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2307),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2305),
.Y(n_2312)
);

INVxp67_ASAP7_75t_L g2313 ( 
.A(n_2312),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2309),
.Y(n_2314)
);

AOI222xp33_ASAP7_75t_SL g2315 ( 
.A1(n_2310),
.A2(n_295),
.B1(n_299),
.B2(n_301),
.C1(n_303),
.C2(n_304),
.Y(n_2315)
);

AOI22xp33_ASAP7_75t_SL g2316 ( 
.A1(n_2308),
.A2(n_301),
.B1(n_304),
.B2(n_305),
.Y(n_2316)
);

XNOR2xp5_ASAP7_75t_L g2317 ( 
.A(n_2311),
.B(n_305),
.Y(n_2317)
);

AOI22xp5_ASAP7_75t_SL g2318 ( 
.A1(n_2313),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_2318)
);

AOI22xp33_ASAP7_75t_L g2319 ( 
.A1(n_2314),
.A2(n_307),
.B1(n_308),
.B2(n_310),
.Y(n_2319)
);

AOI22xp5_ASAP7_75t_SL g2320 ( 
.A1(n_2317),
.A2(n_314),
.B1(n_316),
.B2(n_318),
.Y(n_2320)
);

AOI22xp33_ASAP7_75t_L g2321 ( 
.A1(n_2316),
.A2(n_316),
.B1(n_319),
.B2(n_322),
.Y(n_2321)
);

AO21x2_ASAP7_75t_L g2322 ( 
.A1(n_2320),
.A2(n_2315),
.B(n_319),
.Y(n_2322)
);

AND3x1_ASAP7_75t_L g2323 ( 
.A(n_2321),
.B(n_324),
.C(n_325),
.Y(n_2323)
);

OAI21xp5_ASAP7_75t_L g2324 ( 
.A1(n_2318),
.A2(n_2319),
.B(n_324),
.Y(n_2324)
);

AOI22xp5_ASAP7_75t_L g2325 ( 
.A1(n_2323),
.A2(n_325),
.B1(n_326),
.B2(n_327),
.Y(n_2325)
);

AOI211xp5_ASAP7_75t_L g2326 ( 
.A1(n_2325),
.A2(n_2324),
.B(n_2322),
.C(n_330),
.Y(n_2326)
);


endmodule