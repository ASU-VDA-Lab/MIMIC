module fake_jpeg_17621_n_124 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_124);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_56),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_60),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_45),
.Y(n_61)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_48),
.B1(n_51),
.B2(n_47),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_72),
.B1(n_73),
.B2(n_3),
.Y(n_85)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_20),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_51),
.B1(n_50),
.B2(n_44),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_49),
.B1(n_46),
.B2(n_42),
.Y(n_73)
);

CKINVDCx12_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_49),
.Y(n_76)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_82),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_66),
.B(n_18),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_69),
.C(n_5),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_83),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_85),
.B(n_6),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_84),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_2),
.Y(n_84)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_86),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_65),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_4),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_5),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_64),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_75),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_80),
.B1(n_86),
.B2(n_6),
.Y(n_102)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_101),
.B(n_104),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_102),
.A2(n_105),
.B(n_91),
.Y(n_107)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_27),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_107),
.B(n_108),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_89),
.B(n_96),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_103),
.A2(n_97),
.B1(n_93),
.B2(n_7),
.Y(n_109)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_26),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_10),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_99),
.C(n_7),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_112),
.B(n_106),
.Y(n_115)
);

AOI321xp33_ASAP7_75t_L g117 ( 
.A1(n_115),
.A2(n_116),
.A3(n_15),
.B1(n_16),
.B2(n_21),
.C(n_22),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_114),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_117),
.B(n_28),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_113),
.C(n_30),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_29),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_33),
.C(n_34),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_35),
.C(n_37),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_38),
.Y(n_124)
);


endmodule