module fake_jpeg_2595_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_4),
.B(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_53),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_54),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_12),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_0),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_55),
.A2(n_36),
.B1(n_41),
.B2(n_43),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_61),
.B1(n_48),
.B2(n_40),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_56),
.A2(n_40),
.B1(n_43),
.B2(n_41),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

CKINVDCx6p67_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_70),
.Y(n_86)
);

AND2x6_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_15),
.Y(n_90)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_75),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_45),
.B1(n_37),
.B2(n_48),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_62),
.B1(n_5),
.B2(n_6),
.Y(n_92)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_38),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_16),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_82),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_71),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_60),
.B(n_59),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_13),
.B(n_17),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_89),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_23),
.Y(n_100)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_4),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_100),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_101),
.B(n_106),
.C(n_34),
.D(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

NOR4xp25_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_14),
.C(n_28),
.D(n_25),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_105),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_84),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_20),
.C(n_21),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_10),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_10),
.B(n_11),
.Y(n_115)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_116),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_92),
.B(n_11),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_119),
.Y(n_122)
);

A2O1A1O1Ixp25_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_95),
.B(n_96),
.C(n_104),
.D(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_123),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_120),
.B(n_113),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_124),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_113),
.C(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_128),
.A2(n_123),
.B(n_114),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_114),
.B1(n_125),
.B2(n_110),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_111),
.Y(n_131)
);


endmodule