module fake_jpeg_30362_n_144 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_12),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_0),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_69),
.Y(n_81)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_1),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_47),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_1),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_2),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_52),
.B1(n_46),
.B2(n_50),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_73),
.A2(n_79),
.B1(n_80),
.B2(n_26),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_76),
.Y(n_92)
);

CKINVDCx11_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_46),
.B1(n_50),
.B2(n_52),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_50),
.B1(n_55),
.B2(n_60),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_51),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_62),
.B(n_61),
.C(n_59),
.Y(n_83)
);

AO22x2_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_67),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_87),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_91),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_SL g89 ( 
.A(n_83),
.B(n_4),
.C(n_5),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_8),
.B(n_9),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_6),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_9),
.B1(n_45),
.B2(n_11),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_7),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_77),
.Y(n_97)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_79),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_10),
.B1(n_14),
.B2(n_15),
.Y(n_116)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_118),
.B(n_34),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_39),
.B1(n_40),
.B2(n_109),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_112),
.Y(n_119)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_23),
.B1(n_25),
.B2(n_29),
.Y(n_121)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_21),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_16),
.B(n_18),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_122),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_128),
.B1(n_130),
.B2(n_109),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_30),
.C(n_31),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_32),
.C(n_33),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_123),
.A2(n_127),
.B(n_110),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_116),
.C(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_36),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_126),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_38),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_132),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_119),
.B(n_129),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_129),
.B1(n_105),
.B2(n_119),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_137),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_134),
.B(n_125),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_106),
.Y(n_144)
);


endmodule