module real_jpeg_2100_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx2_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_1),
.A2(n_64),
.B1(n_65),
.B2(n_82),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_1),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_1),
.A2(n_49),
.B1(n_50),
.B2(n_82),
.Y(n_118)
);

BUFx4f_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_3),
.A2(n_49),
.B1(n_50),
.B2(n_58),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_3),
.A2(n_58),
.B1(n_64),
.B2(n_65),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_4),
.B(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_4),
.B(n_48),
.C(n_50),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_4),
.B(n_47),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_4),
.B(n_64),
.C(n_68),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_4),
.A2(n_38),
.B1(n_49),
.B2(n_50),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_4),
.B(n_85),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_4),
.B(n_119),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_5),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_6),
.A2(n_29),
.B1(n_49),
.B2(n_50),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_6),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_6),
.A2(n_29),
.B1(n_64),
.B2(n_65),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_9),
.Y(n_88)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_12),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_12),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_14),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_55),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_14),
.A2(n_49),
.B1(n_50),
.B2(n_55),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_14),
.A2(n_55),
.B1(n_64),
.B2(n_65),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_123),
.B1(n_202),
.B2(n_203),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_18),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_121),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_98),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_20),
.B(n_98),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.C(n_89),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_21),
.B(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_43),
.B2(n_73),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_22),
.B(n_44),
.C(n_59),
.Y(n_120)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_26),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_42)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_38),
.Y(n_39)
);

AOI32xp33_ASAP7_75t_L g76 ( 
.A1(n_27),
.A2(n_32),
.A3(n_34),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_30),
.A2(n_106),
.B(n_108),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_31),
.A2(n_32),
.B1(n_48),
.B2(n_52),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_31),
.B(n_35),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_31),
.B(n_137),
.Y(n_136)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_38),
.A2(n_114),
.B(n_152),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_39),
.Y(n_77)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_41),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_59),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_45),
.A2(n_57),
.B(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_45),
.A2(n_104),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_53),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_47),
.B(n_92),
.Y(n_104)
);

AO22x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_47)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_50),
.B1(n_67),
.B2(n_68),
.Y(n_71)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_50),
.B(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_56),
.B(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B(n_69),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_61),
.A2(n_70),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_63),
.A2(n_69),
.B(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_63),
.A2(n_131),
.B1(n_158),
.B2(n_166),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_64),
.B(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_70),
.A2(n_130),
.B(n_132),
.Y(n_129)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_70),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_72),
.B(n_119),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_74),
.B(n_89),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_79),
.B2(n_80),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_83),
.B1(n_84),
.B2(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_83),
.B(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_83),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_83),
.A2(n_84),
.B1(n_150),
.B2(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_84),
.A2(n_97),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_84),
.B(n_141),
.Y(n_152)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_87),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_85),
.A2(n_140),
.B(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.C(n_96),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_111),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_110),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_120),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_144),
.B(n_201),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_142),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_125),
.B(n_142),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.C(n_134),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_126),
.B(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_129),
.B(n_134),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_133),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_135),
.A2(n_136),
.B1(n_138),
.B2(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_138),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_196),
.B(n_200),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_186),
.B(n_195),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_168),
.B(n_185),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_161),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_161),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_153),
.B1(n_159),
.B2(n_160),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_156),
.C(n_159),
.Y(n_187)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_179),
.B(n_184),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_174),
.B(n_178),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_177),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_176),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_182),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_188),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_192),
.C(n_193),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_199),
.Y(n_200)
);


endmodule