module fake_jpeg_300_n_149 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_149);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_9),
.B(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_28),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_0),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

AND2x6_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_61),
.Y(n_68)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_1),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_40),
.B1(n_52),
.B2(n_45),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_16),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_52),
.B1(n_48),
.B2(n_41),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_70),
.A2(n_72),
.B(n_1),
.Y(n_78)
);

AO22x2_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_53),
.B1(n_18),
.B2(n_21),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_48),
.B1(n_42),
.B2(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_46),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_78),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_51),
.B(n_43),
.C(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_76),
.Y(n_92)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_3),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_2),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_83),
.Y(n_88)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_3),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_22),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_86),
.A2(n_78),
.B1(n_65),
.B2(n_71),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_91),
.B1(n_94),
.B2(n_7),
.Y(n_116)
);

AOI32xp33_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_71),
.A3(n_74),
.B1(n_81),
.B2(n_84),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_25),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_65),
.B1(n_64),
.B2(n_71),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_64),
.B1(n_4),
.B2(n_5),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_96),
.B(n_99),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_101),
.B(n_4),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_23),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_6),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_104),
.B(n_109),
.Y(n_128)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_107),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_112),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_87),
.Y(n_107)
);

AND2x6_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_15),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_110),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_5),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_102),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_116),
.B1(n_120),
.B2(n_37),
.Y(n_125)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_114),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_6),
.B(n_7),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_115),
.A2(n_118),
.B(n_119),
.Y(n_129)
);

CKINVDCx12_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_117),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_120),
.B1(n_113),
.B2(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_30),
.C(n_36),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_124),
.B(n_31),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_26),
.C(n_35),
.Y(n_124)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

BUFx12f_ASAP7_75t_SL g134 ( 
.A(n_123),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_129),
.B1(n_121),
.B2(n_126),
.Y(n_140)
);

XOR2x2_ASAP7_75t_SL g137 ( 
.A(n_127),
.B(n_108),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_132),
.B1(n_131),
.B2(n_130),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_140),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_139),
.A2(n_135),
.B1(n_136),
.B2(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_141),
.B(n_138),
.Y(n_143)
);

AOI322xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_142),
.A3(n_137),
.B1(n_131),
.B2(n_128),
.C1(n_124),
.C2(n_8),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_145),
.B(n_122),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_34),
.C(n_11),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_147),
.A2(n_10),
.B(n_11),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_10),
.Y(n_149)
);


endmodule