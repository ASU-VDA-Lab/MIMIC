module fake_jpeg_18314_n_101 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_101);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx2_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_15),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_11),
.Y(n_42)
);

INVx5_ASAP7_75t_SL g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_30),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_18),
.B1(n_12),
.B2(n_13),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_29),
.B1(n_31),
.B2(n_28),
.Y(n_51)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_26),
.B(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_15),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_13),
.B(n_10),
.Y(n_44)
);

HAxp5_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_14),
.CON(n_62),
.SN(n_62)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_11),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_33),
.B1(n_29),
.B2(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_14),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_47),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_13),
.Y(n_69)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_27),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_29),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_41),
.C(n_28),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_61),
.C(n_27),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_27),
.C(n_35),
.Y(n_61)
);

NOR4xp25_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_52),
.C(n_48),
.D(n_10),
.Y(n_64)
);

XOR2x1_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_35),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_63),
.B(n_36),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_65),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_49),
.C(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_45),
.B(n_54),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_72),
.B1(n_73),
.B2(n_33),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_25),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_60),
.C(n_62),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_76),
.C(n_77),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_37),
.C(n_18),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_37),
.C(n_18),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_29),
.B1(n_12),
.B2(n_17),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_81),
.A2(n_68),
.B1(n_17),
.B2(n_25),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_12),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_84),
.B(n_87),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_0),
.C(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_86),
.Y(n_89)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_79),
.B(n_3),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_2),
.B(n_3),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_88),
.A2(n_82),
.B1(n_17),
.B2(n_4),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_93),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_2),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_89),
.B(n_6),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_88),
.A2(n_17),
.B1(n_5),
.B2(n_6),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_97),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_8),
.B1(n_97),
.B2(n_98),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_8),
.Y(n_101)
);


endmodule