module fake_jpeg_24699_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_1),
.Y(n_13)
);

OAI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_14),
.A2(n_10),
.B1(n_9),
.B2(n_8),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_8),
.A2(n_5),
.B(n_9),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_15),
.A2(n_16),
.B(n_7),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_10),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_5),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_19),
.B(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_15),
.A2(n_7),
.B(n_16),
.C(n_17),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_18),
.B1(n_19),
.B2(n_25),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_24),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_22),
.A2(n_21),
.B1(n_25),
.B2(n_23),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_28),
.B(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_34),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_29),
.C(n_26),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_29),
.Y(n_36)
);


endmodule