module fake_ariane_1636_n_2048 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2048);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2048;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_263;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_95),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_208),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_33),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_13),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_72),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_188),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_40),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_31),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_149),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_81),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_145),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_71),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_100),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_168),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_25),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_55),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_18),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_0),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_76),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_96),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_0),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_61),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_1),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_115),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_9),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_12),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g242 ( 
.A(n_92),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_67),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_203),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_182),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_140),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_17),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_134),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_144),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_150),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_24),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_13),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_108),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_73),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_158),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_177),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_3),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_166),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_60),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_98),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_36),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_122),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_170),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_102),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_87),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_41),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_47),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_35),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_24),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_190),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_83),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_110),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_36),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_7),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_3),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_156),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_43),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_74),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_77),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_86),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_17),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_10),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_136),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_202),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_127),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_152),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_14),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_118),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_58),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_189),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_52),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_157),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_85),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_4),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_184),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_180),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_205),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_19),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_185),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_7),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_174),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_179),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_32),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_28),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_142),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_121),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_107),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_42),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_93),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_78),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_30),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_5),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_113),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_41),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_186),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_63),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_61),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_15),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_44),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_14),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_129),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_89),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_133),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_204),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_126),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_60),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_159),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_51),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_51),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_153),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_33),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_32),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_111),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_198),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_105),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_120),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_181),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_69),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_54),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_26),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_135),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_200),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_101),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_161),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_21),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_66),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_207),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_28),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_27),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_178),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_154),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_117),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_31),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_146),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_23),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_21),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_70),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_193),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_147),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_16),
.Y(n_360)
);

BUFx2_ASAP7_75t_SL g361 ( 
.A(n_114),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_80),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_103),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_187),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_23),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_88),
.Y(n_366)
);

INVxp33_ASAP7_75t_L g367 ( 
.A(n_56),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_46),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_12),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_55),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_56),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_176),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_35),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_57),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_169),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_91),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_155),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_47),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_39),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_191),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_183),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_54),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_124),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_165),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_128),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_167),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_9),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_90),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_27),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_8),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_15),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_195),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_210),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_138),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_196),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_112),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_64),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_1),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_39),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_50),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_104),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_130),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_63),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_40),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_30),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_11),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_82),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g408 ( 
.A(n_44),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_151),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_123),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_45),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_18),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_75),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_143),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_160),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_6),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_139),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_252),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_408),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_339),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_371),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_238),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_238),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_221),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_238),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_240),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_353),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_270),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_266),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_238),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_271),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_286),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_288),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_343),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_367),
.B(n_2),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_238),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_407),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_398),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_398),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_414),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_417),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_259),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_267),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_398),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_266),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_398),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_268),
.Y(n_447)
);

NOR2xp67_ASAP7_75t_L g448 ( 
.A(n_318),
.B(n_2),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_282),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_213),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_269),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_398),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_273),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_300),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_214),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_311),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_281),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_314),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_289),
.Y(n_459)
);

INVxp33_ASAP7_75t_L g460 ( 
.A(n_217),
.Y(n_460)
);

NOR2xp67_ASAP7_75t_L g461 ( 
.A(n_318),
.B(n_4),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_329),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_298),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_329),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_356),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_303),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_304),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_308),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_316),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_356),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_374),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_317),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_282),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_378),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_319),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_326),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_225),
.B(n_5),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_226),
.B(n_6),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_379),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_378),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_403),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_403),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_328),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_218),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_234),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_332),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_231),
.B(n_8),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_214),
.Y(n_488)
);

CKINVDCx14_ASAP7_75t_R g489 ( 
.A(n_285),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_234),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_355),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_360),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_228),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_282),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_227),
.B(n_230),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_416),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_285),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_285),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_295),
.Y(n_499)
);

NOR2xp67_ASAP7_75t_L g500 ( 
.A(n_227),
.B(n_10),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_212),
.B(n_11),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_302),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_236),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_230),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_247),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_247),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_302),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_251),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_305),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_305),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_295),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_251),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_295),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_313),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_257),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_257),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_313),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_365),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_365),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_333),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_333),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_383),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_237),
.B(n_16),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_485),
.B(n_232),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_422),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_485),
.B(n_490),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_422),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_423),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_426),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_490),
.B(n_233),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_423),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_501),
.B(n_223),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_425),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_425),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_430),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_430),
.Y(n_536)
);

BUFx8_ASAP7_75t_L g537 ( 
.A(n_455),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_436),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_436),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_438),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_438),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_439),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_501),
.B(n_429),
.Y(n_543)
);

NAND2xp33_ASAP7_75t_R g544 ( 
.A(n_504),
.B(n_368),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_439),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_444),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_445),
.B(n_385),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_444),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_502),
.B(n_239),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_446),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_420),
.A2(n_390),
.B1(n_275),
.B2(n_412),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_446),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_427),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_452),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_452),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_502),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_507),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_507),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_460),
.B(n_212),
.Y(n_559)
);

INVx6_ASAP7_75t_L g560 ( 
.A(n_523),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_509),
.B(n_385),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_509),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_510),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_510),
.Y(n_564)
);

OA21x2_ASAP7_75t_L g565 ( 
.A1(n_514),
.A2(n_260),
.B(n_258),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_514),
.B(n_262),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_517),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_419),
.B(n_383),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_517),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_455),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_520),
.B(n_248),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_520),
.B(n_276),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_521),
.Y(n_573)
);

INVxp33_ASAP7_75t_SL g574 ( 
.A(n_442),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_521),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_522),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_522),
.Y(n_577)
);

AND2x6_ASAP7_75t_L g578 ( 
.A(n_477),
.B(n_223),
.Y(n_578)
);

OA21x2_ASAP7_75t_L g579 ( 
.A1(n_478),
.A2(n_487),
.B(n_283),
.Y(n_579)
);

AND2x6_ASAP7_75t_L g580 ( 
.A(n_450),
.B(n_223),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_462),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_462),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_484),
.B(n_503),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_464),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_464),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_493),
.B(n_278),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_465),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_465),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_470),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_470),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_474),
.B(n_248),
.Y(n_591)
);

OAI21x1_ASAP7_75t_L g592 ( 
.A1(n_523),
.A2(n_315),
.B(n_293),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_474),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_480),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_480),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_481),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_481),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_482),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_482),
.B(n_321),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_435),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_443),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_447),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_448),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_518),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_451),
.B(n_211),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_518),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_461),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_488),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_600),
.B(n_489),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_601),
.B(n_453),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_562),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_562),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_590),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_536),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_562),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_601),
.B(n_457),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_600),
.B(n_459),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_536),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_532),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_560),
.B(n_500),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_600),
.B(n_463),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_543),
.B(n_466),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_562),
.Y(n_623)
);

AND2x6_ASAP7_75t_L g624 ( 
.A(n_601),
.B(n_363),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_L g625 ( 
.A(n_532),
.B(n_242),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_601),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_536),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_601),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_601),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_590),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_605),
.B(n_467),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_536),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_536),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_562),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_560),
.B(n_449),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_543),
.B(n_468),
.Y(n_636)
);

AO22x2_ASAP7_75t_L g637 ( 
.A1(n_583),
.A2(n_370),
.B1(n_312),
.B2(n_229),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_601),
.B(n_469),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_545),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_562),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_559),
.Y(n_641)
);

BUFx6f_ASAP7_75t_SL g642 ( 
.A(n_601),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_545),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_545),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_545),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_562),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_543),
.B(n_472),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_562),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_569),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_605),
.B(n_475),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_602),
.B(n_583),
.Y(n_651)
);

INVxp67_ASAP7_75t_SL g652 ( 
.A(n_524),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_545),
.Y(n_653)
);

AND2x6_ASAP7_75t_L g654 ( 
.A(n_602),
.B(n_363),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_543),
.B(n_476),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_550),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_528),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_550),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_550),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_550),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_602),
.B(n_583),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_559),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_602),
.B(n_483),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_543),
.B(n_547),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_556),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_556),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_SL g667 ( 
.A(n_574),
.B(n_497),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_558),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_547),
.B(n_495),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_547),
.B(n_486),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_558),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_547),
.B(n_491),
.Y(n_672)
);

AND2x4_ASAP7_75t_SL g673 ( 
.A(n_602),
.B(n_498),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_568),
.B(n_492),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_550),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_583),
.B(n_323),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_559),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_SL g678 ( 
.A(n_544),
.B(n_499),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_525),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_529),
.Y(n_680)
);

BUFx4f_ASAP7_75t_L g681 ( 
.A(n_532),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_563),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_583),
.B(n_505),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_574),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_532),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_592),
.B(n_324),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_592),
.B(n_606),
.Y(n_687)
);

CKINVDCx6p67_ASAP7_75t_R g688 ( 
.A(n_529),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_532),
.B(n_506),
.Y(n_689)
);

OR2x6_ASAP7_75t_L g690 ( 
.A(n_560),
.B(n_361),
.Y(n_690)
);

BUFx4f_ASAP7_75t_L g691 ( 
.A(n_532),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_525),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_591),
.B(n_571),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_568),
.B(n_508),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_525),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_560),
.B(n_512),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_563),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_570),
.B(n_473),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_560),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_569),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_560),
.B(n_241),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_532),
.B(n_515),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_571),
.B(n_261),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_SL g704 ( 
.A1(n_537),
.A2(n_511),
.B1(n_513),
.B2(n_418),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_567),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_525),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_532),
.B(n_516),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_533),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_533),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_532),
.B(n_519),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_528),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_567),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_573),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_533),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_544),
.A2(n_494),
.B1(n_368),
.B2(n_373),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_539),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_537),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_570),
.B(n_421),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_573),
.Y(n_719)
);

BUFx10_ASAP7_75t_L g720 ( 
.A(n_532),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_539),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_529),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_575),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_604),
.B(n_432),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_606),
.B(n_382),
.C(n_373),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_569),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_539),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_575),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_592),
.B(n_325),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_569),
.Y(n_730)
);

OAI21xp33_ASAP7_75t_SL g731 ( 
.A1(n_606),
.A2(n_277),
.B(n_274),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_537),
.Y(n_732)
);

BUFx8_ASAP7_75t_SL g733 ( 
.A(n_553),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_569),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_577),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_R g736 ( 
.A(n_553),
.B(n_434),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_577),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_576),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_546),
.Y(n_739)
);

INVx5_ASAP7_75t_L g740 ( 
.A(n_580),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_606),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_546),
.Y(n_742)
);

AND2x6_ASAP7_75t_L g743 ( 
.A(n_561),
.B(n_571),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_546),
.Y(n_744)
);

AND2x6_ASAP7_75t_L g745 ( 
.A(n_561),
.B(n_366),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_582),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_591),
.B(n_287),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_576),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_528),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_604),
.B(n_608),
.C(n_537),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_528),
.Y(n_751)
);

NAND2xp33_ASAP7_75t_L g752 ( 
.A(n_578),
.B(n_242),
.Y(n_752)
);

INVx4_ASAP7_75t_SL g753 ( 
.A(n_580),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_L g754 ( 
.A1(n_551),
.A2(n_391),
.B1(n_397),
.B2(n_399),
.Y(n_754)
);

BUFx10_ASAP7_75t_L g755 ( 
.A(n_561),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_579),
.A2(n_291),
.B1(n_349),
.B2(n_348),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_579),
.A2(n_411),
.B1(n_387),
.B2(n_345),
.Y(n_757)
);

INVx5_ASAP7_75t_L g758 ( 
.A(n_580),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_738),
.Y(n_759)
);

INVx8_ASAP7_75t_L g760 ( 
.A(n_743),
.Y(n_760)
);

INVx8_ASAP7_75t_L g761 ( 
.A(n_743),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_617),
.B(n_604),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_621),
.B(n_652),
.Y(n_763)
);

O2A1O1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_664),
.A2(n_586),
.B(n_585),
.C(n_608),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_741),
.B(n_608),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_696),
.B(n_537),
.Y(n_766)
);

OR2x6_ASAP7_75t_L g767 ( 
.A(n_635),
.B(n_553),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_L g768 ( 
.A1(n_690),
.A2(n_551),
.B1(n_586),
.B2(n_530),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_741),
.B(n_579),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_651),
.B(n_579),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_651),
.A2(n_579),
.B1(n_578),
.B2(n_561),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_661),
.B(n_561),
.Y(n_772)
);

NAND2xp33_ASAP7_75t_L g773 ( 
.A(n_654),
.B(n_578),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_661),
.B(n_591),
.Y(n_774)
);

OAI221xp5_ASAP7_75t_L g775 ( 
.A1(n_641),
.A2(n_369),
.B1(n_405),
.B2(n_294),
.C(n_320),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_738),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_743),
.A2(n_578),
.B1(n_580),
.B2(n_441),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_649),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_701),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_641),
.B(n_585),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_743),
.A2(n_578),
.B1(n_580),
.B2(n_437),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_738),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_609),
.B(n_603),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_662),
.B(n_585),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_662),
.B(n_585),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_685),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_680),
.B(n_440),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_SL g788 ( 
.A1(n_704),
.A2(n_454),
.B1(n_456),
.B2(n_458),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_637),
.A2(n_578),
.B1(n_565),
.B2(n_580),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_708),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_708),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_677),
.B(n_585),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_685),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_722),
.B(n_718),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_649),
.Y(n_795)
);

INVx6_ASAP7_75t_L g796 ( 
.A(n_755),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_677),
.B(n_603),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_SL g798 ( 
.A(n_717),
.B(n_424),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_698),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_649),
.Y(n_800)
);

NOR2xp67_ASAP7_75t_L g801 ( 
.A(n_684),
.B(n_750),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_700),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_709),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_631),
.B(n_211),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_743),
.A2(n_578),
.B1(n_580),
.B2(n_215),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_700),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_683),
.B(n_607),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_693),
.B(n_607),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_700),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_650),
.B(n_215),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_743),
.A2(n_578),
.B1(n_580),
.B2(n_216),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_701),
.Y(n_812)
);

OR2x6_ASAP7_75t_L g813 ( 
.A(n_635),
.B(n_599),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_622),
.B(n_389),
.C(n_382),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_709),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_726),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_693),
.B(n_578),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_669),
.B(n_578),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_636),
.B(n_647),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_670),
.B(n_219),
.Y(n_820)
);

BUFx8_ASAP7_75t_L g821 ( 
.A(n_724),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_699),
.A2(n_404),
.B1(n_400),
.B2(n_399),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_669),
.B(n_582),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_669),
.B(n_584),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_714),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_655),
.B(n_524),
.Y(n_826)
);

INVxp67_ASAP7_75t_L g827 ( 
.A(n_736),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_676),
.B(n_584),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_619),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_676),
.B(n_587),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_699),
.B(n_587),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_673),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_726),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_672),
.B(n_530),
.Y(n_834)
);

NAND2xp33_ASAP7_75t_L g835 ( 
.A(n_654),
.B(n_580),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_SL g836 ( 
.A(n_717),
.B(n_428),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_635),
.Y(n_837)
);

NOR2xp67_ASAP7_75t_SL g838 ( 
.A(n_619),
.B(n_389),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_681),
.B(n_691),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_694),
.B(n_549),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_726),
.B(n_593),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_716),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_619),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_681),
.B(n_219),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_730),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_674),
.B(n_549),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_730),
.B(n_593),
.Y(n_847)
);

BUFx6f_ASAP7_75t_SL g848 ( 
.A(n_703),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_681),
.B(n_222),
.Y(n_849)
);

INVx4_ASAP7_75t_L g850 ( 
.A(n_691),
.Y(n_850)
);

NAND2x1p5_ASAP7_75t_L g851 ( 
.A(n_691),
.B(n_565),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_730),
.B(n_598),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_665),
.B(n_598),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_613),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_663),
.B(n_755),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_666),
.B(n_557),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_668),
.B(n_557),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_663),
.B(n_566),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_620),
.A2(n_580),
.B1(n_375),
.B2(n_372),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_671),
.B(n_557),
.Y(n_860)
);

NOR3xp33_ASAP7_75t_L g861 ( 
.A(n_725),
.B(n_397),
.C(n_391),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_SL g862 ( 
.A(n_732),
.B(n_431),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_716),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_SL g864 ( 
.A1(n_637),
.A2(n_433),
.B1(n_496),
.B2(n_479),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_755),
.B(n_222),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_635),
.B(n_566),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_682),
.B(n_564),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_610),
.B(n_572),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_697),
.B(n_564),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_715),
.B(n_224),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_SL g871 ( 
.A(n_732),
.B(n_471),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_701),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_687),
.A2(n_572),
.B(n_576),
.C(n_534),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_720),
.B(n_224),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_610),
.B(n_599),
.Y(n_875)
);

NAND2xp33_ASAP7_75t_L g876 ( 
.A(n_654),
.B(n_235),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_705),
.B(n_564),
.Y(n_877)
);

INVx8_ASAP7_75t_L g878 ( 
.A(n_745),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_712),
.B(n_576),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_721),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_713),
.B(n_581),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_688),
.B(n_581),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_688),
.B(n_581),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_720),
.B(n_626),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_701),
.Y(n_885)
);

NOR2x1p5_ASAP7_75t_L g886 ( 
.A(n_684),
.B(n_400),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_630),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_719),
.B(n_588),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_723),
.B(n_588),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_728),
.B(n_588),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_721),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_616),
.B(n_526),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_690),
.A2(n_404),
.B1(n_340),
.B2(n_331),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_735),
.B(n_589),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_720),
.B(n_235),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_626),
.B(n_243),
.Y(n_896)
);

NOR2xp67_ASAP7_75t_L g897 ( 
.A(n_616),
.B(n_526),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_638),
.B(n_589),
.Y(n_898)
);

NOR2x1p5_ASAP7_75t_SL g899 ( 
.A(n_614),
.B(n_242),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_737),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_727),
.Y(n_901)
);

AND2x6_ASAP7_75t_L g902 ( 
.A(n_753),
.B(n_366),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_746),
.B(n_589),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_637),
.A2(n_757),
.B1(n_756),
.B2(n_625),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_734),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_727),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_626),
.B(n_243),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_638),
.B(n_594),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_734),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_620),
.B(n_594),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_620),
.B(n_338),
.Y(n_911)
);

INVxp67_ASAP7_75t_SL g912 ( 
.A(n_625),
.Y(n_912)
);

NAND2xp33_ASAP7_75t_L g913 ( 
.A(n_654),
.B(n_244),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_618),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_620),
.B(n_594),
.Y(n_915)
);

O2A1O1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_687),
.A2(n_406),
.B(n_597),
.C(n_595),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_673),
.Y(n_917)
);

AND2x2_ASAP7_75t_SL g918 ( 
.A(n_752),
.B(n_565),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_747),
.B(n_595),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_747),
.B(n_595),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_739),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_689),
.B(n_244),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_702),
.B(n_245),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_745),
.B(n_596),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_745),
.B(n_596),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_618),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_760),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_787),
.B(n_667),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_846),
.B(n_703),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_763),
.B(n_707),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_900),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_846),
.B(n_703),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_840),
.B(n_826),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_840),
.B(n_690),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_760),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_819),
.B(n_678),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_826),
.B(n_690),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_819),
.B(n_678),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_SL g939 ( 
.A(n_798),
.B(n_733),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_834),
.B(n_745),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_794),
.Y(n_941)
);

INVx4_ASAP7_75t_L g942 ( 
.A(n_760),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_799),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_827),
.B(n_733),
.Y(n_944)
);

O2A1O1Ixp33_ASAP7_75t_SL g945 ( 
.A1(n_817),
.A2(n_873),
.B(n_710),
.C(n_855),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_834),
.B(n_745),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_762),
.B(n_745),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_SL g948 ( 
.A1(n_896),
.A2(n_907),
.B(n_849),
.C(n_844),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_912),
.A2(n_629),
.B(n_628),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_922),
.A2(n_729),
.B(n_686),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_821),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_837),
.B(n_740),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_759),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_837),
.B(n_740),
.Y(n_954)
);

INVxp67_ASAP7_75t_R g955 ( 
.A(n_882),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_821),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_858),
.B(n_654),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_866),
.B(n_740),
.Y(n_958)
);

NOR3xp33_ASAP7_75t_L g959 ( 
.A(n_804),
.B(n_754),
.C(n_731),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_858),
.A2(n_658),
.B(n_656),
.C(n_627),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_770),
.A2(n_729),
.B(n_686),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_866),
.B(n_740),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_807),
.B(n_654),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_914),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_926),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_807),
.B(n_748),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_769),
.A2(n_752),
.B(n_632),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_783),
.B(n_748),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_841),
.A2(n_632),
.B(n_627),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_783),
.B(n_633),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_847),
.A2(n_639),
.B(n_633),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_827),
.B(n_639),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_852),
.A2(n_644),
.B(n_643),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_765),
.B(n_643),
.Y(n_974)
);

NOR3xp33_ASAP7_75t_L g975 ( 
.A(n_810),
.B(n_645),
.C(n_644),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_780),
.A2(n_653),
.B(n_645),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_784),
.A2(n_656),
.B(n_653),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_785),
.A2(n_659),
.B(n_658),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_792),
.A2(n_892),
.B(n_919),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_767),
.B(n_596),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_923),
.A2(n_660),
.B(n_659),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_767),
.B(n_597),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_892),
.A2(n_675),
.B(n_660),
.Y(n_983)
);

AOI22x1_ASAP7_75t_L g984 ( 
.A1(n_778),
.A2(n_675),
.B1(n_640),
.B2(n_634),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_911),
.B(n_739),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_920),
.A2(n_623),
.B(n_612),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_767),
.B(n_597),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_868),
.A2(n_623),
.B(n_612),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_836),
.B(n_642),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_808),
.A2(n_612),
.B(n_634),
.C(n_640),
.Y(n_990)
);

NAND2x1p5_ASAP7_75t_L g991 ( 
.A(n_786),
.B(n_740),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_761),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_868),
.B(n_742),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_773),
.A2(n_634),
.B(n_623),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_875),
.B(n_768),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_879),
.A2(n_640),
.B(n_642),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_831),
.A2(n_642),
.B(n_615),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_875),
.B(n_742),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_768),
.B(n_744),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_774),
.B(n_744),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_883),
.B(n_565),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_793),
.B(n_679),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_771),
.A2(n_695),
.B(n_692),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_761),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_SL g1005 ( 
.A1(n_865),
.A2(n_706),
.B(n_695),
.C(n_692),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_761),
.Y(n_1006)
);

NAND2x1_ASAP7_75t_L g1007 ( 
.A(n_850),
.B(n_796),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_823),
.B(n_706),
.Y(n_1008)
);

AOI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_893),
.A2(n_565),
.B(n_611),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_786),
.Y(n_1010)
);

NOR2xp67_ASAP7_75t_L g1011 ( 
.A(n_832),
.B(n_527),
.Y(n_1011)
);

O2A1O1Ixp5_ASAP7_75t_L g1012 ( 
.A1(n_838),
.A2(n_541),
.B(n_527),
.C(n_531),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_856),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_857),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_824),
.B(n_624),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_860),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_916),
.A2(n_624),
.B(n_758),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_898),
.A2(n_624),
.B(n_758),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_917),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_839),
.A2(n_615),
.B(n_611),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_910),
.B(n_624),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_898),
.A2(n_624),
.B(n_758),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_876),
.A2(n_615),
.B(n_611),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_913),
.A2(n_615),
.B(n_611),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_867),
.A2(n_648),
.B(n_646),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_869),
.Y(n_1026)
);

NOR2xp67_ASAP7_75t_L g1027 ( 
.A(n_801),
.B(n_531),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_862),
.B(n_534),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_871),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_764),
.A2(n_538),
.B(n_535),
.C(n_540),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_813),
.A2(n_624),
.B1(n_646),
.B2(n_648),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_877),
.A2(n_648),
.B(n_646),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_870),
.B(n_646),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_910),
.A2(n_381),
.B(n_377),
.C(n_376),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_881),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_779),
.B(n_758),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_888),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_779),
.B(n_753),
.Y(n_1038)
);

AND2x6_ASAP7_75t_L g1039 ( 
.A(n_829),
.B(n_753),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_889),
.A2(n_648),
.B(n_751),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_812),
.B(n_758),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_890),
.A2(n_751),
.B(n_749),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_915),
.B(n_657),
.Y(n_1043)
);

INVx5_ASAP7_75t_L g1044 ( 
.A(n_878),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_915),
.A2(n_359),
.B(n_347),
.C(n_401),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_772),
.B(n_657),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_797),
.B(n_657),
.Y(n_1047)
);

BUFx4f_ASAP7_75t_L g1048 ( 
.A(n_813),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_894),
.A2(n_751),
.B(n_749),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_903),
.A2(n_751),
.B(n_749),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_812),
.A2(n_375),
.B1(n_246),
.B2(n_249),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_776),
.A2(n_749),
.B(n_711),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_854),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_788),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_796),
.A2(n_711),
.B1(n_657),
.B2(n_327),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_782),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_SL g1057 ( 
.A1(n_795),
.A2(n_330),
.B(n_336),
.C(n_337),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_796),
.A2(n_711),
.B1(n_402),
.B2(n_256),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_872),
.B(n_711),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_886),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_872),
.B(n_245),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_904),
.B(n_897),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_790),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_878),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_820),
.B(n_362),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_885),
.B(n_541),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_814),
.B(n_542),
.Y(n_1067)
);

CKINVDCx10_ASAP7_75t_R g1068 ( 
.A(n_848),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_885),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_800),
.A2(n_253),
.B(n_413),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_814),
.B(n_548),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_850),
.B(n_548),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_828),
.B(n_830),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_853),
.B(n_552),
.Y(n_1074)
);

NAND2x1_ASAP7_75t_L g1075 ( 
.A(n_829),
.B(n_552),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_848),
.B(n_246),
.Y(n_1076)
);

NOR2x1p5_ASAP7_75t_L g1077 ( 
.A(n_818),
.B(n_249),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_802),
.A2(n_554),
.B(n_555),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_806),
.A2(n_554),
.B(n_555),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_905),
.B(n_250),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_905),
.B(n_250),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_809),
.A2(n_528),
.B(n_253),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_777),
.B(n_254),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_816),
.A2(n_528),
.B(n_254),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_833),
.B(n_255),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_789),
.A2(n_415),
.B1(n_392),
.B2(n_413),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_843),
.A2(n_255),
.B1(n_310),
.B2(n_410),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_887),
.A2(n_415),
.B(n_20),
.C(n_22),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_861),
.A2(n_310),
.B1(n_410),
.B2(n_409),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_845),
.B(n_256),
.Y(n_1090)
);

INVx4_ASAP7_75t_L g1091 ( 
.A(n_878),
.Y(n_1091)
);

CKINVDCx10_ASAP7_75t_R g1092 ( 
.A(n_864),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_908),
.A2(n_528),
.B(n_409),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_909),
.B(n_372),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_835),
.A2(n_918),
.B(n_884),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_766),
.B(n_380),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_918),
.A2(n_380),
.B(n_396),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_805),
.A2(n_384),
.B(n_396),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_R g1099 ( 
.A(n_902),
.B(n_384),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_811),
.A2(n_386),
.B(n_395),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_843),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_822),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_851),
.A2(n_386),
.B(n_395),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_924),
.A2(n_925),
.B(n_874),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_791),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_803),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_775),
.B(n_388),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_815),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_859),
.B(n_825),
.Y(n_1109)
);

AOI21x1_ASAP7_75t_L g1110 ( 
.A1(n_895),
.A2(n_528),
.B(n_242),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_842),
.A2(n_921),
.B(n_906),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_936),
.B(n_781),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_933),
.A2(n_861),
.B(n_899),
.C(n_789),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_927),
.Y(n_1114)
);

AO21x2_ASAP7_75t_L g1115 ( 
.A1(n_1009),
.A2(n_901),
.B(n_891),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_928),
.B(n_864),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_995),
.B(n_863),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_938),
.B(n_851),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_931),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_927),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_929),
.B(n_880),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_932),
.A2(n_19),
.B(n_20),
.C(n_22),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_927),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_937),
.B(n_388),
.Y(n_1124)
);

NOR3xp33_ASAP7_75t_L g1125 ( 
.A(n_1088),
.B(n_392),
.C(n_393),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1053),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1013),
.B(n_902),
.Y(n_1127)
);

OA21x2_ASAP7_75t_L g1128 ( 
.A1(n_1003),
.A2(n_393),
.B(n_394),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_979),
.A2(n_309),
.B(n_264),
.Y(n_1129)
);

OAI22x1_ASAP7_75t_L g1130 ( 
.A1(n_1054),
.A2(n_394),
.B1(n_322),
.B2(n_364),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1063),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_SL g1132 ( 
.A1(n_990),
.A2(n_25),
.B(n_26),
.C(n_29),
.Y(n_1132)
);

AO22x1_ASAP7_75t_L g1133 ( 
.A1(n_944),
.A2(n_956),
.B1(n_951),
.B2(n_1107),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1006),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_941),
.B(n_29),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1102),
.B(n_902),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_982),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_1038),
.B(n_902),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_942),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_934),
.A2(n_940),
.B(n_946),
.C(n_959),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_1069),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_1006),
.Y(n_1142)
);

INVx4_ASAP7_75t_L g1143 ( 
.A(n_1006),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1065),
.A2(n_306),
.B(n_358),
.C(n_357),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_979),
.A2(n_301),
.B(n_354),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_970),
.A2(n_299),
.B(n_352),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1106),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_1019),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1097),
.A2(n_296),
.B(n_351),
.C(n_350),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1067),
.A2(n_1071),
.B(n_1090),
.C(n_1085),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_963),
.A2(n_292),
.B(n_346),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_966),
.A2(n_290),
.B(n_344),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1038),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_943),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_968),
.A2(n_284),
.B(n_342),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1014),
.B(n_902),
.Y(n_1156)
);

INVx5_ASAP7_75t_L g1157 ( 
.A(n_1039),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_955),
.B(n_34),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_957),
.A2(n_341),
.B(n_335),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_987),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_930),
.A2(n_334),
.B(n_307),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1016),
.B(n_34),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1029),
.B(n_297),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_964),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1062),
.A2(n_280),
.B1(n_279),
.B2(n_272),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_980),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1026),
.B(n_242),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1074),
.A2(n_263),
.B1(n_265),
.B2(n_220),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_SL g1169 ( 
.A1(n_988),
.A2(n_37),
.B(n_38),
.C(n_42),
.Y(n_1169)
);

OAI22x1_ASAP7_75t_L g1170 ( 
.A1(n_1089),
.A2(n_37),
.B1(n_38),
.B2(n_43),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1035),
.B(n_242),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1037),
.B(n_1073),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_939),
.A2(n_242),
.B1(n_220),
.B2(n_48),
.Y(n_1173)
);

BUFx12f_ASAP7_75t_L g1174 ( 
.A(n_1060),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_945),
.A2(n_220),
.B(n_109),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1076),
.B(n_942),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_993),
.B(n_998),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_972),
.B(n_45),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_965),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1001),
.B(n_46),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_1028),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1064),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1048),
.B(n_220),
.Y(n_1183)
);

O2A1O1Ixp5_ASAP7_75t_L g1184 ( 
.A1(n_1103),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_994),
.A2(n_119),
.B(n_192),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1066),
.B(n_49),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1000),
.B(n_52),
.Y(n_1187)
);

OR2x6_ASAP7_75t_L g1188 ( 
.A(n_1041),
.B(n_53),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1041),
.B(n_53),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1048),
.B(n_57),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1105),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1108),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_1044),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_SL g1194 ( 
.A1(n_1092),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1066),
.B(n_59),
.Y(n_1195)
);

INVx3_ASAP7_75t_SL g1196 ( 
.A(n_1068),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_953),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_967),
.A2(n_132),
.B(n_175),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1094),
.A2(n_1098),
.B(n_1100),
.C(n_948),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_960),
.A2(n_62),
.B(n_65),
.C(n_68),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1056),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1010),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_947),
.A2(n_65),
.B(n_79),
.C(n_84),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_967),
.A2(n_94),
.B(n_97),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1010),
.Y(n_1205)
);

INVxp67_ASAP7_75t_L g1206 ( 
.A(n_1061),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1008),
.Y(n_1207)
);

INVx3_ASAP7_75t_SL g1208 ( 
.A(n_1059),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_SL g1209 ( 
.A(n_1072),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1087),
.A2(n_1081),
.B(n_1080),
.C(n_1034),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1051),
.B(n_209),
.Y(n_1211)
);

O2A1O1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1045),
.A2(n_99),
.B(n_106),
.C(n_116),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_989),
.B(n_125),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1044),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1096),
.B(n_131),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_974),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_950),
.A2(n_137),
.B(n_141),
.Y(n_1217)
);

INVx4_ASAP7_75t_L g1218 ( 
.A(n_1044),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1007),
.Y(n_1219)
);

BUFx4f_ASAP7_75t_L g1220 ( 
.A(n_935),
.Y(n_1220)
);

AND3x1_ASAP7_75t_SL g1221 ( 
.A(n_1077),
.B(n_173),
.C(n_162),
.Y(n_1221)
);

BUFx12f_ASAP7_75t_L g1222 ( 
.A(n_1064),
.Y(n_1222)
);

NOR2xp67_ASAP7_75t_L g1223 ( 
.A(n_985),
.B(n_148),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1011),
.B(n_163),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1020),
.A2(n_164),
.B(n_171),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_935),
.B(n_172),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1044),
.B(n_1091),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_992),
.B(n_1004),
.Y(n_1228)
);

AO21x1_ASAP7_75t_L g1229 ( 
.A1(n_999),
.A2(n_1095),
.B(n_1104),
.Y(n_1229)
);

NOR3xp33_ASAP7_75t_SL g1230 ( 
.A(n_1070),
.B(n_1058),
.C(n_1082),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_1043),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_992),
.B(n_1004),
.Y(n_1232)
);

AOI221xp5_ASAP7_75t_L g1233 ( 
.A1(n_1086),
.A2(n_1057),
.B1(n_1083),
.B2(n_1079),
.C(n_983),
.Y(n_1233)
);

NAND2xp33_ASAP7_75t_L g1234 ( 
.A(n_1039),
.B(n_1101),
.Y(n_1234)
);

AND2x6_ASAP7_75t_SL g1235 ( 
.A(n_1033),
.B(n_1072),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_1099),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1002),
.B(n_1047),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1036),
.A2(n_954),
.B1(n_952),
.B2(n_1109),
.Y(n_1238)
);

INVx3_ASAP7_75t_SL g1239 ( 
.A(n_1091),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1039),
.Y(n_1240)
);

INVx6_ASAP7_75t_L g1241 ( 
.A(n_1039),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1027),
.B(n_1046),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1078),
.Y(n_1243)
);

HAxp5_ASAP7_75t_L g1244 ( 
.A(n_975),
.B(n_1082),
.CON(n_1244),
.SN(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1030),
.A2(n_1005),
.B(n_983),
.C(n_1084),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1101),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1039),
.B(n_1095),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_976),
.B(n_977),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_958),
.A2(n_962),
.B1(n_1055),
.B2(n_1031),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1078),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1025),
.A2(n_1042),
.B(n_1040),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_991),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1021),
.B(n_991),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1084),
.A2(n_1093),
.B(n_981),
.C(n_978),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_976),
.B(n_978),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_977),
.B(n_969),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_969),
.B(n_971),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_971),
.B(n_973),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_973),
.B(n_986),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_986),
.B(n_1111),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1111),
.B(n_961),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1015),
.B(n_1075),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1093),
.B(n_1052),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1018),
.A2(n_1022),
.B1(n_949),
.B2(n_1017),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_984),
.Y(n_1265)
);

NAND2x1p5_ASAP7_75t_L g1266 ( 
.A(n_997),
.B(n_1032),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1012),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1049),
.B(n_1050),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1251),
.A2(n_996),
.B(n_1110),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1154),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1141),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1209),
.B(n_1023),
.Y(n_1272)
);

AOI21xp33_ASAP7_75t_L g1273 ( 
.A1(n_1199),
.A2(n_1112),
.B(n_1178),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1234),
.A2(n_1024),
.B(n_1177),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1148),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1177),
.A2(n_1258),
.B(n_1257),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1174),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1116),
.A2(n_1194),
.B1(n_1211),
.B2(n_1189),
.Y(n_1278)
);

AOI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1268),
.A2(n_1258),
.B(n_1257),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1256),
.A2(n_1255),
.B(n_1248),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1178),
.A2(n_1188),
.B1(n_1172),
.B2(n_1189),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1166),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1188),
.A2(n_1162),
.B1(n_1180),
.B2(n_1149),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1209),
.A2(n_1206),
.B1(n_1163),
.B2(n_1188),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1181),
.B(n_1207),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_SL g1286 ( 
.A1(n_1169),
.A2(n_1132),
.B(n_1113),
.C(n_1226),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1259),
.A2(n_1247),
.B(n_1260),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1181),
.B(n_1216),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1247),
.A2(n_1237),
.B(n_1264),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1231),
.B(n_1137),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1231),
.B(n_1160),
.Y(n_1291)
);

O2A1O1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1150),
.A2(n_1144),
.B(n_1125),
.C(n_1122),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1126),
.Y(n_1293)
);

O2A1O1Ixp33_ASAP7_75t_SL g1294 ( 
.A1(n_1228),
.A2(n_1232),
.B(n_1210),
.C(n_1187),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1175),
.A2(n_1261),
.B(n_1254),
.Y(n_1295)
);

BUFx8_ASAP7_75t_L g1296 ( 
.A(n_1158),
.Y(n_1296)
);

NAND2xp33_ASAP7_75t_SL g1297 ( 
.A(n_1239),
.B(n_1240),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1261),
.A2(n_1245),
.B(n_1204),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1196),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1240),
.B(n_1157),
.Y(n_1300)
);

AOI221x1_ASAP7_75t_L g1301 ( 
.A1(n_1170),
.A2(n_1203),
.B1(n_1168),
.B2(n_1198),
.C(n_1267),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1243),
.A2(n_1250),
.B(n_1225),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1186),
.B(n_1195),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1265),
.A2(n_1118),
.B(n_1117),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_1222),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1190),
.A2(n_1133),
.B1(n_1130),
.B2(n_1215),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1117),
.A2(n_1185),
.B(n_1233),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1180),
.A2(n_1187),
.B1(n_1173),
.B2(n_1168),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1131),
.Y(n_1309)
);

NAND2x1p5_ASAP7_75t_L g1310 ( 
.A(n_1157),
.B(n_1240),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1153),
.Y(n_1311)
);

AOI221xp5_ASAP7_75t_SL g1312 ( 
.A1(n_1200),
.A2(n_1129),
.B1(n_1145),
.B2(n_1155),
.C(n_1152),
.Y(n_1312)
);

NOR3xp33_ASAP7_75t_L g1313 ( 
.A(n_1184),
.B(n_1124),
.C(n_1176),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1262),
.A2(n_1217),
.B(n_1157),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1153),
.Y(n_1315)
);

AO21x2_ASAP7_75t_L g1316 ( 
.A1(n_1115),
.A2(n_1136),
.B(n_1167),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1164),
.B(n_1179),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1253),
.A2(n_1127),
.B(n_1121),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1171),
.A2(n_1156),
.B(n_1249),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1192),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1135),
.A2(n_1230),
.B1(n_1238),
.B2(n_1241),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_SL g1322 ( 
.A1(n_1213),
.A2(n_1224),
.B(n_1227),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1171),
.A2(n_1252),
.B(n_1212),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1151),
.A2(n_1115),
.B(n_1159),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1114),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1220),
.A2(n_1146),
.B(n_1128),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1128),
.A2(n_1242),
.B(n_1223),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1208),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1165),
.A2(n_1161),
.B(n_1205),
.C(n_1202),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1220),
.A2(n_1246),
.B(n_1183),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1246),
.A2(n_1182),
.B(n_1139),
.Y(n_1331)
);

AOI221x1_ASAP7_75t_L g1332 ( 
.A1(n_1197),
.A2(n_1201),
.B1(n_1244),
.B2(n_1147),
.C(n_1221),
.Y(n_1332)
);

AO21x1_ASAP7_75t_L g1333 ( 
.A1(n_1218),
.A2(n_1227),
.B(n_1138),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1114),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1218),
.A2(n_1143),
.A3(n_1235),
.B(n_1241),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1114),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1139),
.A2(n_1182),
.B1(n_1138),
.B2(n_1236),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1120),
.Y(n_1338)
);

AOI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1219),
.A2(n_1193),
.B(n_1214),
.Y(n_1339)
);

AO31x2_ASAP7_75t_L g1340 ( 
.A1(n_1143),
.A2(n_1193),
.A3(n_1214),
.B(n_1134),
.Y(n_1340)
);

O2A1O1Ixp33_ASAP7_75t_SL g1341 ( 
.A1(n_1193),
.A2(n_1214),
.B(n_1123),
.C(n_1134),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1120),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1120),
.B(n_1142),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1142),
.B(n_1123),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1142),
.A2(n_1123),
.B(n_1134),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1140),
.A2(n_933),
.B(n_995),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1241),
.Y(n_1347)
);

O2A1O1Ixp5_ASAP7_75t_L g1348 ( 
.A1(n_1229),
.A2(n_616),
.B(n_638),
.C(n_610),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1137),
.B(n_928),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1119),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1251),
.A2(n_1266),
.B(n_1258),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1148),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1234),
.A2(n_933),
.B(n_934),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1154),
.B(n_684),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1251),
.A2(n_1266),
.B(n_1258),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1251),
.A2(n_1266),
.B(n_1258),
.Y(n_1356)
);

NAND3xp33_ASAP7_75t_L g1357 ( 
.A(n_1199),
.B(n_933),
.C(n_936),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1194),
.A2(n_667),
.B1(n_680),
.B2(n_936),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1154),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1251),
.A2(n_1266),
.B(n_1258),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1234),
.A2(n_933),
.B(n_934),
.Y(n_1361)
);

OA22x2_ASAP7_75t_L g1362 ( 
.A1(n_1194),
.A2(n_767),
.B1(n_788),
.B2(n_1188),
.Y(n_1362)
);

BUFx12f_ASAP7_75t_L g1363 ( 
.A(n_1174),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1251),
.A2(n_1266),
.B(n_1258),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1154),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1137),
.B(n_928),
.Y(n_1366)
);

CKINVDCx8_ASAP7_75t_R g1367 ( 
.A(n_1235),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1194),
.A2(n_667),
.B1(n_680),
.B2(n_936),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_1141),
.Y(n_1369)
);

NOR3xp33_ASAP7_75t_L g1370 ( 
.A(n_1194),
.B(n_933),
.C(n_684),
.Y(n_1370)
);

OAI22x1_ASAP7_75t_L g1371 ( 
.A1(n_1173),
.A2(n_1189),
.B1(n_938),
.B2(n_936),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1140),
.A2(n_933),
.B(n_995),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1172),
.B(n_933),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1196),
.Y(n_1374)
);

A2O1A1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1199),
.A2(n_933),
.B(n_938),
.C(n_936),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1234),
.A2(n_933),
.B(n_934),
.Y(n_1376)
);

AOI221x1_ASAP7_75t_L g1377 ( 
.A1(n_1170),
.A2(n_995),
.B1(n_1125),
.B2(n_1175),
.C(n_1113),
.Y(n_1377)
);

AO31x2_ASAP7_75t_L g1378 ( 
.A1(n_1229),
.A2(n_1263),
.A3(n_1260),
.B(n_1257),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1172),
.B(n_933),
.Y(n_1379)
);

INVxp67_ASAP7_75t_L g1380 ( 
.A(n_1141),
.Y(n_1380)
);

INVxp67_ASAP7_75t_SL g1381 ( 
.A(n_1141),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1251),
.A2(n_1266),
.B(n_1258),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1234),
.A2(n_933),
.B(n_934),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1172),
.B(n_933),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1259),
.A2(n_1255),
.B(n_1248),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1194),
.A2(n_667),
.B1(n_680),
.B2(n_936),
.Y(n_1386)
);

AOI221x1_ASAP7_75t_L g1387 ( 
.A1(n_1170),
.A2(n_995),
.B1(n_1125),
.B2(n_1175),
.C(n_1113),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1199),
.A2(n_933),
.B(n_650),
.C(n_631),
.Y(n_1388)
);

A2O1A1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1199),
.A2(n_933),
.B(n_938),
.C(n_936),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1172),
.B(n_933),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1137),
.B(n_794),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1172),
.B(n_933),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1148),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1234),
.A2(n_933),
.B(n_934),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1140),
.A2(n_933),
.B(n_995),
.Y(n_1395)
);

NAND3xp33_ASAP7_75t_L g1396 ( 
.A(n_1199),
.B(n_933),
.C(n_936),
.Y(n_1396)
);

AOI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1268),
.A2(n_1258),
.B(n_1257),
.Y(n_1397)
);

O2A1O1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1199),
.A2(n_933),
.B(n_650),
.C(n_631),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1251),
.A2(n_1266),
.B(n_1258),
.Y(n_1399)
);

NAND3xp33_ASAP7_75t_SL g1400 ( 
.A(n_1173),
.B(n_684),
.C(n_667),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1234),
.A2(n_933),
.B(n_934),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1178),
.A2(n_933),
.B1(n_995),
.B2(n_932),
.Y(n_1402)
);

AO31x2_ASAP7_75t_L g1403 ( 
.A1(n_1229),
.A2(n_1263),
.A3(n_1260),
.B(n_1257),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1194),
.A2(n_667),
.B1(n_680),
.B2(n_936),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1154),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1234),
.A2(n_933),
.B(n_934),
.Y(n_1406)
);

NOR2xp67_ASAP7_75t_L g1407 ( 
.A(n_1236),
.B(n_827),
.Y(n_1407)
);

INVx1_ASAP7_75t_SL g1408 ( 
.A(n_1154),
.Y(n_1408)
);

AO31x2_ASAP7_75t_L g1409 ( 
.A1(n_1229),
.A2(n_1263),
.A3(n_1260),
.B(n_1257),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1251),
.A2(n_1266),
.B(n_1258),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1178),
.A2(n_933),
.B1(n_995),
.B2(n_932),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1140),
.A2(n_933),
.B(n_995),
.Y(n_1412)
);

AOI221xp5_ASAP7_75t_SL g1413 ( 
.A1(n_1122),
.A2(n_933),
.B1(n_1088),
.B2(n_1199),
.C(n_995),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1116),
.A2(n_864),
.B1(n_788),
.B2(n_1054),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1251),
.A2(n_1266),
.B(n_1258),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1154),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1191),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1153),
.Y(n_1418)
);

BUFx10_ASAP7_75t_L g1419 ( 
.A(n_1209),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1140),
.A2(n_933),
.B(n_995),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1234),
.A2(n_933),
.B(n_934),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1234),
.A2(n_933),
.B(n_934),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1251),
.A2(n_1266),
.B(n_1258),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_SL g1424 ( 
.A(n_1299),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1347),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1405),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1414),
.A2(n_1362),
.B1(n_1278),
.B2(n_1370),
.Y(n_1427)
);

INVx4_ASAP7_75t_L g1428 ( 
.A(n_1275),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1378),
.Y(n_1429)
);

NAND2x1p5_ASAP7_75t_L g1430 ( 
.A(n_1300),
.B(n_1270),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1346),
.A2(n_1372),
.B1(n_1412),
.B2(n_1395),
.Y(n_1431)
);

CKINVDCx11_ASAP7_75t_R g1432 ( 
.A(n_1374),
.Y(n_1432)
);

INVx6_ASAP7_75t_L g1433 ( 
.A(n_1419),
.Y(n_1433)
);

INVx6_ASAP7_75t_L g1434 ( 
.A(n_1419),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1362),
.A2(n_1281),
.B1(n_1308),
.B2(n_1402),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_SL g1436 ( 
.A1(n_1281),
.A2(n_1308),
.B1(n_1411),
.B2(n_1402),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1303),
.B(n_1349),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1317),
.Y(n_1438)
);

BUFx4_ASAP7_75t_SL g1439 ( 
.A(n_1277),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_1352),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1366),
.B(n_1391),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1293),
.Y(n_1442)
);

BUFx4f_ASAP7_75t_SL g1443 ( 
.A(n_1363),
.Y(n_1443)
);

CKINVDCx11_ASAP7_75t_R g1444 ( 
.A(n_1270),
.Y(n_1444)
);

CKINVDCx11_ASAP7_75t_R g1445 ( 
.A(n_1408),
.Y(n_1445)
);

INVx4_ASAP7_75t_SL g1446 ( 
.A(n_1335),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1411),
.B(n_1346),
.Y(n_1447)
);

BUFx4f_ASAP7_75t_SL g1448 ( 
.A(n_1408),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1358),
.A2(n_1368),
.B1(n_1404),
.B2(n_1386),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1311),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1371),
.A2(n_1400),
.B1(n_1283),
.B2(n_1306),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1350),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1359),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1283),
.A2(n_1420),
.B1(n_1372),
.B2(n_1395),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1412),
.A2(n_1420),
.B1(n_1309),
.B2(n_1417),
.Y(n_1455)
);

INVx6_ASAP7_75t_L g1456 ( 
.A(n_1311),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1392),
.A2(n_1288),
.B1(n_1285),
.B2(n_1379),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1320),
.Y(n_1458)
);

BUFx10_ASAP7_75t_L g1459 ( 
.A(n_1354),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1375),
.A2(n_1389),
.B1(n_1357),
.B2(n_1396),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1282),
.B(n_1271),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1392),
.A2(n_1390),
.B1(n_1384),
.B2(n_1373),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1276),
.B(n_1378),
.Y(n_1463)
);

BUFx12f_ASAP7_75t_L g1464 ( 
.A(n_1296),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1290),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1403),
.B(n_1409),
.Y(n_1466)
);

CKINVDCx11_ASAP7_75t_R g1467 ( 
.A(n_1328),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1365),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1291),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1357),
.A2(n_1396),
.B1(n_1321),
.B2(n_1313),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1381),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1334),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1388),
.A2(n_1398),
.B1(n_1321),
.B2(n_1292),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_1296),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1336),
.Y(n_1475)
);

BUFx4_ASAP7_75t_SL g1476 ( 
.A(n_1338),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1284),
.A2(n_1328),
.B1(n_1337),
.B2(n_1407),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1342),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1273),
.A2(n_1327),
.B1(n_1369),
.B2(n_1380),
.Y(n_1479)
);

INVx6_ASAP7_75t_L g1480 ( 
.A(n_1315),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1418),
.Y(n_1481)
);

BUFx10_ASAP7_75t_L g1482 ( 
.A(n_1393),
.Y(n_1482)
);

OAI22xp33_ASAP7_75t_SL g1483 ( 
.A1(n_1367),
.A2(n_1337),
.B1(n_1272),
.B2(n_1416),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1279),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1397),
.Y(n_1485)
);

INVx6_ASAP7_75t_L g1486 ( 
.A(n_1325),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1273),
.A2(n_1421),
.B1(n_1361),
.B2(n_1383),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1327),
.A2(n_1353),
.B1(n_1394),
.B2(n_1401),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1376),
.A2(n_1406),
.B1(n_1422),
.B2(n_1316),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1316),
.A2(n_1318),
.B1(n_1307),
.B2(n_1304),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1347),
.A2(n_1319),
.B1(n_1326),
.B2(n_1333),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1305),
.Y(n_1492)
);

CKINVDCx6p67_ASAP7_75t_R g1493 ( 
.A(n_1325),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1297),
.A2(n_1289),
.B1(n_1323),
.B2(n_1385),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1340),
.Y(n_1495)
);

CKINVDCx11_ASAP7_75t_R g1496 ( 
.A(n_1341),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1343),
.B(n_1344),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1340),
.B(n_1335),
.Y(n_1498)
);

BUFx4_ASAP7_75t_SL g1499 ( 
.A(n_1332),
.Y(n_1499)
);

OAI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1377),
.A2(n_1387),
.B1(n_1301),
.B2(n_1287),
.Y(n_1500)
);

BUFx6f_ASAP7_75t_L g1501 ( 
.A(n_1310),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1345),
.Y(n_1502)
);

NAND2x1p5_ASAP7_75t_L g1503 ( 
.A(n_1339),
.B(n_1331),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_SL g1504 ( 
.A1(n_1413),
.A2(n_1385),
.B1(n_1310),
.B2(n_1295),
.Y(n_1504)
);

INVx6_ASAP7_75t_L g1505 ( 
.A(n_1340),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1274),
.A2(n_1324),
.B1(n_1330),
.B2(n_1280),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1322),
.Y(n_1507)
);

INVx5_ASAP7_75t_SL g1508 ( 
.A(n_1294),
.Y(n_1508)
);

CKINVDCx11_ASAP7_75t_R g1509 ( 
.A(n_1286),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1329),
.Y(n_1510)
);

CKINVDCx20_ASAP7_75t_R g1511 ( 
.A(n_1314),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1302),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1413),
.A2(n_1298),
.B1(n_1360),
.B2(n_1364),
.Y(n_1513)
);

OAI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1312),
.A2(n_1348),
.B1(n_1382),
.B2(n_1351),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1312),
.A2(n_1355),
.B1(n_1356),
.B2(n_1399),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1410),
.A2(n_1415),
.B1(n_1423),
.B2(n_1269),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1317),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_SL g1518 ( 
.A1(n_1362),
.A2(n_1194),
.B1(n_1281),
.B2(n_1116),
.Y(n_1518)
);

INVx4_ASAP7_75t_L g1519 ( 
.A(n_1275),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1275),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1317),
.Y(n_1521)
);

CKINVDCx11_ASAP7_75t_R g1522 ( 
.A(n_1374),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1317),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1317),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1275),
.Y(n_1525)
);

OAI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1358),
.A2(n_1386),
.B1(n_1404),
.B2(n_1368),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1275),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1414),
.A2(n_1362),
.B1(n_864),
.B2(n_788),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1275),
.Y(n_1529)
);

CKINVDCx11_ASAP7_75t_R g1530 ( 
.A(n_1374),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1346),
.A2(n_933),
.B1(n_995),
.B2(n_1372),
.Y(n_1531)
);

INVx8_ASAP7_75t_L g1532 ( 
.A(n_1363),
.Y(n_1532)
);

INVx6_ASAP7_75t_L g1533 ( 
.A(n_1419),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1414),
.A2(n_1362),
.B1(n_864),
.B2(n_788),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1405),
.Y(n_1535)
);

CKINVDCx20_ASAP7_75t_R g1536 ( 
.A(n_1374),
.Y(n_1536)
);

CKINVDCx11_ASAP7_75t_R g1537 ( 
.A(n_1374),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_1374),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1317),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1362),
.A2(n_1194),
.B1(n_1281),
.B2(n_1116),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1414),
.A2(n_1362),
.B1(n_864),
.B2(n_788),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1414),
.A2(n_1362),
.B1(n_864),
.B2(n_788),
.Y(n_1542)
);

INVx4_ASAP7_75t_L g1543 ( 
.A(n_1275),
.Y(n_1543)
);

INVx6_ASAP7_75t_L g1544 ( 
.A(n_1419),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1317),
.Y(n_1545)
);

INVxp67_ASAP7_75t_SL g1546 ( 
.A(n_1385),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1317),
.Y(n_1547)
);

BUFx4f_ASAP7_75t_SL g1548 ( 
.A(n_1374),
.Y(n_1548)
);

BUFx10_ASAP7_75t_L g1549 ( 
.A(n_1354),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1414),
.A2(n_1362),
.B1(n_864),
.B2(n_788),
.Y(n_1550)
);

INVx8_ASAP7_75t_L g1551 ( 
.A(n_1363),
.Y(n_1551)
);

OAI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1375),
.A2(n_1389),
.B(n_1388),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1317),
.Y(n_1553)
);

CKINVDCx6p67_ASAP7_75t_R g1554 ( 
.A(n_1299),
.Y(n_1554)
);

INVx4_ASAP7_75t_L g1555 ( 
.A(n_1275),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1414),
.A2(n_1362),
.B1(n_864),
.B2(n_788),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1317),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1374),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1275),
.Y(n_1559)
);

INVx8_ASAP7_75t_L g1560 ( 
.A(n_1363),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1402),
.B(n_1411),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1317),
.Y(n_1562)
);

BUFx8_ASAP7_75t_SL g1563 ( 
.A(n_1374),
.Y(n_1563)
);

CKINVDCx11_ASAP7_75t_R g1564 ( 
.A(n_1374),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1414),
.A2(n_1362),
.B1(n_864),
.B2(n_788),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1484),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1471),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1461),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1485),
.Y(n_1569)
);

CKINVDCx11_ASAP7_75t_R g1570 ( 
.A(n_1432),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1446),
.B(n_1498),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1446),
.B(n_1495),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1429),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1435),
.A2(n_1518),
.B1(n_1540),
.B2(n_1526),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1429),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1468),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1466),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1466),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1447),
.Y(n_1579)
);

OA21x2_ASAP7_75t_L g1580 ( 
.A1(n_1463),
.A2(n_1506),
.B(n_1552),
.Y(n_1580)
);

AOI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1531),
.A2(n_1561),
.B(n_1431),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1447),
.Y(n_1582)
);

NAND2x1p5_ASAP7_75t_L g1583 ( 
.A(n_1510),
.B(n_1502),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1426),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1535),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1436),
.B(n_1442),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1463),
.Y(n_1587)
);

AO31x2_ASAP7_75t_L g1588 ( 
.A1(n_1431),
.A2(n_1473),
.A3(n_1487),
.B(n_1531),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1505),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_1511),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1472),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1546),
.Y(n_1592)
);

INVxp67_ASAP7_75t_L g1593 ( 
.A(n_1437),
.Y(n_1593)
);

OA21x2_ASAP7_75t_L g1594 ( 
.A1(n_1552),
.A2(n_1490),
.B(n_1489),
.Y(n_1594)
);

NAND4xp25_ASAP7_75t_SL g1595 ( 
.A(n_1518),
.B(n_1540),
.C(n_1427),
.D(n_1436),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1452),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1546),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1458),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1475),
.Y(n_1599)
);

INVx6_ASAP7_75t_L g1600 ( 
.A(n_1428),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1465),
.B(n_1469),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1454),
.B(n_1435),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1478),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1441),
.B(n_1497),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1438),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1517),
.B(n_1521),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1503),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1503),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1512),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1523),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1449),
.A2(n_1451),
.B1(n_1526),
.B2(n_1470),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1524),
.B(n_1539),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1508),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1545),
.B(n_1547),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1553),
.Y(n_1615)
);

INVx4_ASAP7_75t_L g1616 ( 
.A(n_1507),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1557),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1562),
.B(n_1479),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1504),
.B(n_1455),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1433),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1528),
.A2(n_1565),
.B1(n_1534),
.B2(n_1541),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1504),
.B(n_1462),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1508),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1514),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1514),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1460),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1453),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1433),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1460),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1448),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1448),
.B(n_1444),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1491),
.B(n_1494),
.Y(n_1632)
);

INVxp67_ASAP7_75t_SL g1633 ( 
.A(n_1500),
.Y(n_1633)
);

AO21x1_ASAP7_75t_L g1634 ( 
.A1(n_1473),
.A2(n_1500),
.B(n_1487),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1457),
.B(n_1513),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1515),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1515),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1516),
.Y(n_1638)
);

BUFx4f_ASAP7_75t_SL g1639 ( 
.A(n_1536),
.Y(n_1639)
);

NAND2x1p5_ASAP7_75t_L g1640 ( 
.A(n_1501),
.B(n_1477),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1499),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1430),
.Y(n_1642)
);

BUFx3_ASAP7_75t_L g1643 ( 
.A(n_1496),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1499),
.Y(n_1644)
);

BUFx3_ASAP7_75t_L g1645 ( 
.A(n_1493),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1483),
.B(n_1508),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1488),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1450),
.B(n_1481),
.Y(n_1648)
);

AO21x2_ASAP7_75t_L g1649 ( 
.A1(n_1509),
.A2(n_1542),
.B(n_1556),
.Y(n_1649)
);

OR2x6_ASAP7_75t_L g1650 ( 
.A(n_1434),
.B(n_1533),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1550),
.A2(n_1440),
.B(n_1425),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1476),
.A2(n_1486),
.B(n_1480),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1445),
.B(n_1459),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1486),
.B(n_1480),
.Y(n_1654)
);

OAI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1464),
.A2(n_1527),
.B1(n_1529),
.B2(n_1525),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1486),
.Y(n_1656)
);

BUFx2_ASAP7_75t_L g1657 ( 
.A(n_1456),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1428),
.B(n_1543),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1434),
.Y(n_1659)
);

NOR2x1p5_ASAP7_75t_L g1660 ( 
.A(n_1520),
.B(n_1559),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1519),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1519),
.B(n_1555),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1459),
.B(n_1549),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1533),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1543),
.A2(n_1555),
.B(n_1532),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1605),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1568),
.B(n_1554),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1570),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1579),
.B(n_1549),
.Y(n_1669)
);

A2O1A1Ixp33_ASAP7_75t_L g1670 ( 
.A1(n_1574),
.A2(n_1532),
.B(n_1551),
.C(n_1560),
.Y(n_1670)
);

AO32x2_ASAP7_75t_L g1671 ( 
.A1(n_1589),
.A2(n_1467),
.A3(n_1544),
.B1(n_1482),
.B2(n_1439),
.Y(n_1671)
);

O2A1O1Ixp33_ASAP7_75t_L g1672 ( 
.A1(n_1611),
.A2(n_1474),
.B(n_1538),
.C(n_1439),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1610),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1660),
.B(n_1492),
.Y(n_1674)
);

AOI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1595),
.A2(n_1424),
.B1(n_1560),
.B2(n_1551),
.C(n_1532),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1567),
.B(n_1558),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_SL g1677 ( 
.A1(n_1574),
.A2(n_1424),
.B(n_1544),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1660),
.B(n_1544),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1604),
.B(n_1482),
.Y(n_1679)
);

OAI211xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1581),
.A2(n_1564),
.B(n_1522),
.C(n_1530),
.Y(n_1680)
);

A2O1A1Ixp33_ASAP7_75t_L g1681 ( 
.A1(n_1602),
.A2(n_1644),
.B(n_1641),
.C(n_1622),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1579),
.B(n_1551),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1582),
.B(n_1560),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1604),
.B(n_1537),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1590),
.B(n_1548),
.Y(n_1685)
);

INVx4_ASAP7_75t_L g1686 ( 
.A(n_1613),
.Y(n_1686)
);

AOI221xp5_ASAP7_75t_L g1687 ( 
.A1(n_1602),
.A2(n_1443),
.B1(n_1548),
.B2(n_1563),
.C(n_1633),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1652),
.B(n_1571),
.Y(n_1688)
);

OAI211xp5_ASAP7_75t_L g1689 ( 
.A1(n_1626),
.A2(n_1629),
.B(n_1622),
.C(n_1586),
.Y(n_1689)
);

OAI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1626),
.A2(n_1629),
.B1(n_1586),
.B2(n_1621),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1576),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1590),
.B(n_1593),
.Y(n_1692)
);

OA21x2_ASAP7_75t_L g1693 ( 
.A1(n_1634),
.A2(n_1625),
.B(n_1624),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1652),
.B(n_1571),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1617),
.B(n_1591),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1599),
.B(n_1603),
.Y(n_1696)
);

INVxp33_ASAP7_75t_L g1697 ( 
.A(n_1653),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1619),
.A2(n_1647),
.B(n_1594),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1590),
.B(n_1584),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1639),
.B(n_1630),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1644),
.A2(n_1643),
.B1(n_1627),
.B2(n_1631),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1598),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1571),
.B(n_1572),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_SL g1704 ( 
.A1(n_1649),
.A2(n_1619),
.B1(n_1632),
.B2(n_1635),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1585),
.B(n_1630),
.Y(n_1705)
);

OAI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1647),
.A2(n_1594),
.B(n_1635),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1627),
.B(n_1663),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1663),
.B(n_1648),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1661),
.Y(n_1709)
);

AO32x2_ASAP7_75t_L g1710 ( 
.A1(n_1589),
.A2(n_1620),
.A3(n_1628),
.B1(n_1616),
.B2(n_1634),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1587),
.B(n_1588),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_SL g1712 ( 
.A1(n_1594),
.A2(n_1643),
.B(n_1616),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1572),
.B(n_1650),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1596),
.Y(n_1714)
);

OR2x6_ASAP7_75t_L g1715 ( 
.A(n_1583),
.B(n_1632),
.Y(n_1715)
);

OR2x6_ASAP7_75t_L g1716 ( 
.A(n_1583),
.B(n_1632),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1657),
.B(n_1654),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1636),
.A2(n_1637),
.B1(n_1624),
.B2(n_1625),
.C(n_1615),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1613),
.B(n_1623),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1654),
.B(n_1659),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1580),
.Y(n_1721)
);

OAI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1580),
.A2(n_1637),
.B(n_1636),
.Y(n_1722)
);

AOI211xp5_ASAP7_75t_L g1723 ( 
.A1(n_1651),
.A2(n_1646),
.B(n_1618),
.C(n_1655),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1588),
.B(n_1577),
.Y(n_1724)
);

AOI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1649),
.A2(n_1638),
.B1(n_1618),
.B2(n_1614),
.C(n_1612),
.Y(n_1725)
);

OAI21x1_ASAP7_75t_SL g1726 ( 
.A1(n_1665),
.A2(n_1616),
.B(n_1628),
.Y(n_1726)
);

A2O1A1Ixp33_ASAP7_75t_L g1727 ( 
.A1(n_1643),
.A2(n_1638),
.B(n_1613),
.C(n_1623),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1601),
.B(n_1588),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1658),
.B(n_1662),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1658),
.B(n_1662),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1606),
.B(n_1612),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1580),
.A2(n_1607),
.B(n_1608),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1728),
.B(n_1588),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1702),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1731),
.B(n_1588),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1690),
.A2(n_1649),
.B1(n_1601),
.B2(n_1578),
.Y(n_1736)
);

INVxp67_ASAP7_75t_SL g1737 ( 
.A(n_1721),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1711),
.B(n_1592),
.Y(n_1738)
);

BUFx3_ASAP7_75t_L g1739 ( 
.A(n_1688),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1711),
.B(n_1592),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1704),
.A2(n_1569),
.B1(n_1640),
.B2(n_1566),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1710),
.B(n_1597),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1710),
.B(n_1597),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1691),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1710),
.B(n_1609),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1696),
.Y(n_1746)
);

BUFx3_ASAP7_75t_L g1747 ( 
.A(n_1694),
.Y(n_1747)
);

OAI221xp5_ASAP7_75t_SL g1748 ( 
.A1(n_1689),
.A2(n_1675),
.B1(n_1687),
.B2(n_1725),
.C(n_1681),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1724),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1714),
.Y(n_1750)
);

NOR2x1p5_ASAP7_75t_L g1751 ( 
.A(n_1686),
.B(n_1623),
.Y(n_1751)
);

BUFx2_ASAP7_75t_L g1752 ( 
.A(n_1671),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1695),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1693),
.B(n_1566),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1693),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1671),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1666),
.B(n_1575),
.Y(n_1757)
);

INVx3_ASAP7_75t_L g1758 ( 
.A(n_1694),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1732),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1671),
.Y(n_1760)
);

INVxp67_ASAP7_75t_SL g1761 ( 
.A(n_1669),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1673),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1754),
.Y(n_1763)
);

AO21x2_ASAP7_75t_L g1764 ( 
.A1(n_1759),
.A2(n_1698),
.B(n_1706),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1761),
.B(n_1669),
.Y(n_1765)
);

NAND4xp25_ASAP7_75t_L g1766 ( 
.A(n_1752),
.B(n_1687),
.C(n_1683),
.D(n_1682),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1754),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1735),
.B(n_1699),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1761),
.B(n_1709),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1736),
.A2(n_1675),
.B1(n_1725),
.B2(n_1723),
.Y(n_1770)
);

OAI321xp33_ASAP7_75t_L g1771 ( 
.A1(n_1748),
.A2(n_1706),
.A3(n_1722),
.B1(n_1718),
.B2(n_1723),
.C(n_1716),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1739),
.B(n_1703),
.Y(n_1772)
);

OAI322xp33_ASAP7_75t_L g1773 ( 
.A1(n_1733),
.A2(n_1712),
.A3(n_1683),
.B1(n_1682),
.B2(n_1701),
.C1(n_1677),
.C2(n_1676),
.Y(n_1773)
);

OAI211xp5_ASAP7_75t_L g1774 ( 
.A1(n_1752),
.A2(n_1672),
.B(n_1680),
.C(n_1722),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1754),
.Y(n_1775)
);

OAI211xp5_ASAP7_75t_SL g1776 ( 
.A1(n_1762),
.A2(n_1667),
.B(n_1707),
.C(n_1700),
.Y(n_1776)
);

OR2x6_ASAP7_75t_L g1777 ( 
.A(n_1760),
.B(n_1715),
.Y(n_1777)
);

OAI221xp5_ASAP7_75t_L g1778 ( 
.A1(n_1748),
.A2(n_1670),
.B1(n_1727),
.B2(n_1701),
.C(n_1715),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1735),
.B(n_1705),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1757),
.Y(n_1780)
);

AOI21xp33_ASAP7_75t_L g1781 ( 
.A1(n_1755),
.A2(n_1697),
.B(n_1656),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1735),
.B(n_1708),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1757),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1757),
.Y(n_1784)
);

AND4x1_ASAP7_75t_L g1785 ( 
.A(n_1741),
.B(n_1685),
.C(n_1684),
.D(n_1692),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1757),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1758),
.B(n_1717),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1758),
.B(n_1730),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1734),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1754),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1742),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1758),
.B(n_1679),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1750),
.Y(n_1793)
);

INVxp67_ASAP7_75t_SL g1794 ( 
.A(n_1755),
.Y(n_1794)
);

NOR3xp33_ASAP7_75t_L g1795 ( 
.A(n_1748),
.B(n_1664),
.C(n_1719),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1758),
.B(n_1729),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1739),
.B(n_1720),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1739),
.B(n_1703),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1744),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1750),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1742),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1744),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1746),
.B(n_1573),
.Y(n_1803)
);

INVx4_ASAP7_75t_L g1804 ( 
.A(n_1760),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1752),
.A2(n_1716),
.B1(n_1713),
.B2(n_1642),
.Y(n_1805)
);

INVx2_ASAP7_75t_SL g1806 ( 
.A(n_1739),
.Y(n_1806)
);

AND2x6_ASAP7_75t_L g1807 ( 
.A(n_1739),
.B(n_1713),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1750),
.Y(n_1808)
);

INVxp67_ASAP7_75t_SL g1809 ( 
.A(n_1749),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1809),
.B(n_1740),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1785),
.B(n_1760),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1791),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1791),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1801),
.B(n_1733),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1801),
.B(n_1738),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1782),
.B(n_1756),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1789),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1793),
.Y(n_1818)
);

AND2x4_ASAP7_75t_SL g1819 ( 
.A(n_1772),
.B(n_1760),
.Y(n_1819)
);

BUFx3_ASAP7_75t_L g1820 ( 
.A(n_1807),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1764),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1800),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1782),
.B(n_1756),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1779),
.B(n_1756),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1779),
.B(n_1760),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1804),
.B(n_1760),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1764),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1804),
.B(n_1768),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1804),
.B(n_1760),
.Y(n_1829)
);

OR2x6_ASAP7_75t_L g1830 ( 
.A(n_1777),
.B(n_1760),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1768),
.B(n_1760),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1806),
.B(n_1760),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1794),
.B(n_1740),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1780),
.Y(n_1834)
);

INVx3_ASAP7_75t_L g1835 ( 
.A(n_1807),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1806),
.B(n_1742),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1783),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1764),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1784),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1800),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1787),
.B(n_1742),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1786),
.B(n_1740),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1787),
.B(n_1743),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1797),
.B(n_1743),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1808),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1799),
.Y(n_1846)
);

INVxp67_ASAP7_75t_L g1847 ( 
.A(n_1802),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1763),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1808),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1763),
.Y(n_1850)
);

BUFx3_ASAP7_75t_L g1851 ( 
.A(n_1807),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1797),
.B(n_1743),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1803),
.Y(n_1853)
);

AND2x4_ASAP7_75t_L g1854 ( 
.A(n_1807),
.B(n_1747),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1846),
.Y(n_1855)
);

NAND2x1p5_ASAP7_75t_L g1856 ( 
.A(n_1835),
.B(n_1751),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1814),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1817),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1811),
.B(n_1772),
.Y(n_1859)
);

NAND3xp33_ASAP7_75t_SL g1860 ( 
.A(n_1811),
.B(n_1774),
.C(n_1770),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1817),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1853),
.B(n_1753),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1816),
.B(n_1772),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1853),
.B(n_1753),
.Y(n_1864)
);

INVxp67_ASAP7_75t_SL g1865 ( 
.A(n_1821),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1816),
.B(n_1798),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1814),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1814),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1816),
.B(n_1798),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1847),
.B(n_1765),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1847),
.B(n_1740),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1817),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1823),
.B(n_1798),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1846),
.B(n_1743),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1810),
.B(n_1769),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1810),
.B(n_1833),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1823),
.B(n_1795),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1834),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1823),
.B(n_1749),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1824),
.B(n_1749),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1824),
.B(n_1796),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1834),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1837),
.Y(n_1883)
);

INVx2_ASAP7_75t_SL g1884 ( 
.A(n_1820),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1824),
.B(n_1796),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1844),
.B(n_1792),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1837),
.Y(n_1887)
);

OR2x6_ASAP7_75t_L g1888 ( 
.A(n_1830),
.B(n_1777),
.Y(n_1888)
);

INVx6_ASAP7_75t_L g1889 ( 
.A(n_1820),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1839),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1836),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1833),
.B(n_1738),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1839),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1850),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1850),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1850),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1844),
.B(n_1792),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_L g1898 ( 
.A(n_1835),
.B(n_1668),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1818),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1844),
.B(n_1788),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1863),
.B(n_1852),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1891),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1855),
.Y(n_1903)
);

INVxp67_ASAP7_75t_L g1904 ( 
.A(n_1898),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1858),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1863),
.B(n_1866),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1858),
.Y(n_1907)
);

AOI221xp5_ASAP7_75t_L g1908 ( 
.A1(n_1860),
.A2(n_1821),
.B1(n_1838),
.B2(n_1827),
.C(n_1771),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1877),
.B(n_1852),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1861),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1870),
.B(n_1852),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1881),
.B(n_1841),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1881),
.B(n_1841),
.Y(n_1913)
);

INVx1_ASAP7_75t_SL g1914 ( 
.A(n_1889),
.Y(n_1914)
);

AND2x2_ASAP7_75t_SL g1915 ( 
.A(n_1859),
.B(n_1678),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1866),
.B(n_1819),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1889),
.A2(n_1821),
.B1(n_1827),
.B2(n_1838),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1875),
.B(n_1842),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1869),
.B(n_1819),
.Y(n_1919)
);

INVxp67_ASAP7_75t_L g1920 ( 
.A(n_1884),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1875),
.B(n_1842),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_SL g1922 ( 
.A(n_1889),
.B(n_1778),
.Y(n_1922)
);

OAI211xp5_ASAP7_75t_SL g1923 ( 
.A1(n_1884),
.A2(n_1827),
.B(n_1838),
.C(n_1821),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1874),
.A2(n_1773),
.B(n_1862),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1889),
.B(n_1776),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1856),
.B(n_1674),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1885),
.B(n_1841),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1861),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1869),
.B(n_1819),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1891),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1872),
.Y(n_1931)
);

NOR2xp67_ASAP7_75t_L g1932 ( 
.A(n_1859),
.B(n_1835),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1872),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1894),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1885),
.B(n_1843),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1873),
.B(n_1819),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1876),
.B(n_1815),
.Y(n_1937)
);

AOI22xp5_ASAP7_75t_L g1938 ( 
.A1(n_1922),
.A2(n_1838),
.B1(n_1827),
.B2(n_1865),
.Y(n_1938)
);

AOI211xp5_ASAP7_75t_L g1939 ( 
.A1(n_1924),
.A2(n_1826),
.B(n_1829),
.C(n_1851),
.Y(n_1939)
);

OAI332xp33_ASAP7_75t_L g1940 ( 
.A1(n_1914),
.A2(n_1879),
.A3(n_1880),
.B1(n_1876),
.B2(n_1871),
.B3(n_1868),
.C1(n_1857),
.C2(n_1892),
.Y(n_1940)
);

AOI21xp33_ASAP7_75t_L g1941 ( 
.A1(n_1908),
.A2(n_1882),
.B(n_1878),
.Y(n_1941)
);

NOR4xp25_ASAP7_75t_SL g1942 ( 
.A(n_1903),
.B(n_1896),
.C(n_1895),
.D(n_1899),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1906),
.B(n_1873),
.Y(n_1943)
);

OAI31xp33_ASAP7_75t_L g1944 ( 
.A1(n_1923),
.A2(n_1826),
.A3(n_1829),
.B(n_1857),
.Y(n_1944)
);

OAI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1925),
.A2(n_1829),
.B(n_1826),
.Y(n_1945)
);

O2A1O1Ixp33_ASAP7_75t_L g1946 ( 
.A1(n_1934),
.A2(n_1883),
.B(n_1890),
.C(n_1878),
.Y(n_1946)
);

OAI21xp33_ASAP7_75t_SL g1947 ( 
.A1(n_1932),
.A2(n_1906),
.B(n_1901),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1905),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1920),
.B(n_1886),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1937),
.B(n_1864),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1937),
.B(n_1882),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1905),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1910),
.Y(n_1953)
);

OAI32xp33_ASAP7_75t_L g1954 ( 
.A1(n_1909),
.A2(n_1856),
.A3(n_1835),
.B1(n_1892),
.B2(n_1851),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1910),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1901),
.Y(n_1956)
);

NAND3xp33_ASAP7_75t_L g1957 ( 
.A(n_1917),
.B(n_1896),
.C(n_1895),
.Y(n_1957)
);

AOI222xp33_ASAP7_75t_L g1958 ( 
.A1(n_1915),
.A2(n_1911),
.B1(n_1934),
.B2(n_1857),
.C1(n_1868),
.C2(n_1867),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1916),
.B(n_1886),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1902),
.B(n_1897),
.Y(n_1960)
);

OAI21xp33_ASAP7_75t_SL g1961 ( 
.A1(n_1915),
.A2(n_1900),
.B(n_1897),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1933),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1902),
.Y(n_1963)
);

INVxp67_ASAP7_75t_SL g1964 ( 
.A(n_1933),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1907),
.Y(n_1965)
);

AOI221xp5_ASAP7_75t_L g1966 ( 
.A1(n_1941),
.A2(n_1931),
.B1(n_1928),
.B2(n_1930),
.C(n_1868),
.Y(n_1966)
);

OAI22xp33_ASAP7_75t_L g1967 ( 
.A1(n_1938),
.A2(n_1830),
.B1(n_1888),
.B2(n_1820),
.Y(n_1967)
);

AOI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1942),
.A2(n_1940),
.B(n_1939),
.Y(n_1968)
);

AOI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1958),
.A2(n_1926),
.B1(n_1904),
.B2(n_1930),
.Y(n_1969)
);

AOI221xp5_ASAP7_75t_L g1970 ( 
.A1(n_1946),
.A2(n_1867),
.B1(n_1893),
.B2(n_1883),
.C(n_1887),
.Y(n_1970)
);

INVx1_ASAP7_75t_SL g1971 ( 
.A(n_1956),
.Y(n_1971)
);

AOI21xp33_ASAP7_75t_SL g1972 ( 
.A1(n_1947),
.A2(n_1856),
.B(n_1912),
.Y(n_1972)
);

OAI21xp33_ASAP7_75t_L g1973 ( 
.A1(n_1961),
.A2(n_1921),
.B(n_1918),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1964),
.B(n_1887),
.Y(n_1974)
);

INVxp67_ASAP7_75t_SL g1975 ( 
.A(n_1964),
.Y(n_1975)
);

AOI22xp33_ASAP7_75t_L g1976 ( 
.A1(n_1963),
.A2(n_1888),
.B1(n_1830),
.B2(n_1759),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1950),
.B(n_1918),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1950),
.B(n_1921),
.Y(n_1978)
);

OAI32xp33_ASAP7_75t_L g1979 ( 
.A1(n_1956),
.A2(n_1935),
.A3(n_1927),
.B1(n_1913),
.B2(n_1835),
.Y(n_1979)
);

INVxp67_ASAP7_75t_SL g1980 ( 
.A(n_1951),
.Y(n_1980)
);

NAND3xp33_ASAP7_75t_SL g1981 ( 
.A(n_1944),
.B(n_1919),
.C(n_1916),
.Y(n_1981)
);

INVxp67_ASAP7_75t_L g1982 ( 
.A(n_1949),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1943),
.B(n_1919),
.Y(n_1983)
);

NAND3xp33_ASAP7_75t_SL g1984 ( 
.A(n_1943),
.B(n_1936),
.C(n_1929),
.Y(n_1984)
);

OR2x2_ASAP7_75t_L g1985 ( 
.A(n_1960),
.B(n_1900),
.Y(n_1985)
);

AOI221xp5_ASAP7_75t_L g1986 ( 
.A1(n_1957),
.A2(n_1893),
.B1(n_1890),
.B2(n_1775),
.C(n_1790),
.Y(n_1986)
);

INVx2_ASAP7_75t_SL g1987 ( 
.A(n_1959),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1968),
.A2(n_1951),
.B1(n_1965),
.B2(n_1962),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1975),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1972),
.B(n_1959),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1987),
.B(n_1963),
.Y(n_1991)
);

XNOR2x1_ASAP7_75t_L g1992 ( 
.A(n_1969),
.B(n_1674),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1977),
.B(n_1948),
.Y(n_1993)
);

NAND2xp33_ASAP7_75t_SL g1994 ( 
.A(n_1983),
.B(n_1929),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1980),
.Y(n_1995)
);

XNOR2x2_ASAP7_75t_L g1996 ( 
.A(n_1966),
.B(n_1952),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1985),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1974),
.Y(n_1998)
);

XNOR2xp5_ASAP7_75t_L g1999 ( 
.A(n_1984),
.B(n_1678),
.Y(n_1999)
);

AOI222xp33_ASAP7_75t_L g2000 ( 
.A1(n_1971),
.A2(n_1955),
.B1(n_1953),
.B2(n_1954),
.C1(n_1945),
.C2(n_1775),
.Y(n_2000)
);

NAND3xp33_ASAP7_75t_L g2001 ( 
.A(n_2000),
.B(n_1982),
.C(n_1970),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_L g2002 ( 
.A(n_1990),
.B(n_1978),
.Y(n_2002)
);

AND4x1_ASAP7_75t_L g2003 ( 
.A(n_1995),
.B(n_1973),
.C(n_1974),
.D(n_1986),
.Y(n_2003)
);

AOI21xp33_ASAP7_75t_L g2004 ( 
.A1(n_1988),
.A2(n_1979),
.B(n_1967),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1997),
.B(n_1831),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_SL g2006 ( 
.A(n_1993),
.B(n_1981),
.Y(n_2006)
);

NOR4xp25_ASAP7_75t_L g2007 ( 
.A(n_1989),
.B(n_1988),
.C(n_1998),
.D(n_1991),
.Y(n_2007)
);

NOR3xp33_ASAP7_75t_L g2008 ( 
.A(n_1996),
.B(n_1899),
.C(n_1936),
.Y(n_2008)
);

INVxp33_ASAP7_75t_L g2009 ( 
.A(n_1992),
.Y(n_2009)
);

O2A1O1Ixp33_ASAP7_75t_L g2010 ( 
.A1(n_2000),
.A2(n_1976),
.B(n_1790),
.C(n_1767),
.Y(n_2010)
);

NOR2x1_ASAP7_75t_L g2011 ( 
.A(n_1999),
.B(n_1820),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_2005),
.Y(n_2012)
);

A2O1A1Ixp33_ASAP7_75t_L g2013 ( 
.A1(n_2001),
.A2(n_1994),
.B(n_1851),
.C(n_1767),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_2002),
.B(n_2008),
.Y(n_2014)
);

AOI211xp5_ASAP7_75t_L g2015 ( 
.A1(n_2007),
.A2(n_1851),
.B(n_1766),
.C(n_1854),
.Y(n_2015)
);

NOR4xp25_ASAP7_75t_L g2016 ( 
.A(n_2004),
.B(n_1832),
.C(n_1828),
.D(n_1848),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_2006),
.B(n_1836),
.Y(n_2017)
);

AOI22x1_ASAP7_75t_L g2018 ( 
.A1(n_2003),
.A2(n_1828),
.B1(n_2009),
.B2(n_1832),
.Y(n_2018)
);

AOI211xp5_ASAP7_75t_L g2019 ( 
.A1(n_2014),
.A2(n_2010),
.B(n_2011),
.C(n_1854),
.Y(n_2019)
);

AND4x1_ASAP7_75t_L g2020 ( 
.A(n_2016),
.B(n_1828),
.C(n_1831),
.D(n_1825),
.Y(n_2020)
);

AOI211xp5_ASAP7_75t_L g2021 ( 
.A1(n_2013),
.A2(n_1854),
.B(n_1831),
.C(n_1825),
.Y(n_2021)
);

AOI221xp5_ASAP7_75t_L g2022 ( 
.A1(n_2017),
.A2(n_1848),
.B1(n_1781),
.B2(n_1759),
.C(n_1825),
.Y(n_2022)
);

AOI221xp5_ASAP7_75t_L g2023 ( 
.A1(n_2015),
.A2(n_1848),
.B1(n_1745),
.B2(n_1737),
.C(n_1813),
.Y(n_2023)
);

BUFx6f_ASAP7_75t_L g2024 ( 
.A(n_2012),
.Y(n_2024)
);

OAI211xp5_ASAP7_75t_L g2025 ( 
.A1(n_2018),
.A2(n_1832),
.B(n_1836),
.C(n_1843),
.Y(n_2025)
);

NAND4xp25_ASAP7_75t_L g2026 ( 
.A(n_2014),
.B(n_1645),
.C(n_1854),
.D(n_1843),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2024),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_L g2028 ( 
.A(n_2024),
.B(n_1848),
.Y(n_2028)
);

AOI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_2019),
.A2(n_1888),
.B1(n_1830),
.B2(n_1812),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_2020),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_2023),
.B(n_1812),
.Y(n_2031)
);

INVxp33_ASAP7_75t_L g2032 ( 
.A(n_2026),
.Y(n_2032)
);

OAI22xp33_ASAP7_75t_L g2033 ( 
.A1(n_2029),
.A2(n_2022),
.B1(n_1888),
.B2(n_1812),
.Y(n_2033)
);

NAND2x1p5_ASAP7_75t_L g2034 ( 
.A(n_2027),
.B(n_1645),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2028),
.B(n_2021),
.Y(n_2035)
);

XNOR2xp5_ASAP7_75t_L g2036 ( 
.A(n_2034),
.B(n_2032),
.Y(n_2036)
);

AOI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_2036),
.A2(n_2030),
.B1(n_2031),
.B2(n_2033),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2037),
.Y(n_2038)
);

INVx4_ASAP7_75t_L g2039 ( 
.A(n_2037),
.Y(n_2039)
);

AOI21xp33_ASAP7_75t_SL g2040 ( 
.A1(n_2038),
.A2(n_2035),
.B(n_2025),
.Y(n_2040)
);

OAI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_2039),
.A2(n_1813),
.B1(n_1812),
.B2(n_1849),
.Y(n_2041)
);

AOI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_2041),
.A2(n_2039),
.B1(n_1813),
.B2(n_1888),
.Y(n_2042)
);

XNOR2xp5_ASAP7_75t_L g2043 ( 
.A(n_2040),
.B(n_1645),
.Y(n_2043)
);

AOI22xp33_ASAP7_75t_L g2044 ( 
.A1(n_2042),
.A2(n_1813),
.B1(n_1849),
.B2(n_1845),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2044),
.B(n_2043),
.Y(n_2045)
);

AOI221xp5_ASAP7_75t_L g2046 ( 
.A1(n_2045),
.A2(n_1822),
.B1(n_1849),
.B2(n_1845),
.C(n_1840),
.Y(n_2046)
);

OAI221xp5_ASAP7_75t_R g2047 ( 
.A1(n_2046),
.A2(n_1805),
.B1(n_1854),
.B2(n_1600),
.C(n_1726),
.Y(n_2047)
);

OAI211xp5_ASAP7_75t_SL g2048 ( 
.A1(n_2047),
.A2(n_1620),
.B(n_1664),
.C(n_1613),
.Y(n_2048)
);


endmodule