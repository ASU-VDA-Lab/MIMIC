module real_aes_15462_n_376 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_1034;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1441;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1225;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1893;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1872;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1583;
wire n_1250;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_1926;
wire n_898;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1914;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_1612;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1580;
wire n_1000;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1899;
wire n_816;
wire n_1470;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1931;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1868;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g1068 ( .A(n_0), .Y(n_1068) );
AOI22xp33_ASAP7_75t_SL g1354 ( .A1(n_1), .A2(n_333), .B1(n_459), .B2(n_1355), .Y(n_1354) );
INVxp67_ASAP7_75t_SL g1377 ( .A(n_1), .Y(n_1377) );
INVx1_ASAP7_75t_L g831 ( .A(n_2), .Y(n_831) );
AO22x1_ASAP7_75t_L g857 ( .A1(n_2), .A2(n_245), .B1(n_511), .B2(n_759), .Y(n_857) );
INVx1_ASAP7_75t_L g389 ( .A(n_3), .Y(n_389) );
AND2x2_ASAP7_75t_L g440 ( .A(n_3), .B(n_271), .Y(n_440) );
AND2x2_ASAP7_75t_L g501 ( .A(n_3), .B(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_3), .B(n_399), .Y(n_616) );
INVx1_ASAP7_75t_L g841 ( .A(n_4), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_4), .A2(n_123), .B1(n_516), .B2(n_755), .Y(n_856) );
AOI22xp33_ASAP7_75t_SL g1910 ( .A1(n_5), .A2(n_42), .B1(n_459), .B2(n_482), .Y(n_1910) );
INVxp67_ASAP7_75t_SL g1931 ( .A(n_5), .Y(n_1931) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_6), .A2(n_210), .B1(n_474), .B2(n_1076), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_6), .A2(n_189), .B1(n_983), .B2(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1174 ( .A(n_7), .Y(n_1174) );
XOR2x2_ASAP7_75t_L g1386 ( .A(n_8), .B(n_1387), .Y(n_1386) );
INVx1_ASAP7_75t_L g1532 ( .A(n_9), .Y(n_1532) );
OAI22xp5_ASAP7_75t_L g1549 ( .A1(n_9), .A2(n_364), .B1(n_554), .B2(n_873), .Y(n_1549) );
CKINVDCx5p33_ASAP7_75t_R g1567 ( .A(n_10), .Y(n_1567) );
OAI22xp5_ASAP7_75t_L g1245 ( .A1(n_11), .A2(n_233), .B1(n_408), .B2(n_1246), .Y(n_1245) );
AOI22xp33_ASAP7_75t_SL g962 ( .A1(n_12), .A2(n_236), .B1(n_963), .B2(n_964), .Y(n_962) );
INVxp67_ASAP7_75t_SL g1001 ( .A(n_12), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_13), .A2(n_308), .B1(n_1263), .B2(n_1266), .Y(n_1265) );
AOI221xp5_ASAP7_75t_L g1270 ( .A1(n_13), .A2(n_82), .B1(n_755), .B2(n_981), .C(n_1044), .Y(n_1270) );
OAI22xp33_ASAP7_75t_L g1870 ( .A1(n_14), .A2(n_163), .B1(n_1871), .B2(n_1872), .Y(n_1870) );
OAI22xp33_ASAP7_75t_L g1875 ( .A1(n_14), .A2(n_163), .B1(n_391), .B2(n_1876), .Y(n_1875) );
INVx2_ASAP7_75t_L g418 ( .A(n_15), .Y(n_418) );
OAI22xp5_ASAP7_75t_SL g1316 ( .A1(n_16), .A2(n_298), .B1(n_1317), .B2(n_1319), .Y(n_1316) );
OAI221xp5_ASAP7_75t_L g1330 ( .A1(n_16), .A2(n_298), .B1(n_990), .B2(n_1039), .C(n_1331), .Y(n_1330) );
XNOR2x1_ASAP7_75t_L g1293 ( .A(n_17), .B(n_1294), .Y(n_1293) );
AOI22xp5_ASAP7_75t_L g1644 ( .A1(n_17), .A2(n_20), .B1(n_1608), .B2(n_1616), .Y(n_1644) );
AOI22xp33_ASAP7_75t_L g1576 ( .A1(n_18), .A2(n_120), .B1(n_468), .B2(n_1024), .Y(n_1576) );
AOI22xp33_ASAP7_75t_L g1589 ( .A1(n_18), .A2(n_174), .B1(n_625), .B2(n_1538), .Y(n_1589) );
INVx1_ASAP7_75t_L g1222 ( .A(n_19), .Y(n_1222) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_21), .A2(n_243), .B1(n_657), .B2(n_1262), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g1271 ( .A1(n_21), .A2(n_140), .B1(n_1272), .B2(n_1273), .Y(n_1271) );
INVx1_ASAP7_75t_L g929 ( .A(n_22), .Y(n_929) );
OAI22xp33_ASAP7_75t_L g1359 ( .A1(n_23), .A2(n_280), .B1(n_931), .B2(n_1031), .Y(n_1359) );
INVx1_ASAP7_75t_L g1372 ( .A(n_23), .Y(n_1372) );
INVx1_ASAP7_75t_L g1220 ( .A(n_24), .Y(n_1220) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_24), .A2(n_71), .B1(n_984), .B2(n_1052), .Y(n_1236) );
INVx1_ASAP7_75t_L g425 ( .A(n_25), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_26), .A2(n_127), .B1(n_474), .B2(n_1024), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_26), .A2(n_310), .B1(n_984), .B2(n_1052), .Y(n_1051) );
OAI22xp33_ASAP7_75t_L g1584 ( .A1(n_27), .A2(n_226), .B1(n_1030), .B2(n_1031), .Y(n_1584) );
INVx1_ASAP7_75t_L g1591 ( .A(n_27), .Y(n_1591) );
AOI22xp33_ASAP7_75t_SL g1580 ( .A1(n_28), .A2(n_89), .B1(n_461), .B2(n_1266), .Y(n_1580) );
AOI22xp33_ASAP7_75t_SL g1597 ( .A1(n_28), .A2(n_258), .B1(n_1182), .B2(n_1273), .Y(n_1597) );
OAI22xp5_ASAP7_75t_L g1129 ( .A1(n_29), .A2(n_326), .B1(n_554), .B2(n_873), .Y(n_1129) );
CKINVDCx5p33_ASAP7_75t_R g1290 ( .A(n_30), .Y(n_1290) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_31), .Y(n_384) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_31), .B(n_382), .Y(n_1609) );
INVx1_ASAP7_75t_L g1329 ( .A(n_32), .Y(n_1329) );
AOI22xp33_ASAP7_75t_L g1689 ( .A1(n_33), .A2(n_206), .B1(n_1616), .B2(n_1640), .Y(n_1689) );
OAI22xp5_ASAP7_75t_SL g894 ( .A1(n_34), .A2(n_311), .B1(n_895), .B2(n_896), .Y(n_894) );
INVxp67_ASAP7_75t_SL g936 ( .A(n_34), .Y(n_936) );
CKINVDCx5p33_ASAP7_75t_R g941 ( .A(n_35), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_36), .A2(n_235), .B1(n_657), .B2(n_1118), .Y(n_1121) );
AOI221xp5_ASAP7_75t_L g1146 ( .A1(n_36), .A2(n_340), .B1(n_1047), .B2(n_1147), .C(n_1149), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_37), .A2(n_49), .B1(n_470), .B2(n_656), .Y(n_718) );
INVx1_ASAP7_75t_L g730 ( .A(n_37), .Y(n_730) );
INVx1_ASAP7_75t_L g1114 ( .A(n_38), .Y(n_1114) );
OAI221xp5_ASAP7_75t_L g1140 ( .A1(n_38), .A2(n_264), .B1(n_1039), .B2(n_1092), .C(n_1141), .Y(n_1140) );
INVx1_ASAP7_75t_L g627 ( .A(n_39), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_40), .A2(n_47), .B1(n_581), .B2(n_587), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_40), .A2(n_168), .B1(n_655), .B2(n_657), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_41), .A2(n_366), .B1(n_449), .B2(n_708), .C(n_709), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_41), .A2(n_116), .B1(n_519), .B2(n_722), .C(n_729), .Y(n_728) );
AOI221xp5_ASAP7_75t_L g1922 ( .A1(n_42), .A2(n_99), .B1(n_1235), .B2(n_1923), .C(n_1924), .Y(n_1922) );
INVx1_ASAP7_75t_L g1834 ( .A(n_43), .Y(n_1834) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_44), .A2(n_297), .B1(n_785), .B2(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g992 ( .A(n_44), .Y(n_992) );
NAND5xp2_ASAP7_75t_L g745 ( .A(n_45), .B(n_746), .C(n_780), .D(n_797), .E(n_805), .Y(n_745) );
INVx1_ASAP7_75t_L g814 ( .A(n_45), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g1362 ( .A1(n_46), .A2(n_153), .B1(n_554), .B2(n_873), .Y(n_1362) );
OAI211xp5_ASAP7_75t_SL g1364 ( .A1(n_46), .A2(n_1132), .B(n_1365), .C(n_1370), .Y(n_1364) );
AOI22xp33_ASAP7_75t_SL g640 ( .A1(n_47), .A2(n_182), .B1(n_641), .B2(n_643), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g1537 ( .A1(n_48), .A2(n_198), .B1(n_1135), .B2(n_1538), .Y(n_1537) );
AOI22xp33_ASAP7_75t_SL g1556 ( .A1(n_48), .A2(n_343), .B1(n_459), .B2(n_1557), .Y(n_1556) );
INVx1_ASAP7_75t_L g724 ( .A(n_49), .Y(n_724) );
INVx1_ASAP7_75t_L g1865 ( .A(n_50), .Y(n_1865) );
INVxp67_ASAP7_75t_L g1565 ( .A(n_51), .Y(n_1565) );
AOI22xp5_ASAP7_75t_L g1638 ( .A1(n_52), .A2(n_228), .B1(n_1608), .B2(n_1613), .Y(n_1638) );
AOI22xp5_ASAP7_75t_L g1624 ( .A1(n_53), .A2(n_354), .B1(n_1616), .B2(n_1625), .Y(n_1624) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_54), .Y(n_396) );
INVx1_ASAP7_75t_L g1825 ( .A(n_55), .Y(n_1825) );
AOI22xp33_ASAP7_75t_SL g1071 ( .A1(n_56), .A2(n_57), .B1(n_459), .B2(n_964), .Y(n_1071) );
INVx1_ASAP7_75t_L g1094 ( .A(n_56), .Y(n_1094) );
AOI221xp5_ASAP7_75t_L g1083 ( .A1(n_57), .A2(n_137), .B1(n_981), .B2(n_1084), .C(n_1086), .Y(n_1083) );
XOR2x2_ASAP7_75t_L g1524 ( .A(n_58), .B(n_1525), .Y(n_1524) );
XOR2xp5_ASAP7_75t_L g1346 ( .A(n_59), .B(n_1347), .Y(n_1346) );
AOI22xp5_ASAP7_75t_L g1639 ( .A1(n_59), .A2(n_334), .B1(n_1616), .B2(n_1640), .Y(n_1639) );
INVx1_ASAP7_75t_L g950 ( .A(n_60), .Y(n_950) );
AOI22xp5_ASAP7_75t_L g1648 ( .A1(n_61), .A2(n_125), .B1(n_1608), .B2(n_1613), .Y(n_1648) );
INVx1_ASAP7_75t_L g1256 ( .A(n_62), .Y(n_1256) );
OAI222xp33_ASAP7_75t_L g1278 ( .A1(n_62), .A2(n_373), .B1(n_1004), .B2(n_1038), .C1(n_1279), .C2(n_1284), .Y(n_1278) );
AOI22xp33_ASAP7_75t_SL g1356 ( .A1(n_63), .A2(n_305), .B1(n_959), .B2(n_1024), .Y(n_1356) );
AOI221xp5_ASAP7_75t_L g1380 ( .A1(n_63), .A2(n_272), .B1(n_977), .B2(n_979), .C(n_1338), .Y(n_1380) );
INVx1_ASAP7_75t_L g1328 ( .A(n_64), .Y(n_1328) );
AOI22xp33_ASAP7_75t_L g1911 ( .A1(n_65), .A2(n_282), .B1(n_474), .B2(n_1912), .Y(n_1911) );
AOI22xp33_ASAP7_75t_L g1925 ( .A1(n_65), .A2(n_142), .B1(n_525), .B2(n_532), .Y(n_1925) );
CKINVDCx5p33_ASAP7_75t_R g1277 ( .A(n_66), .Y(n_1277) );
AOI221xp5_ASAP7_75t_L g754 ( .A1(n_67), .A2(n_178), .B1(n_516), .B2(n_755), .C(n_757), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_67), .A2(n_251), .B1(n_657), .B2(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g489 ( .A(n_68), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_69), .A2(n_251), .B1(n_753), .B2(n_759), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_69), .A2(n_178), .B1(n_657), .B2(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g1400 ( .A(n_70), .Y(n_1400) );
INVx1_ASAP7_75t_L g1209 ( .A(n_71), .Y(n_1209) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_72), .A2(n_353), .B1(n_591), .B2(n_594), .C(n_598), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_72), .A2(n_313), .B1(n_647), .B2(n_649), .C(n_652), .Y(n_646) );
AOI22xp33_ASAP7_75t_SL g458 ( .A1(n_73), .A2(n_304), .B1(n_459), .B2(n_461), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_73), .A2(n_324), .B1(n_525), .B2(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g953 ( .A1(n_74), .A2(n_185), .B1(n_647), .B2(n_954), .Y(n_953) );
INVxp67_ASAP7_75t_SL g998 ( .A(n_74), .Y(n_998) );
OAI211xp5_ASAP7_75t_SL g698 ( .A1(n_75), .A2(n_666), .B(n_673), .C(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g735 ( .A(n_75), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g1430 ( .A1(n_76), .A2(n_270), .B1(n_1431), .B2(n_1435), .Y(n_1430) );
OAI22xp5_ASAP7_75t_L g1468 ( .A1(n_76), .A2(n_270), .B1(n_1469), .B2(n_1471), .Y(n_1468) );
CKINVDCx5p33_ASAP7_75t_R g770 ( .A(n_77), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_78), .A2(n_249), .B1(n_482), .B2(n_963), .Y(n_1166) );
AOI22xp33_ASAP7_75t_SL g1192 ( .A1(n_78), .A2(n_306), .B1(n_523), .B2(n_1089), .Y(n_1192) );
INVxp67_ASAP7_75t_SL g633 ( .A(n_79), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_79), .A2(n_362), .B1(n_659), .B2(n_662), .Y(n_658) );
AOI22xp33_ASAP7_75t_SL g1122 ( .A1(n_80), .A2(n_369), .B1(n_459), .B2(n_1123), .Y(n_1122) );
AOI221xp5_ASAP7_75t_L g1136 ( .A1(n_80), .A2(n_147), .B1(n_515), .B2(n_762), .C(n_1045), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1914 ( .A1(n_81), .A2(n_99), .B1(n_482), .B2(n_1021), .Y(n_1914) );
INVxp67_ASAP7_75t_SL g1932 ( .A(n_81), .Y(n_1932) );
AOI22xp33_ASAP7_75t_L g1261 ( .A1(n_82), .A2(n_130), .B1(n_1262), .B2(n_1263), .Y(n_1261) );
AOI22xp33_ASAP7_75t_SL g1165 ( .A1(n_83), .A2(n_240), .B1(n_643), .B2(n_1163), .Y(n_1165) );
INVx1_ASAP7_75t_L g1188 ( .A(n_83), .Y(n_1188) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_84), .A2(n_554), .B(n_563), .Y(n_553) );
AOI22xp33_ASAP7_75t_SL g1504 ( .A1(n_85), .A2(n_218), .B1(n_657), .B2(n_785), .Y(n_1504) );
AOI22xp33_ASAP7_75t_L g1515 ( .A1(n_85), .A2(n_94), .B1(n_523), .B2(n_526), .Y(n_1515) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_86), .A2(n_166), .B1(n_511), .B2(n_900), .Y(n_899) );
INVxp67_ASAP7_75t_SL g925 ( .A(n_86), .Y(n_925) );
INVx1_ASAP7_75t_L g1297 ( .A(n_87), .Y(n_1297) );
AOI22xp33_ASAP7_75t_SL g1306 ( .A1(n_88), .A2(n_299), .B1(n_783), .B2(n_927), .Y(n_1306) );
AOI221xp5_ASAP7_75t_L g1323 ( .A1(n_88), .A2(n_95), .B1(n_515), .B2(n_762), .C(n_980), .Y(n_1323) );
AOI221xp5_ASAP7_75t_L g1588 ( .A1(n_89), .A2(n_338), .B1(n_520), .B2(n_755), .C(n_1149), .Y(n_1588) );
INVx1_ASAP7_75t_L g1008 ( .A(n_90), .Y(n_1008) );
AOI22xp5_ASAP7_75t_L g1629 ( .A1(n_91), .A2(n_367), .B1(n_1608), .B2(n_1613), .Y(n_1629) );
OAI21xp33_ASAP7_75t_L g1287 ( .A1(n_92), .A2(n_1246), .B(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1300 ( .A(n_93), .Y(n_1300) );
AOI22xp33_ASAP7_75t_SL g1507 ( .A1(n_94), .A2(n_307), .B1(n_657), .B2(n_785), .Y(n_1507) );
AOI22xp33_ASAP7_75t_L g1314 ( .A1(n_95), .A2(n_202), .B1(n_647), .B2(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1397 ( .A(n_96), .Y(n_1397) );
INVx1_ASAP7_75t_L g1219 ( .A(n_97), .Y(n_1219) );
AOI221xp5_ASAP7_75t_L g1230 ( .A1(n_97), .A2(n_242), .B1(n_1044), .B2(n_1047), .C(n_1086), .Y(n_1230) );
CKINVDCx5p33_ASAP7_75t_R g1500 ( .A(n_98), .Y(n_1500) );
AOI22xp5_ASAP7_75t_SL g1630 ( .A1(n_100), .A2(n_238), .B1(n_1616), .B2(n_1625), .Y(n_1630) );
INVx1_ASAP7_75t_L g1829 ( .A(n_101), .Y(n_1829) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_102), .A2(n_335), .B1(n_463), .B2(n_468), .Y(n_462) );
AOI221xp5_ASAP7_75t_L g533 ( .A1(n_102), .A2(n_359), .B1(n_534), .B2(n_538), .C(n_542), .Y(n_533) );
OAI211xp5_ASAP7_75t_L g764 ( .A1(n_103), .A2(n_765), .B(n_767), .C(n_769), .Y(n_764) );
INVx1_ASAP7_75t_L g810 ( .A(n_103), .Y(n_810) );
INVx1_ASAP7_75t_L g1066 ( .A(n_104), .Y(n_1066) );
OAI221xp5_ASAP7_75t_L g1091 ( .A1(n_104), .A2(n_139), .B1(n_1039), .B2(n_1092), .C(n_1093), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_105), .A2(n_250), .B1(n_511), .B2(n_752), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_105), .A2(n_274), .B1(n_482), .B2(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g1411 ( .A(n_106), .Y(n_1411) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_107), .A2(n_324), .B1(n_459), .B2(n_482), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g514 ( .A1(n_107), .A2(n_304), .B1(n_515), .B2(n_518), .C(n_520), .Y(n_514) );
INVx1_ASAP7_75t_L g886 ( .A(n_108), .Y(n_886) );
INVx1_ASAP7_75t_L g1069 ( .A(n_109), .Y(n_1069) );
INVx1_ASAP7_75t_L g382 ( .A(n_110), .Y(n_382) );
INVx1_ASAP7_75t_L g1496 ( .A(n_111), .Y(n_1496) );
INVx1_ASAP7_75t_L g1495 ( .A(n_112), .Y(n_1495) );
AOI22xp33_ASAP7_75t_SL g1358 ( .A1(n_113), .A2(n_303), .B1(n_459), .B2(n_461), .Y(n_1358) );
INVxp67_ASAP7_75t_SL g1379 ( .A(n_113), .Y(n_1379) );
AOI221xp5_ASAP7_75t_L g1502 ( .A1(n_114), .A2(n_301), .B1(n_461), .B2(n_1315), .C(n_1503), .Y(n_1502) );
AOI221xp5_ASAP7_75t_L g1514 ( .A1(n_114), .A2(n_247), .B1(n_540), .B2(n_762), .C(n_1180), .Y(n_1514) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_115), .A2(n_195), .B1(n_785), .B2(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g996 ( .A(n_115), .Y(n_996) );
INVx1_ASAP7_75t_L g714 ( .A(n_116), .Y(n_714) );
OAI22xp33_ASAP7_75t_L g1204 ( .A1(n_117), .A2(n_322), .B1(n_931), .B2(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1238 ( .A(n_117), .Y(n_1238) );
AOI22xp5_ASAP7_75t_L g1632 ( .A1(n_118), .A2(n_348), .B1(n_1613), .B2(n_1625), .Y(n_1632) );
OAI222xp33_ASAP7_75t_L g847 ( .A1(n_119), .A2(n_352), .B1(n_669), .B2(n_671), .C1(n_848), .C2(n_850), .Y(n_847) );
INVx1_ASAP7_75t_L g860 ( .A(n_119), .Y(n_860) );
AOI21xp33_ASAP7_75t_L g1596 ( .A1(n_120), .A2(n_757), .B(n_761), .Y(n_1596) );
INVx1_ASAP7_75t_L g1908 ( .A(n_121), .Y(n_1908) );
OAI221xp5_ASAP7_75t_L g1929 ( .A1(n_121), .A2(n_122), .B1(n_1039), .B2(n_1092), .C(n_1930), .Y(n_1929) );
INVx1_ASAP7_75t_L g1907 ( .A(n_122), .Y(n_1907) );
INVx1_ASAP7_75t_L g837 ( .A(n_123), .Y(n_837) );
OAI211xp5_ASAP7_75t_L g888 ( .A1(n_124), .A2(n_889), .B(n_890), .C(n_891), .Y(n_888) );
INVxp33_ASAP7_75t_SL g911 ( .A(n_124), .Y(n_911) );
OAI22xp33_ASAP7_75t_L g676 ( .A1(n_126), .A2(n_175), .B1(n_677), .B2(n_680), .Y(n_676) );
INVxp67_ASAP7_75t_SL g685 ( .A(n_126), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g1043 ( .A1(n_127), .A2(n_257), .B1(n_1044), .B2(n_1045), .C(n_1047), .Y(n_1043) );
INVx1_ASAP7_75t_L g1211 ( .A(n_128), .Y(n_1211) );
AOI221xp5_ASAP7_75t_L g1233 ( .A1(n_128), .A2(n_294), .B1(n_1044), .B2(n_1234), .C(n_1235), .Y(n_1233) );
INVxp67_ASAP7_75t_SL g1541 ( .A(n_129), .Y(n_1541) );
AOI22xp33_ASAP7_75t_L g1558 ( .A1(n_129), .A2(n_277), .B1(n_1120), .B2(n_1559), .Y(n_1558) );
INVx1_ASAP7_75t_L g1282 ( .A(n_130), .Y(n_1282) );
INVx1_ASAP7_75t_L g1831 ( .A(n_131), .Y(n_1831) );
OAI211xp5_ASAP7_75t_L g1859 ( .A1(n_132), .A2(n_1439), .B(n_1860), .C(n_1863), .Y(n_1859) );
INVx1_ASAP7_75t_L g1890 ( .A(n_132), .Y(n_1890) );
INVx1_ASAP7_75t_L g945 ( .A(n_133), .Y(n_945) );
OAI222xp33_ASAP7_75t_L g987 ( .A1(n_133), .A2(n_221), .B1(n_988), .B2(n_991), .C1(n_997), .C2(n_1004), .Y(n_987) );
INVx1_ASAP7_75t_L g1531 ( .A(n_134), .Y(n_1531) );
OAI22xp33_ASAP7_75t_L g1563 ( .A1(n_134), .A2(n_187), .B1(n_1030), .B2(n_1205), .Y(n_1563) );
XOR2x2_ASAP7_75t_L g1012 ( .A(n_135), .B(n_1013), .Y(n_1012) );
INVxp67_ASAP7_75t_SL g1535 ( .A(n_136), .Y(n_1535) );
AOI22xp33_ASAP7_75t_SL g1560 ( .A1(n_136), .A2(n_213), .B1(n_474), .B2(n_1163), .Y(n_1560) );
AOI22xp33_ASAP7_75t_SL g1078 ( .A1(n_137), .A2(n_143), .B1(n_461), .B2(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1843 ( .A(n_138), .Y(n_1843) );
INVx1_ASAP7_75t_L g1065 ( .A(n_139), .Y(n_1065) );
AOI22xp33_ASAP7_75t_SL g1260 ( .A1(n_140), .A2(n_244), .B1(n_657), .B2(n_963), .Y(n_1260) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_141), .A2(n_372), .B1(n_677), .B2(n_680), .Y(n_697) );
INVxp33_ASAP7_75t_SL g739 ( .A(n_141), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g1913 ( .A1(n_142), .A2(n_184), .B1(n_474), .B2(n_1912), .Y(n_1913) );
INVxp67_ASAP7_75t_SL g1095 ( .A(n_143), .Y(n_1095) );
INVx1_ASAP7_75t_L g1156 ( .A(n_144), .Y(n_1156) );
OAI221xp5_ASAP7_75t_L g1186 ( .A1(n_144), .A2(n_145), .B1(n_1005), .B2(n_1038), .C(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g1157 ( .A(n_145), .Y(n_1157) );
CKINVDCx5p33_ASAP7_75t_R g700 ( .A(n_146), .Y(n_700) );
AOI22xp33_ASAP7_75t_SL g1116 ( .A1(n_147), .A2(n_203), .B1(n_459), .B2(n_482), .Y(n_1116) );
OA21x2_ASAP7_75t_L g1295 ( .A1(n_148), .A2(n_427), .B(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g704 ( .A(n_149), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_149), .A2(n_267), .B1(n_519), .B2(n_722), .C(n_723), .Y(n_721) );
AOI22xp33_ASAP7_75t_SL g1020 ( .A1(n_150), .A2(n_176), .B1(n_461), .B2(n_1021), .Y(n_1020) );
AOI221xp5_ASAP7_75t_L g1053 ( .A1(n_150), .A2(n_204), .B1(n_520), .B2(n_534), .C(n_979), .Y(n_1053) );
OAI22xp33_ASAP7_75t_L g1029 ( .A1(n_151), .A2(n_319), .B1(n_1030), .B2(n_1031), .Y(n_1029) );
INVx1_ASAP7_75t_L g1055 ( .A(n_151), .Y(n_1055) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_152), .A2(n_168), .B1(n_587), .B2(n_610), .C(n_612), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g644 ( .A1(n_152), .A2(n_353), .B1(n_459), .B2(n_482), .C(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_154), .A2(n_340), .B1(n_1118), .B2(n_1120), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_154), .A2(n_235), .B1(n_983), .B2(n_1135), .Y(n_1134) );
OAI22xp33_ASAP7_75t_L g1915 ( .A1(n_155), .A2(n_296), .B1(n_931), .B2(n_1031), .Y(n_1915) );
INVx1_ASAP7_75t_L g1928 ( .A(n_155), .Y(n_1928) );
INVx1_ASAP7_75t_L g969 ( .A(n_156), .Y(n_969) );
INVx1_ASAP7_75t_L g1570 ( .A(n_157), .Y(n_1570) );
OAI221xp5_ASAP7_75t_SL g1593 ( .A1(n_157), .A2(n_278), .B1(n_1004), .B2(n_1092), .C(n_1594), .Y(n_1593) );
CKINVDCx5p33_ASAP7_75t_R g1128 ( .A(n_158), .Y(n_1128) );
OAI22xp33_ASAP7_75t_L g1451 ( .A1(n_159), .A2(n_169), .B1(n_1452), .B2(n_1455), .Y(n_1451) );
OAI22xp33_ASAP7_75t_L g1463 ( .A1(n_159), .A2(n_169), .B1(n_1464), .B2(n_1465), .Y(n_1463) );
INVx1_ASAP7_75t_L g1291 ( .A(n_160), .Y(n_1291) );
INVx1_ASAP7_75t_L g804 ( .A(n_161), .Y(n_804) );
INVx1_ASAP7_75t_L g1838 ( .A(n_162), .Y(n_1838) );
CKINVDCx5p33_ASAP7_75t_R g1034 ( .A(n_164), .Y(n_1034) );
INVx1_ASAP7_75t_L g1442 ( .A(n_165), .Y(n_1442) );
INVx1_ASAP7_75t_L g919 ( .A(n_166), .Y(n_919) );
CKINVDCx5p33_ASAP7_75t_R g1361 ( .A(n_167), .Y(n_1361) );
OAI22xp5_ASAP7_75t_L g1035 ( .A1(n_170), .A2(n_360), .B1(n_554), .B2(n_873), .Y(n_1035) );
INVx1_ASAP7_75t_L g1405 ( .A(n_171), .Y(n_1405) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_172), .A2(n_309), .B1(n_554), .B2(n_873), .Y(n_1062) );
CKINVDCx5p33_ASAP7_75t_R g893 ( .A(n_173), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g1577 ( .A1(n_174), .A2(n_329), .B1(n_468), .B2(n_1578), .Y(n_1577) );
INVxp67_ASAP7_75t_SL g621 ( .A(n_175), .Y(n_621) );
INVxp67_ASAP7_75t_SL g1041 ( .A(n_176), .Y(n_1041) );
OAI22xp5_ASAP7_75t_L g1918 ( .A1(n_177), .A2(n_200), .B1(n_554), .B2(n_873), .Y(n_1918) );
OAI211xp5_ASAP7_75t_L g1920 ( .A1(n_177), .A2(n_1049), .B(n_1921), .C(n_1926), .Y(n_1920) );
INVx1_ASAP7_75t_L g834 ( .A(n_179), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_179), .A2(n_283), .B1(n_753), .B2(n_759), .Y(n_868) );
INVx1_ASAP7_75t_L g569 ( .A(n_180), .Y(n_569) );
INVx1_ASAP7_75t_L g1686 ( .A(n_181), .Y(n_1686) );
INVx1_ASAP7_75t_L g613 ( .A(n_182), .Y(n_613) );
AOI22xp5_ASAP7_75t_SL g1647 ( .A1(n_183), .A2(n_194), .B1(n_1616), .B2(n_1625), .Y(n_1647) );
AOI221xp5_ASAP7_75t_L g1933 ( .A1(n_184), .A2(n_282), .B1(n_1044), .B2(n_1047), .C(n_1934), .Y(n_1933) );
AOI221xp5_ASAP7_75t_L g976 ( .A1(n_185), .A2(n_236), .B1(n_977), .B2(n_979), .C(n_981), .Y(n_976) );
CKINVDCx5p33_ASAP7_75t_R g892 ( .A(n_186), .Y(n_892) );
INVx1_ASAP7_75t_L g1529 ( .A(n_187), .Y(n_1529) );
INVx1_ASAP7_75t_L g903 ( .A(n_188), .Y(n_903) );
AOI22xp33_ASAP7_75t_SL g1072 ( .A1(n_189), .A2(n_288), .B1(n_1073), .B2(n_1074), .Y(n_1072) );
OAI22xp33_ASAP7_75t_L g1867 ( .A1(n_190), .A2(n_357), .B1(n_1868), .B2(n_1869), .Y(n_1867) );
OAI22xp33_ASAP7_75t_L g1877 ( .A1(n_190), .A2(n_357), .B1(n_1878), .B2(n_1880), .Y(n_1877) );
AOI22xp33_ASAP7_75t_SL g1162 ( .A1(n_191), .A2(n_314), .B1(n_643), .B2(n_1163), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_191), .A2(n_240), .B1(n_526), .B2(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g1305 ( .A(n_192), .Y(n_1305) );
AOI221xp5_ASAP7_75t_L g1337 ( .A1(n_192), .A2(n_239), .B1(n_534), .B2(n_540), .C(n_1338), .Y(n_1337) );
OAI211xp5_ASAP7_75t_L g747 ( .A1(n_193), .A2(n_748), .B(n_750), .C(n_763), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_193), .B(n_408), .Y(n_779) );
XNOR2x2_ASAP7_75t_L g1108 ( .A(n_194), .B(n_1109), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_195), .A2(n_297), .B1(n_983), .B2(n_984), .Y(n_982) );
AOI221xp5_ASAP7_75t_L g1505 ( .A1(n_196), .A2(n_247), .B1(n_647), .B2(n_1315), .C(n_1506), .Y(n_1505) );
AOI22xp33_ASAP7_75t_L g1517 ( .A1(n_196), .A2(n_301), .B1(n_526), .B2(n_900), .Y(n_1517) );
INVx1_ASAP7_75t_L g1018 ( .A(n_197), .Y(n_1018) );
OAI221xp5_ASAP7_75t_L g1037 ( .A1(n_197), .A2(n_336), .B1(n_1038), .B2(n_1039), .C(n_1040), .Y(n_1037) );
AOI22xp33_ASAP7_75t_SL g1561 ( .A1(n_198), .A2(n_371), .B1(n_459), .B2(n_1562), .Y(n_1561) );
INVx2_ASAP7_75t_L g1611 ( .A(n_199), .Y(n_1611) );
AND2x2_ASAP7_75t_L g1614 ( .A(n_199), .B(n_1612), .Y(n_1614) );
AND2x2_ASAP7_75t_L g1619 ( .A(n_199), .B(n_318), .Y(n_1619) );
AOI22xp5_ASAP7_75t_SL g1643 ( .A1(n_201), .A2(n_275), .B1(n_1613), .B2(n_1618), .Y(n_1643) );
INVx1_ASAP7_75t_L g1336 ( .A(n_202), .Y(n_1336) );
INVxp67_ASAP7_75t_SL g1142 ( .A(n_203), .Y(n_1142) );
AOI22xp33_ASAP7_75t_SL g1028 ( .A1(n_204), .A2(n_312), .B1(n_482), .B2(n_921), .Y(n_1028) );
INVx1_ASAP7_75t_L g503 ( .A(n_205), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g1615 ( .A1(n_207), .A2(n_344), .B1(n_1616), .B2(n_1618), .Y(n_1615) );
OAI22xp33_ASAP7_75t_L g1125 ( .A1(n_208), .A2(n_285), .B1(n_1030), .B2(n_1031), .Y(n_1125) );
INVx1_ASAP7_75t_L g1138 ( .A(n_208), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_209), .A2(n_359), .B1(n_463), .B2(n_474), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_209), .A2(n_335), .B1(n_523), .B2(n_525), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g1096 ( .A1(n_210), .A2(n_288), .B1(n_755), .B2(n_757), .C(n_1097), .Y(n_1096) );
INVx1_ASAP7_75t_L g1583 ( .A(n_211), .Y(n_1583) );
AOI22xp5_ASAP7_75t_L g1623 ( .A1(n_212), .A2(n_281), .B1(n_1608), .B2(n_1613), .Y(n_1623) );
INVxp67_ASAP7_75t_SL g1542 ( .A(n_213), .Y(n_1542) );
INVx1_ASAP7_75t_L g876 ( .A(n_214), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g1544 ( .A(n_215), .B(n_1038), .Y(n_1544) );
INVx1_ASAP7_75t_L g1554 ( .A(n_215), .Y(n_1554) );
INVx1_ASAP7_75t_L g968 ( .A(n_216), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_217), .A2(n_293), .B1(n_752), .B2(n_753), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g789 ( .A1(n_217), .A2(n_317), .B1(n_459), .B2(n_790), .Y(n_789) );
AOI221xp5_ASAP7_75t_L g1518 ( .A1(n_218), .A2(n_307), .B1(n_540), .B2(n_722), .C(n_1047), .Y(n_1518) );
INVx1_ASAP7_75t_L g1215 ( .A(n_219), .Y(n_1215) );
INVx1_ASAP7_75t_L g1313 ( .A(n_220), .Y(n_1313) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_220), .A2(n_287), .B1(n_753), .B2(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g947 ( .A(n_221), .Y(n_947) );
INVx1_ASAP7_75t_L g1258 ( .A(n_222), .Y(n_1258) );
OAI211xp5_ASAP7_75t_L g1268 ( .A1(n_222), .A2(n_1049), .B(n_1269), .C(n_1275), .Y(n_1268) );
OAI211xp5_ASAP7_75t_L g1438 ( .A1(n_223), .A2(n_1424), .B(n_1439), .C(n_1441), .Y(n_1438) );
INVx1_ASAP7_75t_L g1484 ( .A(n_223), .Y(n_1484) );
AOI22xp5_ASAP7_75t_L g1633 ( .A1(n_224), .A2(n_292), .B1(n_1608), .B2(n_1616), .Y(n_1633) );
XNOR2xp5_ASAP7_75t_L g1900 ( .A(n_225), .B(n_1901), .Y(n_1900) );
INVx1_ASAP7_75t_L g1592 ( .A(n_226), .Y(n_1592) );
CKINVDCx5p33_ASAP7_75t_R g836 ( .A(n_227), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_229), .A2(n_370), .B1(n_1030), .B2(n_1031), .Y(n_1175) );
INVx1_ASAP7_75t_L g1184 ( .A(n_229), .Y(n_1184) );
CKINVDCx5p33_ASAP7_75t_R g773 ( .A(n_230), .Y(n_773) );
INVx2_ASAP7_75t_L g420 ( .A(n_231), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_231), .B(n_418), .Y(n_435) );
INVx1_ASAP7_75t_L g480 ( .A(n_231), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g1276 ( .A(n_232), .Y(n_1276) );
OAI211xp5_ASAP7_75t_L g1231 ( .A1(n_233), .A2(n_1049), .B(n_1232), .C(n_1237), .Y(n_1231) );
INVx1_ASAP7_75t_L g845 ( .A(n_234), .Y(n_845) );
NAND2xp33_ASAP7_75t_SL g869 ( .A(n_234), .B(n_516), .Y(n_869) );
INVx1_ASAP7_75t_L g1410 ( .A(n_237), .Y(n_1410) );
INVx1_ASAP7_75t_L g1310 ( .A(n_239), .Y(n_1310) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_241), .A2(n_323), .B1(n_765), .B2(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g808 ( .A(n_241), .Y(n_808) );
INVx1_ASAP7_75t_L g1217 ( .A(n_242), .Y(n_1217) );
INVx1_ASAP7_75t_L g1281 ( .A(n_243), .Y(n_1281) );
INVx1_ASAP7_75t_L g1285 ( .A(n_244), .Y(n_1285) );
AOI21xp5_ASAP7_75t_L g846 ( .A1(n_245), .A2(n_645), .B(n_656), .Y(n_846) );
INVx1_ASAP7_75t_L g871 ( .A(n_246), .Y(n_871) );
BUFx3_ASAP7_75t_L g412 ( .A(n_248), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g1179 ( .A1(n_249), .A2(n_261), .B1(n_519), .B2(n_520), .C(n_1180), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_250), .A2(n_289), .B1(n_482), .B2(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g1512 ( .A(n_252), .Y(n_1512) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_253), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g701 ( .A(n_254), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g1201 ( .A1(n_255), .A2(n_262), .B1(n_486), .B2(n_1202), .Y(n_1201) );
OAI221xp5_ASAP7_75t_L g1227 ( .A1(n_255), .A2(n_262), .B1(n_1004), .B2(n_1092), .C(n_1228), .Y(n_1227) );
INVx1_ASAP7_75t_L g1866 ( .A(n_256), .Y(n_1866) );
OAI211xp5_ASAP7_75t_L g1883 ( .A1(n_256), .A2(n_1884), .B(n_1886), .C(n_1887), .Y(n_1883) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_257), .A2(n_310), .B1(n_474), .B2(n_651), .Y(n_1026) );
AOI22xp33_ASAP7_75t_SL g1575 ( .A1(n_258), .A2(n_338), .B1(n_964), .B2(n_1266), .Y(n_1575) );
AOI22xp5_ASAP7_75t_L g1607 ( .A1(n_259), .A2(n_290), .B1(n_1608), .B2(n_1613), .Y(n_1607) );
INVx1_ASAP7_75t_L g824 ( .A(n_260), .Y(n_824) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_260), .B(n_677), .Y(n_826) );
AOI22xp33_ASAP7_75t_SL g1161 ( .A1(n_261), .A2(n_306), .B1(n_482), .B2(n_954), .Y(n_1161) );
AOI21xp33_ASAP7_75t_L g906 ( .A1(n_263), .A2(n_519), .B(n_757), .Y(n_906) );
INVx1_ASAP7_75t_L g917 ( .A(n_263), .Y(n_917) );
INVx1_ASAP7_75t_L g1113 ( .A(n_264), .Y(n_1113) );
INVx1_ASAP7_75t_L g497 ( .A(n_265), .Y(n_497) );
INVx1_ASAP7_75t_L g1198 ( .A(n_266), .Y(n_1198) );
AOI21xp33_ASAP7_75t_L g717 ( .A1(n_267), .A2(n_651), .B(n_652), .Y(n_717) );
XOR2x2_ASAP7_75t_L g881 ( .A(n_268), .B(n_882), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_269), .B(n_1152), .Y(n_1151) );
AOI22xp5_ASAP7_75t_L g1169 ( .A1(n_269), .A2(n_1170), .B1(n_1171), .B2(n_1193), .Y(n_1169) );
INVx1_ASAP7_75t_L g1195 ( .A(n_269), .Y(n_1195) );
BUFx3_ASAP7_75t_L g399 ( .A(n_271), .Y(n_399) );
INVx1_ASAP7_75t_L g502 ( .A(n_271), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g1357 ( .A1(n_272), .A2(n_327), .B1(n_959), .B2(n_1024), .Y(n_1357) );
XNOR2x1_ASAP7_75t_L g1492 ( .A(n_273), .B(n_1493), .Y(n_1492) );
NAND2xp5_ASAP7_75t_SL g898 ( .A(n_274), .B(n_519), .Y(n_898) );
INVxp67_ASAP7_75t_SL g1573 ( .A(n_276), .Y(n_1573) );
OAI211xp5_ASAP7_75t_SL g1586 ( .A1(n_276), .A2(n_1132), .B(n_1587), .C(n_1590), .Y(n_1586) );
AOI21xp5_ASAP7_75t_L g1539 ( .A1(n_277), .A2(n_757), .B(n_1086), .Y(n_1539) );
INVx1_ASAP7_75t_L g1571 ( .A(n_278), .Y(n_1571) );
CKINVDCx5p33_ASAP7_75t_R g706 ( .A(n_279), .Y(n_706) );
INVx1_ASAP7_75t_L g1371 ( .A(n_280), .Y(n_1371) );
INVx1_ASAP7_75t_L g843 ( .A(n_283), .Y(n_843) );
INVx1_ASAP7_75t_L g1511 ( .A(n_284), .Y(n_1511) );
INVx1_ASAP7_75t_L g1139 ( .A(n_285), .Y(n_1139) );
CKINVDCx5p33_ASAP7_75t_R g1168 ( .A(n_286), .Y(n_1168) );
NAND2xp33_ASAP7_75t_SL g1307 ( .A(n_287), .B(n_957), .Y(n_1307) );
NAND2xp5_ASAP7_75t_SL g901 ( .A(n_289), .B(n_515), .Y(n_901) );
INVx1_ASAP7_75t_L g688 ( .A(n_291), .Y(n_688) );
AOI22xp33_ASAP7_75t_SL g782 ( .A1(n_293), .A2(n_374), .B1(n_459), .B2(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g1223 ( .A(n_294), .Y(n_1223) );
INVx1_ASAP7_75t_L g415 ( .A(n_295), .Y(n_415) );
INVx1_ASAP7_75t_L g432 ( .A(n_295), .Y(n_432) );
INVx1_ASAP7_75t_L g1927 ( .A(n_296), .Y(n_1927) );
INVx1_ASAP7_75t_L g1333 ( .A(n_299), .Y(n_1333) );
CKINVDCx5p33_ASAP7_75t_R g1061 ( .A(n_300), .Y(n_1061) );
INVx1_ASAP7_75t_L g1836 ( .A(n_302), .Y(n_1836) );
AOI221xp5_ASAP7_75t_L g1366 ( .A1(n_303), .A2(n_333), .B1(n_518), .B2(n_981), .C(n_1367), .Y(n_1366) );
AOI22xp33_ASAP7_75t_L g1369 ( .A1(n_305), .A2(n_327), .B1(n_523), .B2(n_525), .Y(n_1369) );
INVx1_ASAP7_75t_L g1286 ( .A(n_308), .Y(n_1286) );
OAI211xp5_ASAP7_75t_L g1081 ( .A1(n_309), .A2(n_1049), .B(n_1082), .C(n_1090), .Y(n_1081) );
OAI21xp33_ASAP7_75t_L g909 ( .A1(n_311), .A2(n_799), .B(n_910), .Y(n_909) );
INVxp67_ASAP7_75t_SL g1042 ( .A(n_312), .Y(n_1042) );
INVx1_ASAP7_75t_L g614 ( .A(n_313), .Y(n_614) );
AOI21xp33_ASAP7_75t_L g1189 ( .A1(n_314), .A2(n_1047), .B(n_1190), .Y(n_1189) );
CKINVDCx5p33_ASAP7_75t_R g823 ( .A(n_315), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g1499 ( .A(n_316), .Y(n_1499) );
AOI221xp5_ASAP7_75t_SL g760 ( .A1(n_317), .A2(n_374), .B1(n_516), .B2(n_761), .C(n_762), .Y(n_760) );
INVx1_ASAP7_75t_L g1612 ( .A(n_318), .Y(n_1612) );
AND2x2_ASAP7_75t_L g1617 ( .A(n_318), .B(n_1611), .Y(n_1617) );
INVx1_ASAP7_75t_L g1056 ( .A(n_319), .Y(n_1056) );
INVx1_ASAP7_75t_L g1447 ( .A(n_320), .Y(n_1447) );
OAI211xp5_ASAP7_75t_L g1477 ( .A1(n_320), .A2(n_1394), .B(n_1478), .C(n_1481), .Y(n_1477) );
OAI211xp5_ASAP7_75t_SL g1533 ( .A1(n_321), .A2(n_1039), .B(n_1534), .C(n_1540), .Y(n_1533) );
INVx1_ASAP7_75t_L g1553 ( .A(n_321), .Y(n_1553) );
INVx1_ASAP7_75t_L g1239 ( .A(n_322), .Y(n_1239) );
INVx1_ASAP7_75t_L g796 ( .A(n_323), .Y(n_796) );
XNOR2xp5_ASAP7_75t_L g689 ( .A(n_325), .B(n_690), .Y(n_689) );
OAI211xp5_ASAP7_75t_L g1131 ( .A1(n_326), .A2(n_1132), .B(n_1133), .C(n_1137), .Y(n_1131) );
INVx1_ASAP7_75t_L g1391 ( .A(n_328), .Y(n_1391) );
INVx1_ASAP7_75t_L g1595 ( .A(n_329), .Y(n_1595) );
INVxp67_ASAP7_75t_SL g1159 ( .A(n_330), .Y(n_1159) );
OAI211xp5_ASAP7_75t_L g1177 ( .A1(n_330), .A2(n_1049), .B(n_1178), .C(n_1183), .Y(n_1177) );
INVx1_ASAP7_75t_L g1688 ( .A(n_331), .Y(n_1688) );
CKINVDCx16_ASAP7_75t_R g849 ( .A(n_332), .Y(n_849) );
INVx1_ASAP7_75t_L g1017 ( .A(n_336), .Y(n_1017) );
OAI21xp33_ASAP7_75t_L g966 ( .A1(n_337), .A2(n_554), .B(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g692 ( .A(n_339), .Y(n_692) );
OAI21xp5_ASAP7_75t_SL g1519 ( .A1(n_341), .A2(n_1299), .B(n_1520), .Y(n_1519) );
INVx1_ASAP7_75t_L g712 ( .A(n_342), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g1543 ( .A1(n_343), .A2(n_371), .B1(n_520), .B2(n_1147), .C(n_1149), .Y(n_1543) );
XNOR2xp5_ASAP7_75t_L g1820 ( .A(n_344), .B(n_1821), .Y(n_1820) );
AOI22xp33_ASAP7_75t_L g1895 ( .A1(n_344), .A2(n_1896), .B1(n_1899), .B2(n_1935), .Y(n_1895) );
INVx1_ASAP7_75t_L g1840 ( .A(n_345), .Y(n_1840) );
INVx1_ASAP7_75t_L g1404 ( .A(n_346), .Y(n_1404) );
INVx1_ASAP7_75t_L g1392 ( .A(n_347), .Y(n_1392) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_349), .Y(n_444) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_350), .Y(n_395) );
INVx1_ASAP7_75t_L g1548 ( .A(n_351), .Y(n_1548) );
NOR2xp33_ASAP7_75t_R g862 ( .A(n_352), .B(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g819 ( .A(n_354), .Y(n_819) );
INVx1_ASAP7_75t_L g1351 ( .A(n_355), .Y(n_1351) );
OAI221xp5_ASAP7_75t_SL g1375 ( .A1(n_355), .A2(n_375), .B1(n_1004), .B2(n_1092), .C(n_1376), .Y(n_1375) );
INVxp67_ASAP7_75t_SL g631 ( .A(n_356), .Y(n_631) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_356), .A2(n_358), .B1(n_669), .B2(n_671), .C(n_673), .Y(n_668) );
OAI221xp5_ASAP7_75t_L g600 ( .A1(n_358), .A2(n_362), .B1(n_601), .B2(n_606), .C(n_607), .Y(n_600) );
OAI211xp5_ASAP7_75t_L g1048 ( .A1(n_360), .A2(n_1049), .B(n_1050), .C(n_1054), .Y(n_1048) );
XOR2x2_ASAP7_75t_L g1058 ( .A(n_361), .B(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g424 ( .A(n_363), .Y(n_424) );
INVx1_ASAP7_75t_L g438 ( .A(n_363), .Y(n_438) );
INVx2_ASAP7_75t_L g457 ( .A(n_363), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g1917 ( .A(n_365), .Y(n_1917) );
INVx1_ASAP7_75t_L g725 ( .A(n_366), .Y(n_725) );
CKINVDCx5p33_ASAP7_75t_R g1244 ( .A(n_368), .Y(n_1244) );
INVxp67_ASAP7_75t_SL g1145 ( .A(n_369), .Y(n_1145) );
INVx1_ASAP7_75t_L g1185 ( .A(n_370), .Y(n_1185) );
INVxp67_ASAP7_75t_SL g695 ( .A(n_372), .Y(n_695) );
INVx1_ASAP7_75t_L g1255 ( .A(n_373), .Y(n_1255) );
INVx1_ASAP7_75t_L g1352 ( .A(n_375), .Y(n_1352) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_400), .B(n_1599), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_385), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g1894 ( .A(n_379), .B(n_388), .Y(n_1894) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g1898 ( .A(n_381), .B(n_384), .Y(n_1898) );
INVx1_ASAP7_75t_L g1936 ( .A(n_381), .Y(n_1936) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g1938 ( .A(n_384), .B(n_1936), .Y(n_1938) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g1489 ( .A(n_388), .B(n_1490), .Y(n_1489) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g521 ( .A(n_389), .B(n_399), .Y(n_521) );
AND2x4_ASAP7_75t_L g543 ( .A(n_389), .B(n_398), .Y(n_543) );
INVx1_ASAP7_75t_L g1464 ( .A(n_390), .Y(n_1464) );
AND2x4_ASAP7_75t_SL g1893 ( .A(n_390), .B(n_1894), .Y(n_1893) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x6_ASAP7_75t_L g391 ( .A(n_392), .B(n_397), .Y(n_391) );
OR2x6_ASAP7_75t_L g1470 ( .A(n_392), .B(n_1467), .Y(n_1470) );
INVx1_ASAP7_75t_L g1857 ( .A(n_392), .Y(n_1857) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g589 ( .A(n_393), .Y(n_589) );
BUFx4f_ASAP7_75t_L g766 ( .A(n_393), .Y(n_766) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx2_ASAP7_75t_L g442 ( .A(n_395), .Y(n_442) );
AND2x2_ASAP7_75t_L g507 ( .A(n_395), .B(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g513 ( .A(n_395), .Y(n_513) );
AND2x2_ASAP7_75t_L g517 ( .A(n_395), .B(n_396), .Y(n_517) );
INVx1_ASAP7_75t_L g558 ( .A(n_395), .Y(n_558) );
NAND2x1_ASAP7_75t_L g597 ( .A(n_395), .B(n_396), .Y(n_597) );
INVx1_ASAP7_75t_L g443 ( .A(n_396), .Y(n_443) );
INVx2_ASAP7_75t_L g508 ( .A(n_396), .Y(n_508) );
AND2x2_ASAP7_75t_L g512 ( .A(n_396), .B(n_513), .Y(n_512) );
BUFx2_ASAP7_75t_L g548 ( .A(n_396), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_396), .B(n_513), .Y(n_586) );
OR2x2_ASAP7_75t_L g593 ( .A(n_396), .B(n_442), .Y(n_593) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g1480 ( .A(n_398), .Y(n_1480) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_L g1476 ( .A(n_399), .Y(n_1476) );
AND2x4_ASAP7_75t_L g1487 ( .A(n_399), .B(n_557), .Y(n_1487) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_1101), .B2(n_1102), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
XNOR2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_571), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_568), .B1(n_569), .B2(n_570), .Y(n_404) );
INVx1_ASAP7_75t_L g570 ( .A(n_405), .Y(n_570) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_494), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_425), .B1(n_426), .B2(n_444), .C(n_445), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g1296 ( .A1(n_407), .A2(n_1297), .B1(n_1298), .B2(n_1300), .Y(n_1296) );
AOI221xp5_ASAP7_75t_L g1494 ( .A1(n_407), .A2(n_426), .B1(n_1495), .B2(n_1496), .C(n_1497), .Y(n_1494) );
INVx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx5_ASAP7_75t_L g937 ( .A(n_408), .Y(n_937) );
OR2x6_ASAP7_75t_L g408 ( .A(n_409), .B(n_421), .Y(n_408) );
INVx2_ASAP7_75t_L g667 ( .A(n_409), .Y(n_667) );
OR2x2_ASAP7_75t_L g873 ( .A(n_409), .B(n_421), .Y(n_873) );
NAND2x1p5_ASAP7_75t_L g409 ( .A(n_410), .B(n_416), .Y(n_409) );
INVx8_ASAP7_75t_L g460 ( .A(n_410), .Y(n_460) );
BUFx3_ASAP7_75t_L g656 ( .A(n_410), .Y(n_656) );
AND2x2_ASAP7_75t_L g660 ( .A(n_410), .B(n_661), .Y(n_660) );
BUFx3_ASAP7_75t_L g921 ( .A(n_410), .Y(n_921) );
HB1xp67_ASAP7_75t_L g927 ( .A(n_410), .Y(n_927) );
AND2x4_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
AND2x4_ASAP7_75t_L g466 ( .A(n_411), .B(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_412), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g449 ( .A(n_412), .B(n_450), .Y(n_449) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_412), .Y(n_471) );
OR2x2_ASAP7_75t_L g830 ( .A(n_412), .B(n_414), .Y(n_830) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g467 ( .A(n_415), .Y(n_467) );
AND2x4_ASAP7_75t_L g451 ( .A(n_416), .B(n_437), .Y(n_451) );
AND2x6_ASAP7_75t_L g670 ( .A(n_416), .B(n_487), .Y(n_670) );
AND2x2_ASAP7_75t_L g672 ( .A(n_416), .B(n_493), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_416), .Y(n_675) );
AND2x4_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
NAND3x1_ASAP7_75t_L g478 ( .A(n_417), .B(n_479), .C(n_480), .Y(n_478) );
NAND2x1p5_ASAP7_75t_L g645 ( .A(n_417), .B(n_480), .Y(n_645) );
INVx1_ASAP7_75t_L g1434 ( .A(n_417), .Y(n_1434) );
OR2x6_ASAP7_75t_L g1437 ( .A(n_417), .B(n_1312), .Y(n_1437) );
AND2x4_ASAP7_75t_L g1440 ( .A(n_417), .B(n_449), .Y(n_1440) );
OR2x4_ASAP7_75t_L g1454 ( .A(n_417), .B(n_830), .Y(n_1454) );
INVx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx3_ASAP7_75t_L g455 ( .A(n_418), .Y(n_455) );
NAND2xp33_ASAP7_75t_SL g653 ( .A(n_418), .B(n_420), .Y(n_653) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND3x4_ASAP7_75t_L g454 ( .A(n_420), .B(n_455), .C(n_456), .Y(n_454) );
AND2x2_ASAP7_75t_L g838 ( .A(n_420), .B(n_455), .Y(n_838) );
HB1xp67_ASAP7_75t_L g1459 ( .A(n_420), .Y(n_1459) );
INVxp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g555 ( .A(n_422), .B(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g606 ( .A(n_422), .B(n_556), .Y(n_606) );
INVx1_ASAP7_75t_L g637 ( .A(n_422), .Y(n_637) );
INVx1_ASAP7_75t_L g1490 ( .A(n_422), .Y(n_1490) );
BUFx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g434 ( .A(n_423), .Y(n_434) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g509 ( .A1(n_425), .A2(n_510), .B1(n_514), .B2(n_522), .C(n_527), .Y(n_509) );
AOI211x1_ASAP7_75t_L g940 ( .A1(n_426), .A2(n_941), .B(n_942), .C(n_966), .Y(n_940) );
AOI21xp33_ASAP7_75t_SL g1033 ( .A1(n_426), .A2(n_1034), .B(n_1035), .Y(n_1033) );
AOI21xp5_ASAP7_75t_L g1060 ( .A1(n_426), .A2(n_1061), .B(n_1062), .Y(n_1060) );
AOI21xp33_ASAP7_75t_SL g1127 ( .A1(n_426), .A2(n_1128), .B(n_1129), .Y(n_1127) );
NAND2xp33_ASAP7_75t_L g1167 ( .A(n_426), .B(n_1168), .Y(n_1167) );
AOI21xp33_ASAP7_75t_L g1243 ( .A1(n_426), .A2(n_1244), .B(n_1245), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_426), .B(n_1290), .Y(n_1289) );
AOI21xp5_ASAP7_75t_L g1360 ( .A1(n_426), .A2(n_1361), .B(n_1362), .Y(n_1360) );
AOI21xp33_ASAP7_75t_SL g1547 ( .A1(n_426), .A2(n_1548), .B(n_1549), .Y(n_1547) );
AOI211x1_ASAP7_75t_L g1566 ( .A1(n_426), .A2(n_1567), .B(n_1568), .C(n_1581), .Y(n_1566) );
AOI21xp33_ASAP7_75t_SL g1916 ( .A1(n_426), .A2(n_1917), .B(n_1918), .Y(n_1916) );
INVx8_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_428), .B(n_436), .Y(n_427) );
INVx1_ASAP7_75t_L g809 ( .A(n_428), .Y(n_809) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_433), .Y(n_428) );
BUFx3_ASAP7_75t_L g705 ( .A(n_429), .Y(n_705) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx6f_ASAP7_75t_L g833 ( .A(n_430), .Y(n_833) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g1312 ( .A(n_431), .Y(n_1312) );
INVx2_ASAP7_75t_L g450 ( .A(n_432), .Y(n_450) );
INVx1_ASAP7_75t_L g562 ( .A(n_432), .Y(n_562) );
OR2x2_ASAP7_75t_L g559 ( .A(n_433), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g566 ( .A(n_433), .Y(n_566) );
INVx1_ASAP7_75t_L g802 ( .A(n_433), .Y(n_802) );
OR2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
AND2x2_ASAP7_75t_SL g599 ( .A(n_434), .B(n_521), .Y(n_599) );
INVx1_ASAP7_75t_L g733 ( .A(n_434), .Y(n_733) );
OR2x2_ASAP7_75t_L g915 ( .A(n_434), .B(n_653), .Y(n_915) );
HB1xp67_ASAP7_75t_L g1461 ( .A(n_434), .Y(n_1461) );
INVx1_ASAP7_75t_L g661 ( .A(n_435), .Y(n_661) );
INVx1_ASAP7_75t_L g679 ( .A(n_435), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_436), .B(n_878), .Y(n_877) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .Y(n_436) );
INVx1_ASAP7_75t_L g619 ( .A(n_437), .Y(n_619) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g479 ( .A(n_438), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_438), .B(n_501), .Y(n_624) );
INVx1_ASAP7_75t_L g620 ( .A(n_439), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
AND2x6_ASAP7_75t_L g527 ( .A(n_440), .B(n_516), .Y(n_527) );
AND2x2_ASAP7_75t_L g546 ( .A(n_440), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_440), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_440), .B(n_457), .Y(n_603) );
INVx1_ASAP7_75t_L g775 ( .A(n_440), .Y(n_775) );
AND2x2_ASAP7_75t_L g500 ( .A(n_441), .B(n_501), .Y(n_500) );
INVx3_ASAP7_75t_L g524 ( .A(n_441), .Y(n_524) );
BUFx6f_ASAP7_75t_L g752 ( .A(n_441), .Y(n_752) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_442), .Y(n_772) );
NAND3xp33_ASAP7_75t_SL g445 ( .A(n_446), .B(n_452), .C(n_483), .Y(n_445) );
AND5x1_ASAP7_75t_L g882 ( .A(n_446), .B(n_883), .C(n_912), .D(n_928), .E(n_935), .Y(n_882) );
INVx2_ASAP7_75t_SL g1032 ( .A(n_446), .Y(n_1032) );
NAND4xp75_ASAP7_75t_L g1059 ( .A(n_446), .B(n_1060), .C(n_1063), .D(n_1080), .Y(n_1059) );
AND4x1_ASAP7_75t_L g1253 ( .A(n_446), .B(n_1254), .C(n_1257), .D(n_1259), .Y(n_1253) );
NAND3xp33_ASAP7_75t_SL g1497 ( .A(n_446), .B(n_1498), .C(n_1501), .Y(n_1497) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g793 ( .A1(n_447), .A2(n_770), .B1(n_794), .B2(n_795), .C(n_796), .Y(n_793) );
INVx3_ASAP7_75t_L g951 ( .A(n_447), .Y(n_951) );
NOR3xp33_ASAP7_75t_SL g1301 ( .A(n_447), .B(n_1302), .C(n_1316), .Y(n_1301) );
AND2x4_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .Y(n_447) );
BUFx2_ASAP7_75t_L g1355 ( .A(n_448), .Y(n_1355) );
BUFx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx2_ASAP7_75t_L g461 ( .A(n_449), .Y(n_461) );
BUFx3_ASAP7_75t_L g482 ( .A(n_449), .Y(n_482) );
INVx2_ASAP7_75t_L g648 ( .A(n_449), .Y(n_648) );
AND2x2_ASAP7_75t_L g663 ( .A(n_449), .B(n_661), .Y(n_663) );
BUFx2_ASAP7_75t_L g783 ( .A(n_449), .Y(n_783) );
BUFx2_ASAP7_75t_L g1123 ( .A(n_449), .Y(n_1123) );
BUFx2_ASAP7_75t_L g1557 ( .A(n_449), .Y(n_1557) );
INVx1_ASAP7_75t_L g472 ( .A(n_450), .Y(n_472) );
NAND2x1_ASAP7_75t_L g486 ( .A(n_451), .B(n_487), .Y(n_486) );
AND2x4_ASAP7_75t_L g490 ( .A(n_451), .B(n_491), .Y(n_490) );
AND2x4_ASAP7_75t_SL g794 ( .A(n_451), .B(n_487), .Y(n_794) );
AND2x4_ASAP7_75t_SL g795 ( .A(n_451), .B(n_491), .Y(n_795) );
AND2x2_ASAP7_75t_L g946 ( .A(n_451), .B(n_487), .Y(n_946) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_451), .B(n_487), .Y(n_1318) );
AOI33xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_458), .A3(n_462), .B1(n_473), .B2(n_475), .B3(n_481), .Y(n_452) );
AOI33xp33_ASAP7_75t_L g952 ( .A1(n_453), .A2(n_953), .A3(n_956), .B1(n_958), .B2(n_960), .B3(n_962), .Y(n_952) );
AOI33xp33_ASAP7_75t_L g1070 ( .A1(n_453), .A2(n_1027), .A3(n_1071), .B1(n_1072), .B2(n_1075), .B3(n_1078), .Y(n_1070) );
AOI33xp33_ASAP7_75t_L g1259 ( .A1(n_453), .A2(n_1027), .A3(n_1260), .B1(n_1261), .B2(n_1264), .B3(n_1265), .Y(n_1259) );
AOI33xp33_ASAP7_75t_L g1353 ( .A1(n_453), .A2(n_475), .A3(n_1354), .B1(n_1356), .B2(n_1357), .B3(n_1358), .Y(n_1353) );
AOI33xp33_ASAP7_75t_L g1574 ( .A1(n_453), .A2(n_477), .A3(n_1575), .B1(n_1576), .B2(n_1577), .B3(n_1580), .Y(n_1574) );
BUFx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI33xp33_ASAP7_75t_L g781 ( .A1(n_454), .A2(n_782), .A3(n_784), .B1(n_787), .B2(n_789), .B3(n_791), .Y(n_781) );
AOI33xp33_ASAP7_75t_L g1019 ( .A1(n_454), .A2(n_1020), .A3(n_1023), .B1(n_1026), .B2(n_1027), .B3(n_1028), .Y(n_1019) );
AOI33xp33_ASAP7_75t_L g1115 ( .A1(n_454), .A2(n_1116), .A3(n_1117), .B1(n_1121), .B2(n_1122), .B3(n_1124), .Y(n_1115) );
AOI33xp33_ASAP7_75t_L g1160 ( .A1(n_454), .A2(n_1027), .A3(n_1161), .B1(n_1162), .B2(n_1165), .B3(n_1166), .Y(n_1160) );
INVx1_ASAP7_75t_L g1506 ( .A(n_454), .Y(n_1506) );
AOI33xp33_ASAP7_75t_L g1555 ( .A1(n_454), .A2(n_1124), .A3(n_1556), .B1(n_1558), .B2(n_1560), .B3(n_1561), .Y(n_1555) );
AOI33xp33_ASAP7_75t_L g1909 ( .A1(n_454), .A2(n_1124), .A3(n_1910), .B1(n_1911), .B2(n_1913), .B3(n_1914), .Y(n_1909) );
INVx3_ASAP7_75t_L g1445 ( .A(n_455), .Y(n_1445) );
INVx1_ASAP7_75t_L g683 ( .A(n_456), .Y(n_683) );
OAI31xp33_ASAP7_75t_SL g696 ( .A1(n_456), .A2(n_697), .A3(n_698), .B(n_702), .Y(n_696) );
OAI31xp33_ASAP7_75t_L g825 ( .A1(n_456), .A2(n_826), .A3(n_827), .B(n_847), .Y(n_825) );
INVx2_ASAP7_75t_SL g1057 ( .A(n_456), .Y(n_1057) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g552 ( .A(n_457), .Y(n_552) );
BUFx2_ASAP7_75t_L g1266 ( .A(n_459), .Y(n_1266) );
INVx8_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g565 ( .A(n_460), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g708 ( .A(n_460), .Y(n_708) );
INVx3_ASAP7_75t_L g963 ( .A(n_460), .Y(n_963) );
INVx2_ASAP7_75t_L g1315 ( .A(n_460), .Y(n_1315) );
INVx1_ASAP7_75t_L g965 ( .A(n_461), .Y(n_965) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g1218 ( .A1(n_464), .A2(n_842), .B1(n_1219), .B2(n_1220), .Y(n_1218) );
INVx2_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
AND2x4_ASAP7_75t_L g567 ( .A(n_465), .B(n_566), .Y(n_567) );
HB1xp67_ASAP7_75t_L g1073 ( .A(n_465), .Y(n_1073) );
INVx3_ASAP7_75t_L g1579 ( .A(n_465), .Y(n_1579) );
INVx3_ASAP7_75t_L g1837 ( .A(n_465), .Y(n_1837) );
BUFx8_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g642 ( .A(n_466), .Y(n_642) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_466), .Y(n_651) );
BUFx6f_ASAP7_75t_L g786 ( .A(n_466), .Y(n_786) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g957 ( .A(n_469), .Y(n_957) );
INVx2_ASAP7_75t_R g1120 ( .A(n_469), .Y(n_1120) );
INVx5_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx3_ASAP7_75t_L g474 ( .A(n_470), .Y(n_474) );
BUFx2_ASAP7_75t_L g643 ( .A(n_470), .Y(n_643) );
BUFx12f_ASAP7_75t_L g657 ( .A(n_470), .Y(n_657) );
AND2x4_ASAP7_75t_L g681 ( .A(n_470), .B(n_679), .Y(n_681) );
BUFx3_ASAP7_75t_L g1074 ( .A(n_470), .Y(n_1074) );
AND2x4_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
INVx2_ASAP7_75t_L g488 ( .A(n_471), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g561 ( .A(n_471), .B(n_562), .Y(n_561) );
BUFx2_ASAP7_75t_L g1446 ( .A(n_471), .Y(n_1446) );
INVx1_ASAP7_75t_L g493 ( .A(n_472), .Y(n_493) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g922 ( .A(n_477), .Y(n_922) );
INVx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx3_ASAP7_75t_L g961 ( .A(n_478), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B1(n_489), .B2(n_490), .Y(n_483) );
AOI222xp33_ASAP7_75t_L g528 ( .A1(n_484), .A2(n_489), .B1(n_529), .B2(n_531), .C1(n_533), .C2(n_544), .Y(n_528) );
AOI221x1_ASAP7_75t_L g912 ( .A1(n_485), .A2(n_490), .B1(n_886), .B2(n_892), .C(n_913), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_485), .A2(n_490), .B1(n_1017), .B2(n_1018), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_485), .A2(n_490), .B1(n_1065), .B2(n_1066), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_485), .A2(n_490), .B1(n_1113), .B2(n_1114), .Y(n_1112) );
AOI22xp5_ASAP7_75t_L g1155 ( .A1(n_485), .A2(n_490), .B1(n_1156), .B2(n_1157), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_485), .A2(n_1203), .B1(n_1255), .B2(n_1256), .Y(n_1254) );
AOI22xp33_ASAP7_75t_L g1906 ( .A1(n_485), .A2(n_490), .B1(n_1907), .B2(n_1908), .Y(n_1906) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AO22x1_ASAP7_75t_L g944 ( .A1(n_490), .A2(n_945), .B1(n_946), .B2(n_947), .Y(n_944) );
HB1xp67_ASAP7_75t_L g1203 ( .A(n_490), .Y(n_1203) );
AOI22xp33_ASAP7_75t_L g1350 ( .A1(n_490), .A2(n_946), .B1(n_1351), .B2(n_1352), .Y(n_1350) );
AOI22xp33_ASAP7_75t_L g1552 ( .A1(n_490), .A2(n_1318), .B1(n_1553), .B2(n_1554), .Y(n_1552) );
AOI22xp5_ASAP7_75t_L g1569 ( .A1(n_490), .A2(n_1318), .B1(n_1570), .B2(n_1571), .Y(n_1569) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_549), .B(n_553), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_509), .C(n_528), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B1(n_503), .B2(n_504), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_497), .A2(n_503), .B1(n_564), .B2(n_567), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_498), .A2(n_1371), .B1(n_1372), .B2(n_1373), .Y(n_1370) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_499), .A2(n_505), .B1(n_1068), .B2(n_1069), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_499), .A2(n_505), .B1(n_1184), .B2(n_1185), .Y(n_1183) );
AOI22xp5_ASAP7_75t_L g1327 ( .A1(n_499), .A2(n_505), .B1(n_1328), .B2(n_1329), .Y(n_1327) );
AOI22xp5_ASAP7_75t_L g1510 ( .A1(n_499), .A2(n_505), .B1(n_1511), .B2(n_1512), .Y(n_1510) );
AOI22xp33_ASAP7_75t_L g1530 ( .A1(n_499), .A2(n_510), .B1(n_1531), .B2(n_1532), .Y(n_1530) );
AOI22xp33_ASAP7_75t_L g1590 ( .A1(n_499), .A2(n_504), .B1(n_1591), .B2(n_1592), .Y(n_1590) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x4_ASAP7_75t_L g636 ( .A(n_500), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g974 ( .A(n_500), .Y(n_974) );
AND2x4_ASAP7_75t_L g505 ( .A(n_501), .B(n_506), .Y(n_505) );
AND2x4_ASAP7_75t_L g510 ( .A(n_501), .B(n_511), .Y(n_510) );
AND2x4_ASAP7_75t_SL g530 ( .A(n_501), .B(n_516), .Y(n_530) );
AND2x2_ASAP7_75t_L g687 ( .A(n_501), .B(n_506), .Y(n_687) );
AND2x2_ASAP7_75t_L g749 ( .A(n_501), .B(n_625), .Y(n_749) );
BUFx2_ASAP7_75t_L g776 ( .A(n_501), .Y(n_776) );
HB1xp67_ASAP7_75t_L g1467 ( .A(n_502), .Y(n_1467) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_504), .A2(n_973), .B1(n_1055), .B2(n_1056), .Y(n_1054) );
AOI22xp5_ASAP7_75t_L g1137 ( .A1(n_504), .A2(n_973), .B1(n_1138), .B2(n_1139), .Y(n_1137) );
AOI21xp5_ASAP7_75t_L g1528 ( .A1(n_504), .A2(n_527), .B(n_1529), .Y(n_1528) );
AOI22xp33_ASAP7_75t_L g1926 ( .A1(n_504), .A2(n_973), .B1(n_1927), .B2(n_1928), .Y(n_1926) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_505), .A2(n_968), .B1(n_969), .B2(n_973), .Y(n_972) );
HB1xp67_ASAP7_75t_L g1240 ( .A(n_505), .Y(n_1240) );
INVx1_ASAP7_75t_L g1374 ( .A(n_505), .Y(n_1374) );
INVx2_ASAP7_75t_L g541 ( .A(n_506), .Y(n_541) );
BUFx6f_ASAP7_75t_L g980 ( .A(n_506), .Y(n_980) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
BUFx3_ASAP7_75t_L g519 ( .A(n_507), .Y(n_519) );
INVx2_ASAP7_75t_L g756 ( .A(n_507), .Y(n_756) );
AND2x4_ASAP7_75t_L g1466 ( .A(n_507), .B(n_1467), .Y(n_1466) );
NAND2xp5_ASAP7_75t_R g986 ( .A(n_510), .B(n_950), .Y(n_986) );
INVx2_ASAP7_75t_SL g1049 ( .A(n_510), .Y(n_1049) );
INVx3_ASAP7_75t_L g1132 ( .A(n_510), .Y(n_1132) );
BUFx2_ASAP7_75t_L g1135 ( .A(n_511), .Y(n_1135) );
INVx1_ASAP7_75t_L g1274 ( .A(n_511), .Y(n_1274) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx3_ASAP7_75t_L g526 ( .A(n_512), .Y(n_526) );
INVx2_ASAP7_75t_L g626 ( .A(n_512), .Y(n_626) );
BUFx3_ASAP7_75t_L g753 ( .A(n_512), .Y(n_753) );
BUFx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx3_ASAP7_75t_L g722 ( .A(n_516), .Y(n_722) );
BUFx3_ASAP7_75t_L g1044 ( .A(n_516), .Y(n_1044) );
INVx1_ASAP7_75t_L g1085 ( .A(n_516), .Y(n_1085) );
BUFx3_ASAP7_75t_L g1149 ( .A(n_516), .Y(n_1149) );
BUFx6f_ASAP7_75t_L g1180 ( .A(n_516), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_516), .B(n_1480), .Y(n_1479) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g537 ( .A(n_517), .Y(n_537) );
BUFx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g1191 ( .A(n_519), .Y(n_1191) );
HB1xp67_ASAP7_75t_SL g1235 ( .A(n_520), .Y(n_1235) );
INVx4_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x4_ASAP7_75t_L g731 ( .A(n_521), .B(n_732), .Y(n_731) );
INVx4_ASAP7_75t_L g762 ( .A(n_521), .Y(n_762) );
NAND4xp25_ASAP7_75t_L g897 ( .A(n_521), .B(n_898), .C(n_899), .D(n_901), .Y(n_897) );
INVx1_ASAP7_75t_SL g981 ( .A(n_521), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g1408 ( .A(n_521), .B(n_732), .Y(n_1408) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_SL g532 ( .A(n_524), .Y(n_532) );
INVx2_ASAP7_75t_L g759 ( .A(n_524), .Y(n_759) );
INVx1_ASAP7_75t_L g900 ( .A(n_524), .Y(n_900) );
INVx2_ASAP7_75t_L g983 ( .A(n_524), .Y(n_983) );
INVx1_ASAP7_75t_L g1052 ( .A(n_524), .Y(n_1052) );
BUFx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_SL g985 ( .A(n_526), .Y(n_985) );
AOI21xp5_ASAP7_75t_L g975 ( .A1(n_527), .A2(n_976), .B(n_982), .Y(n_975) );
AOI21xp5_ASAP7_75t_L g1050 ( .A1(n_527), .A2(n_1051), .B(n_1053), .Y(n_1050) );
AOI21xp5_ASAP7_75t_SL g1082 ( .A1(n_527), .A2(n_1083), .B(n_1088), .Y(n_1082) );
AOI21xp5_ASAP7_75t_L g1133 ( .A1(n_527), .A2(n_1134), .B(n_1136), .Y(n_1133) );
AOI21xp5_ASAP7_75t_L g1178 ( .A1(n_527), .A2(n_1179), .B(n_1181), .Y(n_1178) );
AOI21xp5_ASAP7_75t_L g1232 ( .A1(n_527), .A2(n_1233), .B(n_1236), .Y(n_1232) );
AOI21xp5_ASAP7_75t_L g1269 ( .A1(n_527), .A2(n_1270), .B(n_1271), .Y(n_1269) );
AOI221xp5_ASAP7_75t_L g1322 ( .A1(n_527), .A2(n_749), .B1(n_1300), .B2(n_1323), .C(n_1324), .Y(n_1322) );
AOI21xp5_ASAP7_75t_L g1365 ( .A1(n_527), .A2(n_1366), .B(n_1369), .Y(n_1365) );
AOI221xp5_ASAP7_75t_L g1513 ( .A1(n_527), .A2(n_749), .B1(n_1495), .B2(n_1514), .C(n_1515), .Y(n_1513) );
AOI21xp5_ASAP7_75t_L g1587 ( .A1(n_527), .A2(n_1588), .B(n_1589), .Y(n_1587) );
AOI21xp5_ASAP7_75t_SL g1921 ( .A1(n_527), .A2(n_1922), .B(n_1925), .Y(n_1921) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_529), .B(n_886), .Y(n_885) );
AOI222xp33_ASAP7_75t_L g1516 ( .A1(n_529), .A2(n_546), .B1(n_1499), .B2(n_1500), .C1(n_1517), .C2(n_1518), .Y(n_1516) );
BUFx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g990 ( .A(n_530), .Y(n_990) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx2_ASAP7_75t_L g978 ( .A(n_537), .Y(n_978) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
HB1xp67_ASAP7_75t_L g1924 ( .A(n_540), .Y(n_1924) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g1046 ( .A(n_541), .Y(n_1046) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx3_ASAP7_75t_L g757 ( .A(n_543), .Y(n_757) );
OAI221xp5_ASAP7_75t_L g991 ( .A1(n_543), .A2(n_595), .B1(n_992), .B2(n_993), .C(n_996), .Y(n_991) );
INVx2_ASAP7_75t_L g1047 ( .A(n_543), .Y(n_1047) );
INVx2_ASAP7_75t_L g1338 ( .A(n_543), .Y(n_1338) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_547), .A2(n_770), .B1(n_771), .B2(n_773), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_547), .A2(n_771), .B1(n_892), .B2(n_893), .Y(n_891) );
BUFx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g605 ( .A(n_548), .Y(n_605) );
INVx1_ASAP7_75t_L g1007 ( .A(n_548), .Y(n_1007) );
AND2x4_ASAP7_75t_L g1483 ( .A(n_548), .B(n_1476), .Y(n_1483) );
OAI21xp5_ASAP7_75t_L g970 ( .A1(n_549), .A2(n_971), .B(n_987), .Y(n_970) );
OAI21xp5_ASAP7_75t_L g1176 ( .A1(n_549), .A2(n_1177), .B(n_1186), .Y(n_1176) );
AOI21xp5_ASAP7_75t_L g1508 ( .A1(n_549), .A2(n_1509), .B(n_1519), .Y(n_1508) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g1339 ( .A(n_550), .Y(n_1339) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_551), .B(n_681), .Y(n_878) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g615 ( .A(n_552), .B(n_616), .Y(n_615) );
OR2x6_ASAP7_75t_L g792 ( .A(n_552), .B(n_645), .Y(n_792) );
OR2x2_ASAP7_75t_L g1503 ( .A(n_552), .B(n_645), .Y(n_1503) );
INVx2_ASAP7_75t_L g1173 ( .A(n_554), .Y(n_1173) );
HB1xp67_ASAP7_75t_L g1246 ( .A(n_554), .Y(n_1246) );
AND2x4_ASAP7_75t_L g554 ( .A(n_555), .B(n_559), .Y(n_554) );
INVx2_ASAP7_75t_SL g737 ( .A(n_555), .Y(n_737) );
AND2x4_ASAP7_75t_L g1299 ( .A(n_555), .B(n_559), .Y(n_1299) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g806 ( .A(n_559), .Y(n_806) );
INVx3_ASAP7_75t_L g716 ( .A(n_560), .Y(n_716) );
BUFx6f_ASAP7_75t_L g1419 ( .A(n_560), .Y(n_1419) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
BUFx2_ASAP7_75t_L g674 ( .A(n_561), .Y(n_674) );
BUFx3_ASAP7_75t_L g1425 ( .A(n_561), .Y(n_1425) );
BUFx2_ASAP7_75t_L g1450 ( .A(n_562), .Y(n_1450) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_564), .A2(n_567), .B1(n_968), .B2(n_969), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g1288 ( .A1(n_564), .A2(n_567), .B1(n_1276), .B2(n_1277), .Y(n_1288) );
AOI22xp5_ASAP7_75t_L g1340 ( .A1(n_564), .A2(n_1328), .B1(n_1329), .B2(n_1341), .Y(n_1340) );
AND2x4_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
AND2x4_ASAP7_75t_L g807 ( .A(n_565), .B(n_566), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g848 ( .A1(n_565), .A2(n_790), .B1(n_823), .B2(n_849), .Y(n_848) );
INVx2_ASAP7_75t_L g1031 ( .A(n_567), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_567), .A2(n_807), .B1(n_1068), .B2(n_1069), .Y(n_1067) );
INVx2_ASAP7_75t_L g1205 ( .A(n_567), .Y(n_1205) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_569), .Y(n_568) );
AO22x2_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_1011), .B1(n_1099), .B2(n_1100), .Y(n_571) );
XOR2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_741), .Y(n_572) );
XNOR2x1_ASAP7_75t_L g1100 ( .A(n_573), .B(n_741), .Y(n_1100) );
BUFx2_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
INVxp67_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
XNOR2x1_ASAP7_75t_L g575 ( .A(n_576), .B(n_689), .Y(n_575) );
XNOR2x1_ASAP7_75t_L g576 ( .A(n_577), .B(n_688), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_638), .Y(n_577) );
NAND3xp33_ASAP7_75t_SL g578 ( .A(n_579), .B(n_617), .C(n_632), .Y(n_578) );
AOI211xp5_ASAP7_75t_SL g579 ( .A1(n_580), .A2(n_590), .B(n_600), .C(n_609), .Y(n_579) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OAI221xp5_ASAP7_75t_L g1093 ( .A1(n_582), .A2(n_588), .B1(n_1094), .B2(n_1095), .C(n_1096), .Y(n_1093) );
BUFx2_ASAP7_75t_L g1229 ( .A(n_582), .Y(n_1229) );
OAI221xp5_ASAP7_75t_L g1930 ( .A1(n_582), .A2(n_999), .B1(n_1931), .B2(n_1932), .C(n_1933), .Y(n_1930) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g726 ( .A(n_584), .Y(n_726) );
INVx4_ASAP7_75t_L g896 ( .A(n_584), .Y(n_896) );
BUFx6f_ASAP7_75t_L g1003 ( .A(n_584), .Y(n_1003) );
INVx2_ASAP7_75t_SL g1144 ( .A(n_584), .Y(n_1144) );
INVx1_ASAP7_75t_L g1335 ( .A(n_584), .Y(n_1335) );
INVx1_ASAP7_75t_L g1378 ( .A(n_584), .Y(n_1378) );
INVx8_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
BUFx2_ASAP7_75t_L g611 ( .A(n_585), .Y(n_611) );
OR2x2_ASAP7_75t_L g1475 ( .A(n_585), .B(n_1476), .Y(n_1475) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI221xp5_ASAP7_75t_L g1141 ( .A1(n_588), .A2(n_1142), .B1(n_1143), .B2(n_1145), .C(n_1146), .Y(n_1141) );
OAI221xp5_ASAP7_75t_SL g1228 ( .A1(n_588), .A2(n_1215), .B1(n_1222), .B2(n_1229), .C(n_1230), .Y(n_1228) );
OAI22xp5_ASAP7_75t_L g1284 ( .A1(n_588), .A2(n_1229), .B1(n_1285), .B2(n_1286), .Y(n_1284) );
OAI221xp5_ASAP7_75t_L g1540 ( .A1(n_588), .A2(n_1143), .B1(n_1541), .B2(n_1542), .C(n_1543), .Y(n_1540) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_589), .A2(n_724), .B1(n_725), .B2(n_726), .Y(n_723) );
OAI22x1_ASAP7_75t_SL g729 ( .A1(n_589), .A2(n_706), .B1(n_726), .B2(n_730), .Y(n_729) );
BUFx3_ASAP7_75t_L g1332 ( .A(n_589), .Y(n_1332) );
INVx2_ASAP7_75t_SL g1399 ( .A(n_589), .Y(n_1399) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OAI221xp5_ASAP7_75t_L g612 ( .A1(n_592), .A2(n_595), .B1(n_613), .B2(n_614), .C(n_615), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g1849 ( .A1(n_592), .A2(n_778), .B1(n_1831), .B2(n_1836), .Y(n_1849) );
BUFx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g867 ( .A(n_593), .Y(n_867) );
BUFx2_ASAP7_75t_L g895 ( .A(n_593), .Y(n_895) );
BUFx2_ASAP7_75t_L g995 ( .A(n_593), .Y(n_995) );
INVxp67_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
BUFx4f_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x6_ASAP7_75t_L g607 ( .A(n_596), .B(n_608), .Y(n_607) );
INVx4_ASAP7_75t_L g768 ( .A(n_596), .Y(n_768) );
BUFx4f_ASAP7_75t_L g778 ( .A(n_596), .Y(n_778) );
BUFx6f_ASAP7_75t_L g1394 ( .A(n_596), .Y(n_1394) );
BUFx4f_ASAP7_75t_L g1536 ( .A(n_596), .Y(n_1536) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx3_ASAP7_75t_L g630 ( .A(n_597), .Y(n_630) );
OAI21xp5_ASAP7_75t_L g864 ( .A1(n_598), .A2(n_607), .B(n_865), .Y(n_864) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g736 ( .A(n_601), .Y(n_736) );
INVx2_ASAP7_75t_SL g861 ( .A(n_601), .Y(n_861) );
NAND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx1_ASAP7_75t_L g608 ( .A(n_602), .Y(n_608) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_SL g859 ( .A(n_606), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_607), .Y(n_740) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_615), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_615), .B(n_856), .Y(n_855) );
INVx2_ASAP7_75t_L g1395 ( .A(n_615), .Y(n_1395) );
INVx1_ASAP7_75t_L g1848 ( .A(n_615), .Y(n_1848) );
AOI222xp33_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_621), .B1(n_622), .B2(n_627), .C1(n_628), .C2(n_631), .Y(n_617) );
AOI21xp33_ASAP7_75t_SL g738 ( .A1(n_618), .A2(n_739), .B(n_740), .Y(n_738) );
AND2x4_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
AOI222xp33_ASAP7_75t_L g734 ( .A1(n_622), .A2(n_700), .B1(n_712), .B2(n_735), .C1(n_736), .C2(n_737), .Y(n_734) );
INVx1_ASAP7_75t_L g874 ( .A(n_622), .Y(n_874) );
AND2x4_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g629 ( .A(n_624), .B(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g863 ( .A(n_624), .B(n_630), .Y(n_863) );
INVx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g1089 ( .A(n_626), .Y(n_1089) );
AOI211xp5_ASAP7_75t_L g664 ( .A1(n_627), .A2(n_665), .B(n_668), .C(n_676), .Y(n_664) );
AOI222xp33_ASAP7_75t_L g720 ( .A1(n_628), .A2(n_701), .B1(n_721), .B2(n_727), .C1(n_728), .C2(n_731), .Y(n_720) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_SL g905 ( .A(n_630), .Y(n_905) );
BUFx2_ASAP7_75t_SL g1280 ( .A(n_630), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_635), .B(n_931), .Y(n_930) );
INVx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_636), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_636), .A2(n_686), .B1(n_823), .B2(n_824), .Y(n_822) );
AND2x4_ASAP7_75t_L g686 ( .A(n_637), .B(n_687), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_664), .B(n_682), .C(n_684), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_644), .B1(n_646), .B2(n_654), .C(n_658), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x6_ASAP7_75t_SL g677 ( .A(n_642), .B(n_678), .Y(n_677) );
INVx3_ASAP7_75t_L g801 ( .A(n_642), .Y(n_801) );
BUFx2_ASAP7_75t_L g1025 ( .A(n_642), .Y(n_1025) );
BUFx2_ASAP7_75t_L g1077 ( .A(n_642), .Y(n_1077) );
INVx3_ASAP7_75t_L g710 ( .A(n_645), .Y(n_710) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g790 ( .A(n_648), .Y(n_790) );
INVx1_ASAP7_75t_L g1263 ( .A(n_648), .Y(n_1263) );
INVx1_ASAP7_75t_L g1562 ( .A(n_648), .Y(n_1562) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI221xp5_ASAP7_75t_L g703 ( .A1(n_650), .A2(n_704), .B1(n_705), .B2(n_706), .C(n_707), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g835 ( .A1(n_650), .A2(n_674), .B1(n_836), .B2(n_837), .C(n_838), .Y(n_835) );
INVx3_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_SL g840 ( .A(n_651), .Y(n_840) );
INVx5_ASAP7_75t_L g924 ( .A(n_651), .Y(n_924) );
INVx2_ASAP7_75t_SL g1164 ( .A(n_651), .Y(n_1164) );
HB1xp67_ASAP7_75t_L g1559 ( .A(n_651), .Y(n_1559) );
BUFx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
BUFx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
BUFx2_ASAP7_75t_L g959 ( .A(n_657), .Y(n_959) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_660), .A2(n_663), .B1(n_692), .B2(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx4_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_670), .A2(n_672), .B1(n_700), .B2(n_701), .Y(n_699) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g827 ( .A1(n_673), .A2(n_828), .B1(n_835), .B2(n_839), .C(n_844), .Y(n_827) );
OR2x6_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g1862 ( .A(n_674), .Y(n_1862) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_679), .Y(n_851) );
INVx3_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
HB1xp67_ASAP7_75t_L g908 ( .A(n_682), .Y(n_908) );
INVx1_ASAP7_75t_L g1242 ( .A(n_682), .Y(n_1242) );
INVx1_ASAP7_75t_L g1546 ( .A(n_682), .Y(n_1546) );
BUFx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI21x1_ASAP7_75t_L g746 ( .A1(n_683), .A2(n_747), .B(n_779), .Y(n_746) );
HB1xp67_ASAP7_75t_L g1098 ( .A(n_683), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_686), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g803 ( .A(n_686), .Y(n_803) );
AOI211x1_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .B(n_693), .C(n_719), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_711), .C(n_713), .Y(n_702) );
OAI221xp5_ASAP7_75t_L g923 ( .A1(n_705), .A2(n_903), .B1(n_924), .B2(n_925), .C(n_926), .Y(n_923) );
INVx3_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
OAI211xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B(n_717), .C(n_718), .Y(n_713) );
OAI21xp5_ASAP7_75t_SL g844 ( .A1(n_715), .A2(n_845), .B(n_846), .Y(n_844) );
INVx3_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g1210 ( .A(n_716), .Y(n_1210) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_734), .C(n_738), .Y(n_719) );
INVx2_ASAP7_75t_L g1852 ( .A(n_731), .Y(n_1852) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AO22x2_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_938), .B1(n_1009), .B2(n_1010), .Y(n_741) );
INVx1_ASAP7_75t_L g1009 ( .A(n_742), .Y(n_1009) );
XNOR2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_881), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_818), .B1(n_879), .B2(n_880), .Y(n_743) );
INVx1_ASAP7_75t_L g880 ( .A(n_744), .Y(n_880) );
NAND3xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_811), .C(n_815), .Y(n_744) );
INVx1_ASAP7_75t_L g812 ( .A(n_746), .Y(n_812) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_754), .B1(n_758), .B2(n_760), .Y(n_750) );
BUFx6f_ASAP7_75t_L g1182 ( .A(n_752), .Y(n_1182) );
INVx3_ASAP7_75t_L g1326 ( .A(n_752), .Y(n_1326) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g761 ( .A(n_756), .Y(n_761) );
INVx2_ASAP7_75t_L g1087 ( .A(n_761), .Y(n_1087) );
INVx1_ASAP7_75t_L g1148 ( .A(n_761), .Y(n_1148) );
HB1xp67_ASAP7_75t_L g1234 ( .A(n_761), .Y(n_1234) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_774), .B1(n_776), .B2(n_777), .Y(n_763) );
INVx3_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx4_ASAP7_75t_L g889 ( .A(n_766), .Y(n_889) );
BUFx6f_ASAP7_75t_L g1000 ( .A(n_766), .Y(n_1000) );
OAI211xp5_ASAP7_75t_L g1187 ( .A1(n_767), .A2(n_1188), .B(n_1189), .C(n_1192), .Y(n_1187) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g890 ( .A(n_768), .Y(n_890) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
AOI222xp33_ASAP7_75t_L g805 ( .A1(n_773), .A2(n_806), .B1(n_807), .B2(n_808), .C1(n_809), .C2(n_810), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g887 ( .A1(n_774), .A2(n_776), .B1(n_888), .B2(n_894), .Y(n_887) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NOR2x1_ASAP7_75t_L g1006 ( .A(n_775), .B(n_1007), .Y(n_1006) );
INVx1_ASAP7_75t_L g813 ( .A(n_780), .Y(n_813) );
AND2x2_ASAP7_75t_L g780 ( .A(n_781), .B(n_793), .Y(n_780) );
BUFx6f_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
BUFx6f_ASAP7_75t_L g788 ( .A(n_786), .Y(n_788) );
INVx2_ASAP7_75t_L g1119 ( .A(n_786), .Y(n_1119) );
INVx2_ASAP7_75t_L g1421 ( .A(n_786), .Y(n_1421) );
AND2x4_ASAP7_75t_L g1456 ( .A(n_786), .B(n_1434), .Y(n_1456) );
INVx1_ASAP7_75t_L g1423 ( .A(n_788), .Y(n_1423) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g1498 ( .A1(n_794), .A2(n_795), .B1(n_1499), .B2(n_1500), .Y(n_1498) );
INVx1_ASAP7_75t_L g1319 ( .A(n_795), .Y(n_1319) );
INVx1_ASAP7_75t_L g817 ( .A(n_797), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_798), .B(n_804), .Y(n_797) );
NAND2x1_ASAP7_75t_L g798 ( .A(n_799), .B(n_803), .Y(n_798) );
INVx2_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g1520 ( .A1(n_800), .A2(n_807), .B1(n_1511), .B2(n_1512), .Y(n_1520) );
AND2x2_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
INVx2_ASAP7_75t_L g1309 ( .A(n_801), .Y(n_1309) );
INVxp67_ASAP7_75t_L g934 ( .A(n_802), .Y(n_934) );
INVx1_ASAP7_75t_L g816 ( .A(n_805), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g910 ( .A1(n_806), .A2(n_809), .B1(n_893), .B2(n_911), .Y(n_910) );
OAI21xp5_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_813), .B(n_814), .Y(n_811) );
OAI21xp33_ASAP7_75t_L g815 ( .A1(n_814), .A2(n_816), .B(n_817), .Y(n_815) );
INVx1_ASAP7_75t_L g879 ( .A(n_818), .Y(n_879) );
XNOR2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
NOR2x1_ASAP7_75t_L g820 ( .A(n_821), .B(n_852), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_825), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_831), .B1(n_832), .B2(n_834), .Y(n_828) );
HB1xp67_ASAP7_75t_L g1416 ( .A(n_829), .Y(n_1416) );
INVx1_ASAP7_75t_L g1428 ( .A(n_829), .Y(n_1428) );
BUFx4f_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g933 ( .A(n_830), .Y(n_933) );
OR2x4_ASAP7_75t_L g1433 ( .A(n_830), .B(n_1434), .Y(n_1433) );
BUFx3_ASAP7_75t_L g1828 ( .A(n_830), .Y(n_1828) );
OAI22xp5_ASAP7_75t_L g1835 ( .A1(n_832), .A2(n_1836), .B1(n_1837), .B2(n_1838), .Y(n_1835) );
INVx3_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx3_ASAP7_75t_L g842 ( .A(n_833), .Y(n_842) );
INVx3_ASAP7_75t_L g918 ( .A(n_833), .Y(n_918) );
OAI211xp5_ASAP7_75t_L g865 ( .A1(n_836), .A2(n_866), .B(n_868), .C(n_869), .Y(n_865) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_840), .A2(n_841), .B1(n_842), .B2(n_843), .Y(n_839) );
OAI221xp5_ASAP7_75t_L g916 ( .A1(n_840), .A2(n_917), .B1(n_918), .B2(n_919), .C(n_920), .Y(n_916) );
OAI211xp5_ASAP7_75t_L g1304 ( .A1(n_840), .A2(n_1305), .B(n_1306), .C(n_1307), .Y(n_1304) );
OAI22xp33_ASAP7_75t_L g1208 ( .A1(n_842), .A2(n_1209), .B1(n_1210), .B2(n_1211), .Y(n_1208) );
OAI22xp5_ASAP7_75t_L g1420 ( .A1(n_842), .A2(n_1391), .B1(n_1404), .B2(n_1421), .Y(n_1420) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_849), .A2(n_859), .B1(n_860), .B2(n_861), .Y(n_858) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
NAND3xp33_ASAP7_75t_L g852 ( .A(n_853), .B(n_870), .C(n_875), .Y(n_852) );
NOR3xp33_ASAP7_75t_SL g853 ( .A(n_854), .B(n_862), .C(n_864), .Y(n_853) );
OAI21xp5_ASAP7_75t_SL g854 ( .A1(n_855), .A2(n_857), .B(n_858), .Y(n_854) );
INVx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_876), .B(n_877), .Y(n_875) );
AOI21xp5_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_908), .B(n_909), .Y(n_883) );
NAND4xp25_ASAP7_75t_L g884 ( .A(n_885), .B(n_887), .C(n_897), .D(n_902), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g1390 ( .A1(n_895), .A2(n_1391), .B1(n_1392), .B2(n_1393), .Y(n_1390) );
OAI22xp5_ASAP7_75t_L g1409 ( .A1(n_895), .A2(n_1401), .B1(n_1410), .B2(n_1411), .Y(n_1409) );
INVx2_ASAP7_75t_L g1402 ( .A(n_896), .Y(n_1402) );
OAI211xp5_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_904), .B(n_906), .C(n_907), .Y(n_902) );
OAI211xp5_ASAP7_75t_L g1594 ( .A1(n_904), .A2(n_1595), .B(n_1596), .C(n_1597), .Y(n_1594) );
OAI22xp5_ASAP7_75t_L g1850 ( .A1(n_904), .A2(n_1829), .B1(n_1843), .B2(n_1851), .Y(n_1850) );
INVx5_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
OAI22xp5_ASAP7_75t_SL g913 ( .A1(n_914), .A2(n_916), .B1(n_922), .B2(n_923), .Y(n_913) );
BUFx2_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
BUFx8_ASAP7_75t_L g1207 ( .A(n_915), .Y(n_1207) );
BUFx4f_ASAP7_75t_L g1303 ( .A(n_915), .Y(n_1303) );
BUFx4f_ASAP7_75t_L g1414 ( .A(n_915), .Y(n_1414) );
OAI22xp5_ASAP7_75t_L g1426 ( .A1(n_918), .A2(n_1400), .B1(n_1411), .B2(n_1427), .Y(n_1426) );
INVx2_ASAP7_75t_SL g955 ( .A(n_921), .Y(n_955) );
INVx1_ASAP7_75t_L g1022 ( .A(n_921), .Y(n_1022) );
BUFx3_ASAP7_75t_L g1079 ( .A(n_921), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g1302 ( .A1(n_922), .A2(n_1303), .B1(n_1304), .B2(n_1308), .Y(n_1302) );
OAI33xp33_ASAP7_75t_L g1823 ( .A1(n_922), .A2(n_1303), .A3(n_1824), .B1(n_1830), .B2(n_1835), .B3(n_1839), .Y(n_1823) );
BUFx3_ASAP7_75t_L g1216 ( .A(n_924), .Y(n_1216) );
INVx8_ASAP7_75t_L g1833 ( .A(n_924), .Y(n_1833) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_929), .B(n_930), .Y(n_928) );
OR2x6_ASAP7_75t_L g931 ( .A(n_932), .B(n_934), .Y(n_931) );
OR2x2_ASAP7_75t_L g1030 ( .A(n_932), .B(n_934), .Y(n_1030) );
INVx2_ASAP7_75t_SL g1214 ( .A(n_932), .Y(n_1214) );
INVx2_ASAP7_75t_SL g932 ( .A(n_933), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_936), .B(n_937), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_937), .B(n_950), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_937), .B(n_1159), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1257 ( .A(n_937), .B(n_1258), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1572 ( .A(n_937), .B(n_1573), .Y(n_1572) );
INVx2_ASAP7_75t_L g1010 ( .A(n_938), .Y(n_1010) );
XOR2x2_ASAP7_75t_L g938 ( .A(n_939), .B(n_1008), .Y(n_938) );
NAND2xp5_ASAP7_75t_SL g939 ( .A(n_940), .B(n_970), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_943), .B(n_952), .Y(n_942) );
NOR2xp33_ASAP7_75t_L g943 ( .A(n_944), .B(n_948), .Y(n_943) );
NAND2xp5_ASAP7_75t_SL g948 ( .A(n_949), .B(n_951), .Y(n_948) );
INVx1_ASAP7_75t_L g1126 ( .A(n_951), .Y(n_1126) );
NAND4xp25_ASAP7_75t_SL g1154 ( .A(n_951), .B(n_1155), .C(n_1158), .D(n_1160), .Y(n_1154) );
NAND4xp25_ASAP7_75t_SL g1568 ( .A(n_951), .B(n_1569), .C(n_1572), .D(n_1574), .Y(n_1568) );
INVx2_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
BUFx2_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
BUFx2_ASAP7_75t_L g1027 ( .A(n_961), .Y(n_1027) );
BUFx2_ASAP7_75t_L g1124 ( .A(n_961), .Y(n_1124) );
BUFx2_ASAP7_75t_L g1225 ( .A(n_961), .Y(n_1225) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
NAND3xp33_ASAP7_75t_SL g971 ( .A(n_972), .B(n_975), .C(n_986), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_973), .A2(n_1238), .B1(n_1239), .B2(n_1240), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g1275 ( .A1(n_973), .A2(n_1240), .B1(n_1276), .B2(n_1277), .Y(n_1275) );
INVx2_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
BUFx3_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
INVx1_ASAP7_75t_SL g984 ( .A(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx2_ASAP7_75t_L g1038 ( .A(n_989), .Y(n_1038) );
INVx2_ASAP7_75t_L g1092 ( .A(n_989), .Y(n_1092) );
INVx4_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
OAI221xp5_ASAP7_75t_L g1279 ( .A1(n_993), .A2(n_1280), .B1(n_1281), .B2(n_1282), .C(n_1283), .Y(n_1279) );
INVx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx2_ASAP7_75t_L g1851 ( .A(n_994), .Y(n_1851) );
INVx4_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g997 ( .A1(n_998), .A2(n_999), .B1(n_1001), .B2(n_1002), .Y(n_997) );
OAI221xp5_ASAP7_75t_L g1040 ( .A1(n_999), .A2(n_1002), .B1(n_1041), .B2(n_1042), .C(n_1043), .Y(n_1040) );
OAI221xp5_ASAP7_75t_L g1376 ( .A1(n_999), .A2(n_1377), .B1(n_1378), .B2(n_1379), .C(n_1380), .Y(n_1376) );
INVx2_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
INVx2_ASAP7_75t_L g1846 ( .A(n_1000), .Y(n_1846) );
OAI22xp33_ASAP7_75t_L g1853 ( .A1(n_1002), .A2(n_1834), .B1(n_1838), .B2(n_1854), .Y(n_1853) );
INVx5_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx6_ASAP7_75t_L g1847 ( .A(n_1003), .Y(n_1847) );
BUFx2_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx2_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx2_ASAP7_75t_L g1039 ( .A(n_1006), .Y(n_1039) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1011), .Y(n_1099) );
XNOR2x1_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1058), .Y(n_1011) );
NAND3xp33_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1033), .C(n_1036), .Y(n_1013) );
NOR3xp33_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1029), .C(n_1032), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1019), .Y(n_1015) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVxp67_ASAP7_75t_L g1341 ( .A(n_1031), .Y(n_1341) );
NOR4xp25_ASAP7_75t_L g1200 ( .A(n_1032), .B(n_1201), .C(n_1204), .D(n_1206), .Y(n_1200) );
NOR3xp33_ASAP7_75t_L g1348 ( .A(n_1032), .B(n_1349), .C(n_1359), .Y(n_1348) );
NOR3xp33_ASAP7_75t_L g1904 ( .A(n_1032), .B(n_1905), .C(n_1915), .Y(n_1904) );
OAI21xp5_ASAP7_75t_L g1036 ( .A1(n_1037), .A2(n_1048), .B(n_1057), .Y(n_1036) );
BUFx2_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1047), .Y(n_1283) );
OAI21xp5_ASAP7_75t_L g1130 ( .A1(n_1057), .A2(n_1131), .B(n_1140), .Y(n_1130) );
O2A1O1Ixp5_ASAP7_75t_L g1267 ( .A1(n_1057), .A2(n_1268), .B(n_1278), .C(n_1287), .Y(n_1267) );
OAI21xp5_ASAP7_75t_L g1919 ( .A1(n_1057), .A2(n_1920), .B(n_1929), .Y(n_1919) );
AND3x1_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1067), .C(n_1070), .Y(n_1063) );
INVx2_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
OAI21xp5_ASAP7_75t_L g1080 ( .A1(n_1081), .A2(n_1091), .B(n_1098), .Y(n_1080) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1085), .Y(n_1097) );
INVx2_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx2_ASAP7_75t_L g1934 ( .A(n_1087), .Y(n_1934) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
XOR2xp5_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1383), .Y(n_1102) );
OAI22xp5_ASAP7_75t_L g1103 ( .A1(n_1104), .A2(n_1248), .B1(n_1249), .B2(n_1382), .Y(n_1103) );
INVx2_ASAP7_75t_L g1382 ( .A(n_1104), .Y(n_1382) );
AO22x2_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1106), .B1(n_1197), .B2(n_1247), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
OAI22xp5_ASAP7_75t_L g1106 ( .A1(n_1107), .A2(n_1108), .B1(n_1150), .B2(n_1196), .Y(n_1106) );
INVx2_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
NAND3xp33_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1127), .C(n_1130), .Y(n_1109) );
NOR3xp33_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1125), .C(n_1126), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1115), .Y(n_1111) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
NOR3xp33_ASAP7_75t_L g1550 ( .A(n_1126), .B(n_1551), .C(n_1563), .Y(n_1550) );
HB1xp67_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1150), .Y(n_1196) );
NAND2x1p5_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1169), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1167), .Y(n_1152) );
INVxp67_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
NOR2xp33_ASAP7_75t_SL g1193 ( .A(n_1154), .B(n_1194), .Y(n_1193) );
INVx2_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1167), .B(n_1195), .Y(n_1194) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1172), .B(n_1176), .Y(n_1171) );
AOI21xp5_ASAP7_75t_L g1172 ( .A1(n_1173), .A2(n_1174), .B(n_1175), .Y(n_1172) );
AOI21xp5_ASAP7_75t_L g1582 ( .A1(n_1173), .A2(n_1583), .B(n_1584), .Y(n_1582) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1180), .Y(n_1368) );
BUFx2_ASAP7_75t_L g1923 ( .A(n_1180), .Y(n_1923) );
HB1xp67_ASAP7_75t_L g1272 ( .A(n_1182), .Y(n_1272) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1197), .Y(n_1247) );
XNOR2xp5_ASAP7_75t_SL g1197 ( .A(n_1198), .B(n_1199), .Y(n_1197) );
AND3x2_ASAP7_75t_L g1199 ( .A(n_1200), .B(n_1226), .C(n_1243), .Y(n_1199) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
OAI33xp33_ASAP7_75t_L g1206 ( .A1(n_1207), .A2(n_1208), .A3(n_1212), .B1(n_1218), .B2(n_1221), .B3(n_1224), .Y(n_1206) );
OAI22xp33_ASAP7_75t_L g1221 ( .A1(n_1210), .A2(n_1213), .B1(n_1222), .B2(n_1223), .Y(n_1221) );
OAI22xp5_ASAP7_75t_L g1212 ( .A1(n_1213), .A2(n_1215), .B1(n_1216), .B2(n_1217), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1216), .Y(n_1262) );
OAI33xp33_ASAP7_75t_L g1412 ( .A1(n_1224), .A2(n_1413), .A3(n_1415), .B1(n_1420), .B2(n_1422), .B3(n_1426), .Y(n_1412) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
OAI21xp5_ASAP7_75t_L g1226 ( .A1(n_1227), .A2(n_1231), .B(n_1241), .Y(n_1226) );
OAI21xp5_ASAP7_75t_L g1363 ( .A1(n_1241), .A2(n_1364), .B(n_1375), .Y(n_1363) );
INVx2_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
AOI22xp5_ASAP7_75t_L g1249 ( .A1(n_1250), .A2(n_1344), .B1(n_1345), .B2(n_1381), .Y(n_1249) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1250), .Y(n_1381) );
OAI22xp5_ASAP7_75t_L g1250 ( .A1(n_1251), .A2(n_1292), .B1(n_1342), .B2(n_1343), .Y(n_1250) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1251), .Y(n_1342) );
XOR2x2_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1291), .Y(n_1251) );
NAND3x1_ASAP7_75t_SL g1252 ( .A(n_1253), .B(n_1267), .C(n_1289), .Y(n_1252) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1292), .Y(n_1343) );
HB1xp67_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
NAND4xp75_ASAP7_75t_L g1294 ( .A(n_1295), .B(n_1301), .C(n_1320), .D(n_1340), .Y(n_1294) );
INVx1_ASAP7_75t_SL g1298 ( .A(n_1299), .Y(n_1298) );
OAI221xp5_ASAP7_75t_L g1308 ( .A1(n_1309), .A2(n_1310), .B1(n_1311), .B2(n_1313), .C(n_1314), .Y(n_1308) );
OAI22xp5_ASAP7_75t_L g1830 ( .A1(n_1311), .A2(n_1831), .B1(n_1832), .B2(n_1834), .Y(n_1830) );
BUFx3_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
OAI21xp5_ASAP7_75t_L g1320 ( .A1(n_1321), .A2(n_1330), .B(n_1339), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1327), .Y(n_1321) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
INVx2_ASAP7_75t_SL g1538 ( .A(n_1326), .Y(n_1538) );
OAI221xp5_ASAP7_75t_L g1331 ( .A1(n_1332), .A2(n_1333), .B1(n_1334), .B2(n_1336), .C(n_1337), .Y(n_1331) );
BUFx3_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
OAI21xp33_ASAP7_75t_L g1585 ( .A1(n_1339), .A2(n_1586), .B(n_1593), .Y(n_1585) );
INVx2_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
INVx2_ASAP7_75t_SL g1345 ( .A(n_1346), .Y(n_1345) );
NAND3xp33_ASAP7_75t_L g1347 ( .A(n_1348), .B(n_1360), .C(n_1363), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1353), .Y(n_1349) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1368), .Y(n_1367) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
OAI22xp5_ASAP7_75t_L g1384 ( .A1(n_1385), .A2(n_1522), .B1(n_1523), .B2(n_1598), .Y(n_1384) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1385), .Y(n_1598) );
AO22x1_ASAP7_75t_L g1385 ( .A1(n_1386), .A2(n_1491), .B1(n_1492), .B2(n_1521), .Y(n_1385) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1386), .Y(n_1521) );
NAND3xp33_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1429), .C(n_1462), .Y(n_1387) );
NOR2xp33_ASAP7_75t_L g1388 ( .A(n_1389), .B(n_1412), .Y(n_1388) );
OAI33xp33_ASAP7_75t_L g1389 ( .A1(n_1390), .A2(n_1395), .A3(n_1396), .B1(n_1403), .B2(n_1406), .B3(n_1409), .Y(n_1389) );
OAI22xp5_ASAP7_75t_L g1422 ( .A1(n_1392), .A2(n_1405), .B1(n_1423), .B2(n_1424), .Y(n_1422) );
HB1xp67_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
OAI22xp33_ASAP7_75t_L g1403 ( .A1(n_1394), .A2(n_1398), .B1(n_1404), .B2(n_1405), .Y(n_1403) );
OAI22xp5_ASAP7_75t_L g1396 ( .A1(n_1397), .A2(n_1398), .B1(n_1400), .B2(n_1401), .Y(n_1396) );
OAI22xp33_ASAP7_75t_L g1415 ( .A1(n_1397), .A2(n_1410), .B1(n_1416), .B2(n_1417), .Y(n_1415) );
INVx2_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
INVx2_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVx2_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
BUFx3_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
INVx2_ASAP7_75t_SL g1417 ( .A(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
OAI22xp33_ASAP7_75t_L g1824 ( .A1(n_1424), .A2(n_1825), .B1(n_1826), .B2(n_1829), .Y(n_1824) );
BUFx6f_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
INVx2_ASAP7_75t_L g1842 ( .A(n_1425), .Y(n_1842) );
INVx2_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
OAI31xp33_ASAP7_75t_L g1429 ( .A1(n_1430), .A2(n_1438), .A3(n_1451), .B(n_1457), .Y(n_1429) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
INVx2_ASAP7_75t_L g1868 ( .A(n_1432), .Y(n_1868) );
INVx2_ASAP7_75t_SL g1432 ( .A(n_1433), .Y(n_1432) );
INVx2_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
INVx2_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
BUFx3_ASAP7_75t_L g1869 ( .A(n_1437), .Y(n_1869) );
CKINVDCx8_ASAP7_75t_R g1439 ( .A(n_1440), .Y(n_1439) );
AOI22xp33_ASAP7_75t_L g1441 ( .A1(n_1442), .A2(n_1443), .B1(n_1447), .B2(n_1448), .Y(n_1441) );
AOI22xp33_ASAP7_75t_L g1481 ( .A1(n_1442), .A2(n_1482), .B1(n_1484), .B2(n_1485), .Y(n_1481) );
BUFx3_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
BUFx3_ASAP7_75t_L g1864 ( .A(n_1444), .Y(n_1864) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1446), .Y(n_1444) );
AND2x4_ASAP7_75t_L g1449 ( .A(n_1445), .B(n_1450), .Y(n_1449) );
AOI22xp33_ASAP7_75t_L g1863 ( .A1(n_1448), .A2(n_1864), .B1(n_1865), .B2(n_1866), .Y(n_1863) );
BUFx6f_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
HB1xp67_ASAP7_75t_L g1871 ( .A(n_1454), .Y(n_1871) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
INVx1_ASAP7_75t_L g1872 ( .A(n_1456), .Y(n_1872) );
AND2x2_ASAP7_75t_SL g1457 ( .A(n_1458), .B(n_1460), .Y(n_1457) );
AND2x4_ASAP7_75t_L g1873 ( .A(n_1458), .B(n_1460), .Y(n_1873) );
INVx1_ASAP7_75t_SL g1458 ( .A(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
OAI31xp33_ASAP7_75t_SL g1462 ( .A1(n_1463), .A2(n_1468), .A3(n_1477), .B(n_1488), .Y(n_1462) );
INVx3_ASAP7_75t_SL g1465 ( .A(n_1466), .Y(n_1465) );
CKINVDCx16_ASAP7_75t_R g1876 ( .A(n_1466), .Y(n_1876) );
HB1xp67_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
INVx1_ASAP7_75t_L g1879 ( .A(n_1470), .Y(n_1879) );
INVx2_ASAP7_75t_L g1471 ( .A(n_1472), .Y(n_1471) );
INVx2_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
INVx2_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
BUFx2_ASAP7_75t_L g1882 ( .A(n_1475), .Y(n_1882) );
INVx3_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1886 ( .A(n_1479), .Y(n_1886) );
AOI22xp33_ASAP7_75t_L g1887 ( .A1(n_1482), .A2(n_1865), .B1(n_1888), .B2(n_1890), .Y(n_1887) );
BUFx3_ASAP7_75t_L g1482 ( .A(n_1483), .Y(n_1482) );
INVx2_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
INVx2_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
INVx2_ASAP7_75t_L g1889 ( .A(n_1487), .Y(n_1889) );
BUFx3_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
BUFx2_ASAP7_75t_SL g1891 ( .A(n_1489), .Y(n_1891) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1494), .B(n_1508), .Y(n_1493) );
AOI22xp5_ASAP7_75t_L g1501 ( .A1(n_1502), .A2(n_1504), .B1(n_1505), .B2(n_1507), .Y(n_1501) );
NAND3xp33_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1513), .C(n_1516), .Y(n_1509) );
INVx2_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
XNOR2x2_ASAP7_75t_L g1523 ( .A(n_1524), .B(n_1564), .Y(n_1523) );
NAND3xp33_ASAP7_75t_L g1525 ( .A(n_1526), .B(n_1547), .C(n_1550), .Y(n_1525) );
OAI31xp33_ASAP7_75t_L g1526 ( .A1(n_1527), .A2(n_1533), .A3(n_1544), .B(n_1545), .Y(n_1526) );
NAND2xp5_ASAP7_75t_L g1527 ( .A(n_1528), .B(n_1530), .Y(n_1527) );
OAI211xp5_ASAP7_75t_L g1534 ( .A1(n_1535), .A2(n_1536), .B(n_1537), .C(n_1539), .Y(n_1534) );
INVx1_ASAP7_75t_L g1885 ( .A(n_1536), .Y(n_1885) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
NAND2xp5_ASAP7_75t_L g1551 ( .A(n_1552), .B(n_1555), .Y(n_1551) );
XNOR2x2_ASAP7_75t_L g1564 ( .A(n_1565), .B(n_1566), .Y(n_1564) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
NAND2xp5_ASAP7_75t_L g1581 ( .A(n_1582), .B(n_1585), .Y(n_1581) );
OAI221xp5_ASAP7_75t_L g1599 ( .A1(n_1600), .A2(n_1814), .B1(n_1818), .B2(n_1892), .C(n_1895), .Y(n_1599) );
AOI21xp5_ASAP7_75t_L g1600 ( .A1(n_1601), .A2(n_1740), .B(n_1788), .Y(n_1600) );
NAND5xp2_ASAP7_75t_L g1601 ( .A(n_1602), .B(n_1690), .C(n_1706), .D(n_1719), .E(n_1732), .Y(n_1601) );
AOI211xp5_ASAP7_75t_L g1602 ( .A1(n_1603), .A2(n_1634), .B(n_1649), .C(n_1674), .Y(n_1602) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1604), .B(n_1620), .Y(n_1603) );
AND2x2_ASAP7_75t_L g1766 ( .A(n_1604), .B(n_1701), .Y(n_1766) );
CKINVDCx5p33_ASAP7_75t_R g1604 ( .A(n_1605), .Y(n_1604) );
OR2x2_ASAP7_75t_L g1692 ( .A(n_1605), .B(n_1658), .Y(n_1692) );
AND2x2_ASAP7_75t_L g1700 ( .A(n_1605), .B(n_1701), .Y(n_1700) );
AOI322xp5_ASAP7_75t_L g1719 ( .A1(n_1605), .A2(n_1676), .A3(n_1720), .B1(n_1724), .B2(n_1725), .C1(n_1729), .C2(n_1730), .Y(n_1719) );
NAND2xp5_ASAP7_75t_L g1758 ( .A(n_1605), .B(n_1759), .Y(n_1758) );
NAND2xp5_ASAP7_75t_L g1775 ( .A(n_1605), .B(n_1776), .Y(n_1775) );
NAND2xp5_ASAP7_75t_L g1804 ( .A(n_1605), .B(n_1666), .Y(n_1804) );
O2A1O1Ixp33_ASAP7_75t_SL g1810 ( .A1(n_1605), .A2(n_1660), .B(n_1675), .C(n_1760), .Y(n_1810) );
INVx4_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
INVx4_ASAP7_75t_L g1656 ( .A(n_1606), .Y(n_1656) );
NAND2xp5_ASAP7_75t_SL g1665 ( .A(n_1606), .B(n_1622), .Y(n_1665) );
AND2x2_ASAP7_75t_L g1693 ( .A(n_1606), .B(n_1694), .Y(n_1693) );
NOR2xp33_ASAP7_75t_L g1709 ( .A(n_1606), .B(n_1641), .Y(n_1709) );
OR2x2_ASAP7_75t_L g1728 ( .A(n_1606), .B(n_1622), .Y(n_1728) );
NOR2xp33_ASAP7_75t_L g1729 ( .A(n_1606), .B(n_1627), .Y(n_1729) );
NAND2xp5_ASAP7_75t_L g1755 ( .A(n_1606), .B(n_1735), .Y(n_1755) );
AND2x2_ASAP7_75t_L g1787 ( .A(n_1606), .B(n_1695), .Y(n_1787) );
AOI321xp33_ASAP7_75t_R g1799 ( .A1(n_1606), .A2(n_1634), .A3(n_1693), .B1(n_1705), .B2(n_1724), .C(n_1800), .Y(n_1799) );
AND2x4_ASAP7_75t_SL g1606 ( .A(n_1607), .B(n_1615), .Y(n_1606) );
AND2x4_ASAP7_75t_L g1608 ( .A(n_1609), .B(n_1610), .Y(n_1608) );
AND2x6_ASAP7_75t_L g1613 ( .A(n_1609), .B(n_1614), .Y(n_1613) );
AND2x6_ASAP7_75t_L g1616 ( .A(n_1609), .B(n_1617), .Y(n_1616) );
AND2x2_ASAP7_75t_L g1618 ( .A(n_1609), .B(n_1619), .Y(n_1618) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_1609), .B(n_1619), .Y(n_1625) );
AND2x2_ASAP7_75t_L g1640 ( .A(n_1609), .B(n_1619), .Y(n_1640) );
NAND2xp5_ASAP7_75t_L g1685 ( .A(n_1609), .B(n_1610), .Y(n_1685) );
AND2x2_ASAP7_75t_L g1610 ( .A(n_1611), .B(n_1612), .Y(n_1610) );
INVx2_ASAP7_75t_L g1687 ( .A(n_1613), .Y(n_1687) );
OAI21xp5_ASAP7_75t_L g1935 ( .A1(n_1619), .A2(n_1936), .B(n_1937), .Y(n_1935) );
AOI221xp5_ASAP7_75t_L g1808 ( .A1(n_1620), .A2(n_1750), .B1(n_1773), .B2(n_1809), .C(n_1810), .Y(n_1808) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_1621), .B(n_1626), .Y(n_1620) );
OR2x2_ASAP7_75t_L g1670 ( .A(n_1621), .B(n_1627), .Y(n_1670) );
AND2x2_ASAP7_75t_L g1694 ( .A(n_1621), .B(n_1695), .Y(n_1694) );
OR2x2_ASAP7_75t_L g1760 ( .A(n_1621), .B(n_1660), .Y(n_1760) );
AND2x2_ASAP7_75t_L g1790 ( .A(n_1621), .B(n_1739), .Y(n_1790) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
NAND2xp5_ASAP7_75t_L g1708 ( .A(n_1622), .B(n_1631), .Y(n_1708) );
OR2x2_ASAP7_75t_L g1712 ( .A(n_1622), .B(n_1628), .Y(n_1712) );
AND2x2_ASAP7_75t_L g1714 ( .A(n_1622), .B(n_1666), .Y(n_1714) );
AND2x2_ASAP7_75t_L g1717 ( .A(n_1622), .B(n_1718), .Y(n_1717) );
AND2x2_ASAP7_75t_L g1771 ( .A(n_1622), .B(n_1696), .Y(n_1771) );
OR2x2_ASAP7_75t_L g1807 ( .A(n_1622), .B(n_1696), .Y(n_1807) );
AND2x2_ASAP7_75t_L g1622 ( .A(n_1623), .B(n_1624), .Y(n_1622) );
AND2x2_ASAP7_75t_L g1659 ( .A(n_1623), .B(n_1624), .Y(n_1659) );
NAND2xp5_ASAP7_75t_L g1699 ( .A(n_1626), .B(n_1700), .Y(n_1699) );
NAND3xp33_ASAP7_75t_L g1753 ( .A(n_1626), .B(n_1745), .C(n_1754), .Y(n_1753) );
NAND2xp5_ASAP7_75t_L g1767 ( .A(n_1626), .B(n_1752), .Y(n_1767) );
AND2x2_ASAP7_75t_L g1798 ( .A(n_1626), .B(n_1664), .Y(n_1798) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1627), .Y(n_1626) );
OR2x2_ASAP7_75t_L g1748 ( .A(n_1627), .B(n_1728), .Y(n_1748) );
OR2x2_ASAP7_75t_L g1627 ( .A(n_1628), .B(n_1631), .Y(n_1627) );
NAND2xp5_ASAP7_75t_L g1660 ( .A(n_1628), .B(n_1661), .Y(n_1660) );
AND2x2_ASAP7_75t_L g1666 ( .A(n_1628), .B(n_1631), .Y(n_1666) );
INVx2_ASAP7_75t_L g1696 ( .A(n_1628), .Y(n_1696) );
NAND2x1p5_ASAP7_75t_L g1628 ( .A(n_1629), .B(n_1630), .Y(n_1628) );
INVx1_ASAP7_75t_L g1661 ( .A(n_1631), .Y(n_1661) );
AND2x2_ASAP7_75t_L g1695 ( .A(n_1631), .B(n_1696), .Y(n_1695) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1631), .Y(n_1718) );
OR2x2_ASAP7_75t_L g1777 ( .A(n_1631), .B(n_1659), .Y(n_1777) );
AND2x2_ASAP7_75t_L g1631 ( .A(n_1632), .B(n_1633), .Y(n_1631) );
AOI221xp5_ASAP7_75t_L g1789 ( .A1(n_1634), .A2(n_1679), .B1(n_1790), .B2(n_1791), .C(n_1792), .Y(n_1789) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1635), .Y(n_1634) );
OR2x2_ASAP7_75t_L g1635 ( .A(n_1636), .B(n_1641), .Y(n_1635) );
AOI221xp5_ASAP7_75t_L g1690 ( .A1(n_1636), .A2(n_1676), .B1(n_1691), .B2(n_1693), .C(n_1697), .Y(n_1690) );
AOI221xp5_ASAP7_75t_L g1706 ( .A1(n_1636), .A2(n_1707), .B1(n_1709), .B2(n_1710), .C(n_1715), .Y(n_1706) );
OAI322xp33_ASAP7_75t_L g1764 ( .A1(n_1636), .A2(n_1659), .A3(n_1765), .B1(n_1767), .B2(n_1768), .C1(n_1769), .C2(n_1770), .Y(n_1764) );
AND2x2_ASAP7_75t_L g1786 ( .A(n_1636), .B(n_1752), .Y(n_1786) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
INVx3_ASAP7_75t_L g1652 ( .A(n_1637), .Y(n_1652) );
AND2x2_ASAP7_75t_L g1668 ( .A(n_1637), .B(n_1669), .Y(n_1668) );
AND2x2_ASAP7_75t_L g1704 ( .A(n_1637), .B(n_1645), .Y(n_1704) );
OR2x2_ASAP7_75t_L g1736 ( .A(n_1637), .B(n_1645), .Y(n_1736) );
AND2x2_ASAP7_75t_L g1637 ( .A(n_1638), .B(n_1639), .Y(n_1637) );
HB1xp67_ASAP7_75t_L g1817 ( .A(n_1640), .Y(n_1817) );
AOI21xp33_ASAP7_75t_L g1813 ( .A1(n_1641), .A2(n_1692), .B(n_1713), .Y(n_1813) );
OR2x2_ASAP7_75t_L g1641 ( .A(n_1642), .B(n_1645), .Y(n_1641) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1642), .Y(n_1657) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1642), .Y(n_1673) );
NAND2xp5_ASAP7_75t_L g1642 ( .A(n_1643), .B(n_1644), .Y(n_1642) );
A2O1A1Ixp33_ASAP7_75t_L g1662 ( .A1(n_1645), .A2(n_1663), .B(n_1667), .C(n_1671), .Y(n_1662) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1645), .Y(n_1669) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1645), .B(n_1652), .Y(n_1676) );
OR2x2_ASAP7_75t_L g1702 ( .A(n_1645), .B(n_1673), .Y(n_1702) );
OAI22xp5_ASAP7_75t_L g1710 ( .A1(n_1645), .A2(n_1711), .B1(n_1712), .B2(n_1713), .Y(n_1710) );
AND2x2_ASAP7_75t_L g1724 ( .A(n_1645), .B(n_1657), .Y(n_1724) );
INVx2_ASAP7_75t_L g1745 ( .A(n_1645), .Y(n_1745) );
INVx2_ASAP7_75t_L g1645 ( .A(n_1646), .Y(n_1645) );
OR2x2_ASAP7_75t_L g1738 ( .A(n_1646), .B(n_1673), .Y(n_1738) );
NAND2xp5_ASAP7_75t_L g1646 ( .A(n_1647), .B(n_1648), .Y(n_1646) );
NAND2xp5_ASAP7_75t_L g1649 ( .A(n_1650), .B(n_1662), .Y(n_1649) );
NAND2xp5_ASAP7_75t_L g1650 ( .A(n_1651), .B(n_1653), .Y(n_1650) );
CKINVDCx14_ASAP7_75t_R g1651 ( .A(n_1652), .Y(n_1651) );
NAND2xp5_ASAP7_75t_L g1731 ( .A(n_1652), .B(n_1657), .Y(n_1731) );
OR2x2_ASAP7_75t_L g1763 ( .A(n_1652), .B(n_1672), .Y(n_1763) );
OR2x2_ASAP7_75t_L g1768 ( .A(n_1652), .B(n_1657), .Y(n_1768) );
OR2x2_ASAP7_75t_L g1769 ( .A(n_1652), .B(n_1702), .Y(n_1769) );
AND2x2_ASAP7_75t_L g1773 ( .A(n_1652), .B(n_1701), .Y(n_1773) );
O2A1O1Ixp33_ASAP7_75t_SL g1792 ( .A1(n_1652), .A2(n_1723), .B(n_1793), .C(n_1795), .Y(n_1792) );
OR2x2_ASAP7_75t_L g1806 ( .A(n_1652), .B(n_1738), .Y(n_1806) );
A2O1A1Ixp33_ASAP7_75t_R g1811 ( .A1(n_1652), .A2(n_1766), .B(n_1812), .C(n_1813), .Y(n_1811) );
AOI221xp5_ASAP7_75t_L g1741 ( .A1(n_1653), .A2(n_1676), .B1(n_1702), .B2(n_1742), .C(n_1747), .Y(n_1741) );
NOR2xp33_ASAP7_75t_L g1653 ( .A(n_1654), .B(n_1658), .Y(n_1653) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1655), .Y(n_1654) );
OAI21xp33_ASAP7_75t_L g1703 ( .A1(n_1655), .A2(n_1704), .B(n_1705), .Y(n_1703) );
AND2x2_ASAP7_75t_L g1655 ( .A(n_1656), .B(n_1657), .Y(n_1655) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1656), .B(n_1680), .Y(n_1679) );
NOR2x1_ASAP7_75t_L g1739 ( .A(n_1656), .B(n_1722), .Y(n_1739) );
NAND2x1_ASAP7_75t_L g1743 ( .A(n_1656), .B(n_1714), .Y(n_1743) );
CKINVDCx5p33_ASAP7_75t_R g1752 ( .A(n_1656), .Y(n_1752) );
NOR2xp33_ASAP7_75t_L g1794 ( .A(n_1656), .B(n_1669), .Y(n_1794) );
INVx2_ASAP7_75t_L g1735 ( .A(n_1657), .Y(n_1735) );
AND2x2_ASAP7_75t_L g1751 ( .A(n_1657), .B(n_1752), .Y(n_1751) );
NAND2xp5_ASAP7_75t_L g1707 ( .A(n_1658), .B(n_1708), .Y(n_1707) );
OR2x2_ASAP7_75t_L g1658 ( .A(n_1659), .B(n_1660), .Y(n_1658) );
AND2x2_ASAP7_75t_L g1705 ( .A(n_1659), .B(n_1695), .Y(n_1705) );
OR2x2_ASAP7_75t_L g1721 ( .A(n_1659), .B(n_1722), .Y(n_1721) );
AOI321xp33_ASAP7_75t_L g1783 ( .A1(n_1659), .A2(n_1681), .A3(n_1730), .B1(n_1784), .B2(n_1786), .C(n_1787), .Y(n_1783) );
OAI221xp5_ASAP7_75t_L g1674 ( .A1(n_1660), .A2(n_1675), .B1(n_1677), .B2(n_1678), .C(n_1681), .Y(n_1674) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1660), .Y(n_1680) );
NAND2xp5_ASAP7_75t_L g1784 ( .A(n_1660), .B(n_1785), .Y(n_1784) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1663), .Y(n_1698) );
AND2x2_ASAP7_75t_L g1663 ( .A(n_1664), .B(n_1666), .Y(n_1663) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1665), .Y(n_1664) );
INVx1_ASAP7_75t_L g1722 ( .A(n_1666), .Y(n_1722) );
NAND2xp5_ASAP7_75t_L g1726 ( .A(n_1666), .B(n_1727), .Y(n_1726) );
OAI31xp33_ASAP7_75t_L g1732 ( .A1(n_1667), .A2(n_1733), .A3(n_1737), .B(n_1739), .Y(n_1732) );
NOR2xp33_ASAP7_75t_L g1667 ( .A(n_1668), .B(n_1670), .Y(n_1667) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1668), .Y(n_1677) );
AOI221xp5_ASAP7_75t_L g1772 ( .A1(n_1668), .A2(n_1773), .B1(n_1774), .B2(n_1778), .C(n_1779), .Y(n_1772) );
OAI22xp5_ASAP7_75t_L g1742 ( .A1(n_1669), .A2(n_1743), .B1(n_1744), .B2(n_1746), .Y(n_1742) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1670), .Y(n_1782) );
OAI211xp5_ASAP7_75t_L g1697 ( .A1(n_1671), .A2(n_1698), .B(n_1699), .C(n_1703), .Y(n_1697) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
NAND2xp5_ASAP7_75t_L g1675 ( .A(n_1672), .B(n_1676), .Y(n_1675) );
INVx1_ASAP7_75t_L g1672 ( .A(n_1673), .Y(n_1672) );
NOR2xp33_ASAP7_75t_L g1796 ( .A(n_1673), .B(n_1797), .Y(n_1796) );
A2O1A1Ixp33_ASAP7_75t_L g1801 ( .A1(n_1673), .A2(n_1704), .B(n_1739), .C(n_1761), .Y(n_1801) );
AND2x2_ASAP7_75t_L g1809 ( .A(n_1676), .B(n_1751), .Y(n_1809) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
INVx2_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1683), .Y(n_1682) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
OAI221xp5_ASAP7_75t_L g1684 ( .A1(n_1685), .A2(n_1686), .B1(n_1687), .B2(n_1688), .C(n_1689), .Y(n_1684) );
INVx1_ASAP7_75t_L g1691 ( .A(n_1692), .Y(n_1691) );
NAND2xp5_ASAP7_75t_L g1746 ( .A(n_1695), .B(n_1727), .Y(n_1746) );
INVx1_ASAP7_75t_L g1785 ( .A(n_1695), .Y(n_1785) );
INVx1_ASAP7_75t_L g1711 ( .A(n_1700), .Y(n_1711) );
NAND2xp5_ASAP7_75t_L g1716 ( .A(n_1700), .B(n_1717), .Y(n_1716) );
CKINVDCx5p33_ASAP7_75t_R g1701 ( .A(n_1702), .Y(n_1701) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1708), .Y(n_1812) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1712), .Y(n_1750) );
INVx1_ASAP7_75t_L g1713 ( .A(n_1714), .Y(n_1713) );
INVxp67_ASAP7_75t_L g1715 ( .A(n_1716), .Y(n_1715) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1717), .Y(n_1723) );
NAND2xp5_ASAP7_75t_SL g1720 ( .A(n_1721), .B(n_1723), .Y(n_1720) );
INVx1_ASAP7_75t_L g1778 ( .A(n_1721), .Y(n_1778) );
INVx1_ASAP7_75t_L g1725 ( .A(n_1726), .Y(n_1725) );
OAI211xp5_ASAP7_75t_L g1802 ( .A1(n_1727), .A2(n_1803), .B(n_1805), .C(n_1807), .Y(n_1802) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1731), .Y(n_1730) );
INVx1_ASAP7_75t_L g1733 ( .A(n_1734), .Y(n_1733) );
OR2x2_ASAP7_75t_L g1734 ( .A(n_1735), .B(n_1736), .Y(n_1734) );
CKINVDCx5p33_ASAP7_75t_R g1737 ( .A(n_1738), .Y(n_1737) );
OAI211xp5_ASAP7_75t_L g1747 ( .A1(n_1738), .A2(n_1748), .B(n_1749), .C(n_1753), .Y(n_1747) );
NAND4xp25_ASAP7_75t_L g1740 ( .A(n_1741), .B(n_1756), .C(n_1772), .D(n_1783), .Y(n_1740) );
NAND3xp33_ASAP7_75t_L g1749 ( .A(n_1744), .B(n_1750), .C(n_1751), .Y(n_1749) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
INVx1_ASAP7_75t_L g1761 ( .A(n_1748), .Y(n_1761) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1755), .Y(n_1754) );
O2A1O1Ixp33_ASAP7_75t_L g1756 ( .A1(n_1757), .A2(n_1761), .B(n_1762), .C(n_1764), .Y(n_1756) );
INVxp67_ASAP7_75t_L g1757 ( .A(n_1758), .Y(n_1757) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1763), .Y(n_1762) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1766), .Y(n_1765) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1768), .Y(n_1781) );
INVx1_ASAP7_75t_L g1791 ( .A(n_1769), .Y(n_1791) );
CKINVDCx14_ASAP7_75t_R g1770 ( .A(n_1771), .Y(n_1770) );
INVx1_ASAP7_75t_L g1774 ( .A(n_1775), .Y(n_1774) );
INVxp67_ASAP7_75t_L g1776 ( .A(n_1777), .Y(n_1776) );
INVx1_ASAP7_75t_L g1779 ( .A(n_1780), .Y(n_1779) );
NAND2xp5_ASAP7_75t_L g1780 ( .A(n_1781), .B(n_1782), .Y(n_1780) );
NAND4xp25_ASAP7_75t_L g1788 ( .A(n_1789), .B(n_1799), .C(n_1808), .D(n_1811), .Y(n_1788) );
INVx1_ASAP7_75t_L g1793 ( .A(n_1794), .Y(n_1793) );
INVx1_ASAP7_75t_L g1795 ( .A(n_1796), .Y(n_1795) );
INVx1_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
NAND2xp5_ASAP7_75t_SL g1800 ( .A(n_1801), .B(n_1802), .Y(n_1800) );
INVxp67_ASAP7_75t_SL g1803 ( .A(n_1804), .Y(n_1803) );
INVx1_ASAP7_75t_L g1805 ( .A(n_1806), .Y(n_1805) );
CKINVDCx20_ASAP7_75t_R g1814 ( .A(n_1815), .Y(n_1814) );
CKINVDCx20_ASAP7_75t_R g1815 ( .A(n_1816), .Y(n_1815) );
INVx4_ASAP7_75t_L g1816 ( .A(n_1817), .Y(n_1816) );
INVx1_ASAP7_75t_L g1818 ( .A(n_1819), .Y(n_1818) );
INVx1_ASAP7_75t_L g1819 ( .A(n_1820), .Y(n_1819) );
AND3x1_ASAP7_75t_L g1821 ( .A(n_1822), .B(n_1858), .C(n_1874), .Y(n_1821) );
NOR2xp33_ASAP7_75t_L g1822 ( .A(n_1823), .B(n_1844), .Y(n_1822) );
OAI22xp33_ASAP7_75t_L g1845 ( .A1(n_1825), .A2(n_1840), .B1(n_1846), .B2(n_1847), .Y(n_1845) );
OAI22xp33_ASAP7_75t_L g1839 ( .A1(n_1826), .A2(n_1840), .B1(n_1841), .B2(n_1843), .Y(n_1839) );
INVx2_ASAP7_75t_L g1826 ( .A(n_1827), .Y(n_1826) );
INVx1_ASAP7_75t_L g1827 ( .A(n_1828), .Y(n_1827) );
INVx2_ASAP7_75t_L g1832 ( .A(n_1833), .Y(n_1832) );
INVx1_ASAP7_75t_L g1912 ( .A(n_1837), .Y(n_1912) );
INVx2_ASAP7_75t_L g1841 ( .A(n_1842), .Y(n_1841) );
OAI33xp33_ASAP7_75t_L g1844 ( .A1(n_1845), .A2(n_1848), .A3(n_1849), .B1(n_1850), .B2(n_1852), .B3(n_1853), .Y(n_1844) );
INVx1_ASAP7_75t_L g1854 ( .A(n_1855), .Y(n_1854) );
INVx1_ASAP7_75t_L g1855 ( .A(n_1856), .Y(n_1855) );
INVx1_ASAP7_75t_L g1856 ( .A(n_1857), .Y(n_1856) );
OAI31xp33_ASAP7_75t_L g1858 ( .A1(n_1859), .A2(n_1867), .A3(n_1870), .B(n_1873), .Y(n_1858) );
HB1xp67_ASAP7_75t_L g1860 ( .A(n_1861), .Y(n_1860) );
INVxp67_ASAP7_75t_SL g1861 ( .A(n_1862), .Y(n_1861) );
OAI31xp33_ASAP7_75t_L g1874 ( .A1(n_1875), .A2(n_1877), .A3(n_1883), .B(n_1891), .Y(n_1874) );
INVx1_ASAP7_75t_L g1878 ( .A(n_1879), .Y(n_1878) );
INVx1_ASAP7_75t_L g1880 ( .A(n_1881), .Y(n_1880) );
INVx2_ASAP7_75t_SL g1881 ( .A(n_1882), .Y(n_1881) );
INVx1_ASAP7_75t_L g1884 ( .A(n_1885), .Y(n_1884) );
INVx2_ASAP7_75t_L g1888 ( .A(n_1889), .Y(n_1888) );
INVx3_ASAP7_75t_L g1892 ( .A(n_1893), .Y(n_1892) );
HB1xp67_ASAP7_75t_L g1896 ( .A(n_1897), .Y(n_1896) );
BUFx3_ASAP7_75t_L g1897 ( .A(n_1898), .Y(n_1897) );
INVxp33_ASAP7_75t_SL g1899 ( .A(n_1900), .Y(n_1899) );
INVx1_ASAP7_75t_L g1901 ( .A(n_1902), .Y(n_1901) );
HB1xp67_ASAP7_75t_L g1902 ( .A(n_1903), .Y(n_1902) );
NAND3xp33_ASAP7_75t_L g1903 ( .A(n_1904), .B(n_1916), .C(n_1919), .Y(n_1903) );
NAND2xp5_ASAP7_75t_L g1905 ( .A(n_1906), .B(n_1909), .Y(n_1905) );
INVx1_ASAP7_75t_L g1937 ( .A(n_1938), .Y(n_1937) );
endmodule