module fake_jpeg_3058_n_555 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_555);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_555;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_10),
.B(n_4),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_52),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_59),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_28),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_60),
.Y(n_105)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_0),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_28),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_62),
.B(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_64),
.B(n_66),
.Y(n_165)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_19),
.B(n_1),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_69),
.B(n_90),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_70),
.Y(n_164)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_21),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_73),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_26),
.B(n_2),
.Y(n_79)
);

BUFx4f_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_37),
.B(n_2),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_87),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_34),
.B(n_18),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g149 ( 
.A(n_86),
.B(n_42),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_25),
.B(n_2),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_37),
.B(n_41),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_95),
.Y(n_127)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_41),
.B(n_2),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_46),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_98),
.B(n_104),
.Y(n_167)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_38),
.Y(n_122)
);

BUFx6f_ASAP7_75t_SL g102 ( 
.A(n_21),
.Y(n_102)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_48),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_78),
.A2(n_34),
.B1(n_51),
.B2(n_43),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_107),
.A2(n_126),
.B1(n_128),
.B2(n_162),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_50),
.B1(n_22),
.B2(n_43),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_111),
.A2(n_133),
.B1(n_15),
.B2(n_139),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_55),
.A2(n_34),
.B1(n_50),
.B2(n_22),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_115),
.A2(n_116),
.B1(n_141),
.B2(n_144),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_67),
.A2(n_50),
.B1(n_35),
.B2(n_22),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_53),
.A2(n_35),
.B1(n_43),
.B2(n_47),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_117),
.A2(n_159),
.B(n_17),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_122),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_65),
.A2(n_51),
.B1(n_35),
.B2(n_38),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_72),
.A2(n_47),
.B1(n_19),
.B2(n_40),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_59),
.A2(n_40),
.B1(n_27),
.B2(n_24),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_27),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_136),
.B(n_7),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_70),
.A2(n_24),
.B1(n_20),
.B2(n_21),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_79),
.A2(n_20),
.B1(n_21),
.B2(n_42),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_86),
.B(n_3),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_148),
.B(n_151),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_75),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_56),
.B(n_3),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_89),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_99),
.Y(n_183)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_52),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_156),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_91),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_54),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_81),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_163),
.A2(n_92),
.B1(n_101),
.B2(n_77),
.Y(n_200)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_168),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_111),
.A2(n_103),
.B1(n_82),
.B2(n_97),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_169),
.A2(n_186),
.B1(n_216),
.B2(n_226),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_170),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_54),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_171),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_109),
.B(n_76),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_172),
.B(n_181),
.Y(n_254)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_174),
.Y(n_268)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_175),
.Y(n_251)
);

INVx4_ASAP7_75t_SL g176 ( 
.A(n_121),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_176),
.B(n_222),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_177),
.B(n_191),
.Y(n_230)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_179),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_127),
.A2(n_100),
.B(n_94),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_180),
.B(n_187),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_124),
.B(n_119),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_183),
.Y(n_283)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_185),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_141),
.A2(n_88),
.B1(n_85),
.B2(n_96),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_105),
.B(n_71),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_165),
.B(n_80),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_189),
.B(n_205),
.Y(n_241)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_166),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_192),
.B(n_195),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_193),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_142),
.A2(n_102),
.B1(n_80),
.B2(n_101),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_194),
.A2(n_208),
.B1(n_146),
.B2(n_135),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_132),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_196),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_132),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_197),
.B(n_201),
.Y(n_260)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_128),
.A2(n_136),
.B(n_138),
.C(n_131),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_198),
.A2(n_107),
.B(n_162),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_199),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_200),
.A2(n_227),
.B1(n_207),
.B2(n_226),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_145),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_137),
.Y(n_202)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_202),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_112),
.B(n_74),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_203),
.B(n_143),
.C(n_158),
.Y(n_243)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_113),
.Y(n_204)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_204),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_68),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_129),
.Y(n_206)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_206),
.Y(n_281)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_134),
.A2(n_84),
.B(n_61),
.C(n_77),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_207),
.B(n_106),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_142),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_153),
.Y(n_209)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_209),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_210),
.B(n_215),
.Y(n_275)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_140),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_211),
.B(n_217),
.Y(n_261)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_212),
.Y(n_237)
);

AND2x4_ASAP7_75t_L g213 ( 
.A(n_160),
.B(n_18),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_214),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_114),
.B(n_8),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_152),
.B(n_9),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_116),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_123),
.B(n_9),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_125),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_218),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_161),
.B(n_9),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_219),
.B(n_213),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_123),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_220),
.B(n_221),
.Y(n_273)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_139),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_130),
.B(n_12),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_223),
.B(n_224),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_130),
.B(n_13),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_108),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_225),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_115),
.A2(n_17),
.B1(n_14),
.B2(n_15),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_163),
.A2(n_14),
.B1(n_15),
.B2(n_126),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_108),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_228),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_229),
.A2(n_164),
.B1(n_147),
.B2(n_135),
.Y(n_247)
);

AO21x1_ASAP7_75t_L g291 ( 
.A1(n_231),
.A2(n_255),
.B(n_265),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_198),
.A2(n_106),
.B(n_157),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_235),
.A2(n_234),
.B(n_231),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_229),
.A2(n_145),
.B1(n_150),
.B2(n_157),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_236),
.A2(n_246),
.B1(n_247),
.B2(n_252),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_242),
.B(n_249),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_243),
.B(n_245),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_245),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_184),
.A2(n_150),
.B1(n_158),
.B2(n_147),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_181),
.B(n_143),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_248),
.B(n_259),
.Y(n_289)
);

OAI32xp33_ASAP7_75t_L g249 ( 
.A1(n_172),
.A2(n_15),
.A3(n_170),
.B1(n_213),
.B2(n_182),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_170),
.A2(n_178),
.B1(n_171),
.B2(n_188),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_171),
.A2(n_221),
.B(n_203),
.Y(n_255)
);

AOI32xp33_ASAP7_75t_L g256 ( 
.A1(n_188),
.A2(n_189),
.A3(n_219),
.B1(n_192),
.B2(n_191),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_202),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_257),
.A2(n_258),
.B1(n_270),
.B2(n_284),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_178),
.A2(n_214),
.B1(n_227),
.B2(n_200),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_182),
.B(n_204),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_213),
.A2(n_220),
.B(n_214),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_262),
.A2(n_278),
.B(n_263),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_264),
.B(n_225),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_201),
.A2(n_213),
.B1(n_212),
.B2(n_196),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_206),
.A2(n_222),
.B1(n_209),
.B2(n_211),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_276),
.A2(n_218),
.B1(n_199),
.B2(n_195),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_190),
.B(n_173),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_175),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_199),
.A2(n_218),
.B1(n_185),
.B2(n_173),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_241),
.B(n_176),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_285),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_286),
.A2(n_268),
.B1(n_251),
.B2(n_271),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_241),
.B(n_176),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_287),
.B(n_292),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_272),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_288),
.Y(n_337)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_260),
.Y(n_290)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_290),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_291),
.A2(n_300),
.B(n_307),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_197),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_293),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_295),
.B(n_299),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_296),
.B(n_302),
.Y(n_356)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_297),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_280),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_298),
.B(n_304),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_242),
.A2(n_228),
.B1(n_174),
.B2(n_168),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_257),
.A2(n_179),
.B1(n_193),
.B2(n_254),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_301),
.A2(n_312),
.B1(n_282),
.B2(n_238),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_254),
.B(n_264),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_278),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_249),
.B(n_253),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_308),
.B(n_309),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_253),
.B(n_262),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_244),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_310),
.B(n_315),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_243),
.B(n_234),
.C(n_248),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_314),
.C(n_318),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_257),
.A2(n_258),
.B1(n_273),
.B2(n_252),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_239),
.A2(n_236),
.B1(n_247),
.B2(n_273),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_313),
.A2(n_327),
.B1(n_333),
.B2(n_282),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_243),
.B(n_255),
.C(n_259),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_256),
.B(n_230),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_277),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_317),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_253),
.B(n_262),
.C(n_244),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_253),
.B(n_230),
.C(n_232),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_319),
.A2(n_323),
.B(n_329),
.Y(n_369)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_281),
.Y(n_320)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_320),
.Y(n_338)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_276),
.Y(n_321)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_321),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_275),
.B(n_274),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_322),
.A2(n_328),
.B(n_330),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_232),
.B(n_261),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_272),
.Y(n_324)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_274),
.B(n_261),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_325),
.Y(n_354)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_326),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_239),
.A2(n_246),
.B1(n_270),
.B2(n_235),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_279),
.B(n_278),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_263),
.A2(n_250),
.B(n_233),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_331),
.A2(n_328),
.B(n_298),
.Y(n_374)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_267),
.Y(n_332)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_332),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_237),
.A2(n_284),
.B1(n_240),
.B2(n_233),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_279),
.B(n_266),
.Y(n_334)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_334),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_306),
.A2(n_237),
.B1(n_240),
.B2(n_250),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_336),
.A2(n_347),
.B1(n_350),
.B2(n_352),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g382 ( 
.A(n_351),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_306),
.A2(n_251),
.B1(n_238),
.B2(n_268),
.Y(n_352)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_297),
.Y(n_357)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_357),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_294),
.A2(n_268),
.B1(n_271),
.B2(n_269),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_358),
.Y(n_383)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_305),
.Y(n_360)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_312),
.A2(n_269),
.B1(n_271),
.B2(n_266),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_361),
.A2(n_365),
.B1(n_333),
.B2(n_321),
.Y(n_384)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_320),
.Y(n_362)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_362),
.Y(n_412)
);

AO22x1_ASAP7_75t_L g363 ( 
.A1(n_316),
.A2(n_301),
.B1(n_290),
.B2(n_293),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_377),
.Y(n_389)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_326),
.Y(n_364)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_364),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_327),
.A2(n_313),
.B1(n_303),
.B2(n_316),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_303),
.A2(n_316),
.B1(n_310),
.B2(n_300),
.Y(n_366)
);

INVxp33_ASAP7_75t_SL g413 ( 
.A(n_366),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_307),
.A2(n_291),
.B(n_329),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_368),
.A2(n_374),
.B(n_288),
.Y(n_407)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_332),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_370),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_308),
.A2(n_317),
.B1(n_302),
.B2(n_295),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_376),
.A2(n_356),
.B1(n_363),
.B2(n_375),
.Y(n_409)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_324),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_296),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_378),
.B(n_289),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_343),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_379),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_353),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_380),
.A2(n_409),
.B1(n_414),
.B2(n_355),
.Y(n_420)
);

INVx5_ASAP7_75t_L g381 ( 
.A(n_349),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_381),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_384),
.A2(n_388),
.B1(n_406),
.B2(n_375),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_354),
.B(n_322),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_386),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_292),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_387),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_365),
.A2(n_330),
.B1(n_309),
.B2(n_304),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_341),
.B(n_285),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_390),
.Y(n_424)
);

FAx1_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_291),
.CI(n_318),
.CON(n_392),
.SN(n_392)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_392),
.A2(n_407),
.B(n_411),
.Y(n_421)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_393),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_374),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_394),
.B(n_398),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_289),
.Y(n_396)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_396),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_331),
.Y(n_397)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_397),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_337),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_337),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_405),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_340),
.B(n_314),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_400),
.B(n_373),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_340),
.B(n_311),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_403),
.C(n_372),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_319),
.Y(n_403)
);

AO22x1_ASAP7_75t_SL g404 ( 
.A1(n_376),
.A2(n_336),
.B1(n_378),
.B2(n_352),
.Y(n_404)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_404),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_353),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_347),
.A2(n_323),
.B1(n_287),
.B2(n_288),
.Y(n_406)
);

XNOR2x2_ASAP7_75t_L g408 ( 
.A(n_339),
.B(n_286),
.Y(n_408)
);

MAJx2_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_360),
.C(n_357),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_371),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_410),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_373),
.A2(n_369),
.B(n_363),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_359),
.B(n_356),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_413),
.A2(n_361),
.B1(n_355),
.B2(n_339),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_416),
.A2(n_442),
.B1(n_394),
.B2(n_389),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_417),
.A2(n_420),
.B1(n_436),
.B2(n_441),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_401),
.B(n_371),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_422),
.B(n_393),
.Y(n_460)
);

NAND2x1_ASAP7_75t_L g426 ( 
.A(n_397),
.B(n_371),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_426),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_428),
.B(n_435),
.C(n_445),
.Y(n_462)
);

MAJx2_ASAP7_75t_L g448 ( 
.A(n_433),
.B(n_438),
.C(n_444),
.Y(n_448)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_395),
.Y(n_434)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_434),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_335),
.C(n_338),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_406),
.A2(n_342),
.B1(n_338),
.B2(n_335),
.Y(n_436)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_395),
.Y(n_439)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_439),
.Y(n_453)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_385),
.Y(n_440)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_440),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_396),
.A2(n_342),
.B1(n_362),
.B2(n_345),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_409),
.A2(n_345),
.B1(n_346),
.B2(n_364),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_385),
.Y(n_443)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_443),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_403),
.B(n_346),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_392),
.B(n_388),
.C(n_410),
.Y(n_445)
);

OAI211xp5_ASAP7_75t_SL g446 ( 
.A1(n_392),
.A2(n_370),
.B(n_344),
.C(n_377),
.Y(n_446)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_446),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_424),
.B(n_418),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_450),
.B(n_456),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_428),
.B(n_411),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g485 ( 
.A(n_452),
.B(n_421),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_454),
.A2(n_436),
.B1(n_429),
.B2(n_417),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_446),
.A2(n_407),
.B(n_389),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_455),
.A2(n_466),
.B(n_454),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_430),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_460),
.B(n_472),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_430),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_461),
.B(n_474),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_381),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_463),
.B(n_473),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_433),
.B(n_408),
.C(n_405),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_470),
.C(n_438),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_423),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_465),
.B(n_469),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_425),
.B(n_398),
.Y(n_467)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_467),
.Y(n_477)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_440),
.Y(n_468)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_468),
.Y(n_486)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_443),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_435),
.B(n_399),
.C(n_404),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_434),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_471),
.B(n_415),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_444),
.B(n_404),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_437),
.B(n_391),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_427),
.B(n_447),
.Y(n_474)
);

NAND3xp33_ASAP7_75t_L g500 ( 
.A(n_475),
.B(n_491),
.C(n_448),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_449),
.A2(n_416),
.B1(n_431),
.B2(n_447),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_476),
.B(n_485),
.Y(n_511)
);

AOI322xp5_ASAP7_75t_L g478 ( 
.A1(n_465),
.A2(n_427),
.A3(n_431),
.B1(n_467),
.B2(n_429),
.C1(n_451),
.C2(n_453),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_478),
.B(n_412),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_451),
.B(n_439),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_479),
.B(n_488),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g480 ( 
.A(n_460),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_480),
.B(n_481),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_422),
.C(n_445),
.Y(n_481)
);

INVxp33_ASAP7_75t_L g482 ( 
.A(n_459),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_482),
.B(n_493),
.Y(n_510)
);

OAI21xp33_ASAP7_75t_L g484 ( 
.A1(n_464),
.A2(n_421),
.B(n_423),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_484),
.A2(n_383),
.B(n_457),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_492),
.Y(n_507)
);

OA21x2_ASAP7_75t_SL g493 ( 
.A1(n_459),
.A2(n_426),
.B(n_442),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_495),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_466),
.A2(n_383),
.B1(n_384),
.B2(n_419),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_453),
.B(n_419),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_496),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_481),
.B(n_462),
.C(n_470),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_497),
.B(n_499),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_490),
.A2(n_455),
.B(n_471),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_500),
.A2(n_506),
.B1(n_514),
.B2(n_486),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_475),
.B(n_448),
.C(n_452),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_501),
.B(n_503),
.C(n_504),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_483),
.B(n_472),
.C(n_426),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_483),
.B(n_402),
.C(n_468),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_477),
.A2(n_469),
.B1(n_458),
.B2(n_457),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_488),
.B(n_402),
.C(n_458),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_513),
.C(n_486),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_495),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_492),
.B(n_344),
.C(n_391),
.Y(n_513)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_502),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_515),
.A2(n_523),
.B1(n_524),
.B2(n_525),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_517),
.B(n_521),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_509),
.B(n_489),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_518),
.B(n_497),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_502),
.B(n_479),
.Y(n_519)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_519),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_510),
.B(n_489),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_520),
.A2(n_522),
.B1(n_526),
.B2(n_505),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_498),
.A2(n_493),
.B(n_477),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_498),
.A2(n_487),
.B(n_496),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_513),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_507),
.A2(n_476),
.B1(n_487),
.B2(n_494),
.Y(n_525)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_508),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_527),
.B(n_507),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_529),
.B(n_531),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_530),
.A2(n_533),
.B(n_517),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_504),
.C(n_501),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g535 ( 
.A(n_521),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_535),
.B(n_537),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_523),
.B(n_505),
.C(n_503),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_520),
.B(n_511),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_538),
.B(n_516),
.Y(n_541)
);

AO21x1_ASAP7_75t_L g548 ( 
.A1(n_541),
.A2(n_544),
.B(n_536),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_537),
.B(n_527),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_542),
.B(n_543),
.Y(n_547)
);

XNOR2x1_ASAP7_75t_L g543 ( 
.A(n_534),
.B(n_516),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_539),
.A2(n_534),
.B(n_532),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_545),
.B(n_546),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_539),
.A2(n_532),
.B(n_519),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_547),
.Y(n_549)
);

OAI321xp33_ASAP7_75t_L g551 ( 
.A1(n_549),
.A2(n_540),
.A3(n_522),
.B1(n_515),
.B2(n_525),
.C(n_524),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_551),
.B(n_552),
.C(n_485),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_550),
.A2(n_511),
.B(n_412),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_553),
.B(n_415),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_554),
.B(n_382),
.Y(n_555)
);


endmodule