module fake_jpeg_4223_n_178 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_37),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_36),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_22),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_31),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_24),
.B1(n_28),
.B2(n_20),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_28),
.B1(n_27),
.B2(n_21),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_28),
.B1(n_14),
.B2(n_22),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_14),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_27),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_55),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_54),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_60),
.B1(n_18),
.B2(n_19),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_62),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_16),
.B1(n_17),
.B2(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_64),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_17),
.B1(n_26),
.B2(n_14),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_22),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_20),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_68),
.B(n_69),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_21),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_23),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_31),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_82),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_74),
.B(n_90),
.Y(n_100)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_88),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_42),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_52),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_31),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_39),
.B1(n_15),
.B2(n_23),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_34),
.B(n_42),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_87),
.A2(n_69),
.B(n_68),
.Y(n_97)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_92),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_30),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_61),
.B1(n_42),
.B2(n_58),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_108),
.B1(n_90),
.B2(n_73),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_74),
.A2(n_69),
.B1(n_68),
.B2(n_67),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_81),
.C(n_79),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_97),
.A2(n_99),
.B(n_107),
.Y(n_118)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_102),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_77),
.B(n_52),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_38),
.Y(n_103)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_39),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_77),
.B(n_19),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_111),
.Y(n_120)
);

AO22x1_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_32),
.B1(n_39),
.B2(n_23),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_15),
.B(n_1),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_121),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_127),
.B1(n_100),
.B2(n_112),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_82),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_97),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_107),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_128),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_126),
.C(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_83),
.B1(n_77),
.B2(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_109),
.B(n_92),
.Y(n_126)
);

AO21x2_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_72),
.B(n_88),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_104),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_133),
.C(n_138),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_110),
.C(n_100),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_140),
.B1(n_135),
.B2(n_130),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_96),
.C(n_102),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_141),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_106),
.B(n_85),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_108),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_111),
.C(n_95),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_118),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_147),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_136),
.A2(n_127),
.B1(n_129),
.B2(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

AOI322xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_127),
.A3(n_125),
.B1(n_115),
.B2(n_120),
.C1(n_117),
.C2(n_15),
.Y(n_147)
);

AOI322xp5_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_127),
.A3(n_15),
.B1(n_89),
.B2(n_78),
.C1(n_8),
.C2(n_10),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_151),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_149),
.B(n_3),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_3),
.B(n_4),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_132),
.B(n_10),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_133),
.B1(n_139),
.B2(n_131),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_155),
.B(n_157),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_11),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_150),
.A2(n_3),
.B(n_4),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_9),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_160),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_157),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_146),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_163),
.B(n_164),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_146),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_4),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_166),
.A2(n_156),
.B(n_144),
.C(n_6),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_169),
.B(n_170),
.Y(n_174)
);

AOI31xp33_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_144),
.A3(n_6),
.B(n_7),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_5),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_168),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_173),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_169),
.B(n_163),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_6),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_175),
.Y(n_178)
);


endmodule